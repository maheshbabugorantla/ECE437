/*
  Mahesh Babu Gorantla
  mgorantl@purdue.edu

  holds datapath request_unit interface signals
*/
`ifndef REQUEST_UNIT_IF_VH
`define REQUEST_UNIT_IF_VH

// types
`include "cpu_types_pkg.vh"

interface request_control_if;

	// import types
	import cpu_types_pkg::*;

		


endinterface

`endif