// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 64-Bit"
// VERSION "Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"

// DATE "08/29/2017 07:59:39"

// 
// Device: Altera EP4CE115F29C8 Package FBGA780
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module register_file (
	clk,
	n_rst,
	\my_rf.rdat2 ,
	\my_rf.rdat1 ,
	\my_rf.wdat ,
	\my_rf.rsel2 ,
	\my_rf.rsel1 ,
	\my_rf.wsel ,
	\my_rf.WEN );
input 	clk;
input 	n_rst;
output 	[31:0] \my_rf.rdat2 ;
output 	[31:0] \my_rf.rdat1 ;
input 	[31:0] \my_rf.wdat ;
input 	[4:0] \my_rf.rsel2 ;
input 	[4:0] \my_rf.rsel1 ;
input 	[4:0] \my_rf.wsel ;
input 	\my_rf.WEN ;

// Design Ports Information
// my_rf.rdat2[0]	=>  Location: PIN_C14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[1]	=>  Location: PIN_AD15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[2]	=>  Location: PIN_AE16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[3]	=>  Location: PIN_P2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[4]	=>  Location: PIN_AG17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[5]	=>  Location: PIN_AB2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[6]	=>  Location: PIN_E15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[7]	=>  Location: PIN_C15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[8]	=>  Location: PIN_C13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[9]	=>  Location: PIN_A17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[10]	=>  Location: PIN_N8,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[11]	=>  Location: PIN_D13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[12]	=>  Location: PIN_AC15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[13]	=>  Location: PIN_AF15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[14]	=>  Location: PIN_AE11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[15]	=>  Location: PIN_H13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[16]	=>  Location: PIN_L2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[17]	=>  Location: PIN_F12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[18]	=>  Location: PIN_AG10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[19]	=>  Location: PIN_C12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[20]	=>  Location: PIN_L1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[21]	=>  Location: PIN_U6,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[22]	=>  Location: PIN_AF11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[23]	=>  Location: PIN_Y4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[24]	=>  Location: PIN_AD14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[25]	=>  Location: PIN_AE12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[26]	=>  Location: PIN_B10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[27]	=>  Location: PIN_U2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[28]	=>  Location: PIN_G13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[29]	=>  Location: PIN_B11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[30]	=>  Location: PIN_N4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat2[31]	=>  Location: PIN_J12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[0]	=>  Location: PIN_F15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[1]	=>  Location: PIN_M8,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[2]	=>  Location: PIN_AH17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[3]	=>  Location: PIN_H14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[4]	=>  Location: PIN_AF10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[5]	=>  Location: PIN_D14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[6]	=>  Location: PIN_H15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[7]	=>  Location: PIN_AE15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[8]	=>  Location: PIN_D15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[9]	=>  Location: PIN_B17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[10]	=>  Location: PIN_J14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[11]	=>  Location: PIN_P21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[12]	=>  Location: PIN_U1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[13]	=>  Location: PIN_AA16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[14]	=>  Location: PIN_M7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[15]	=>  Location: PIN_D10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[16]	=>  Location: PIN_AB1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[17]	=>  Location: PIN_A12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[18]	=>  Location: PIN_F14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[19]	=>  Location: PIN_W1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[20]	=>  Location: PIN_AE9,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[21]	=>  Location: PIN_AE10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[22]	=>  Location: PIN_M1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[23]	=>  Location: PIN_P1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[24]	=>  Location: PIN_W2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[25]	=>  Location: PIN_C10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[26]	=>  Location: PIN_M2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[27]	=>  Location: PIN_J13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[28]	=>  Location: PIN_A10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[29]	=>  Location: PIN_AB11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[30]	=>  Location: PIN_AF16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rdat1[31]	=>  Location: PIN_A11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rsel2[3]	=>  Location: PIN_V2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rsel2[2]	=>  Location: PIN_AB14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rsel2[0]	=>  Location: PIN_D12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rsel2[1]	=>  Location: PIN_V4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rsel2[4]	=>  Location: PIN_R1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rsel1[3]	=>  Location: PIN_AH12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rsel1[2]	=>  Location: PIN_V3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rsel1[0]	=>  Location: PIN_AG11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rsel1[1]	=>  Location: PIN_AH11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.rsel1[4]	=>  Location: PIN_AC10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[0]	=>  Location: PIN_AC14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// clk	=>  Location: PIN_J1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// n_rst	=>  Location: PIN_Y2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wsel[3]	=>  Location: PIN_AH10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wsel[4]	=>  Location: PIN_AF12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wsel[0]	=>  Location: PIN_T7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.WEN	=>  Location: PIN_U5,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wsel[1]	=>  Location: PIN_Y3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wsel[2]	=>  Location: PIN_V1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[1]	=>  Location: PIN_AA14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[2]	=>  Location: PIN_Y12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[3]	=>  Location: PIN_AF14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[4]	=>  Location: PIN_AE14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[5]	=>  Location: PIN_AD11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[6]	=>  Location: PIN_Y15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[7]	=>  Location: PIN_AG12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[8]	=>  Location: PIN_Y14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[9]	=>  Location: PIN_AA13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[10]	=>  Location: PIN_AD12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[11]	=>  Location: PIN_U3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[12]	=>  Location: PIN_R6,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[13]	=>  Location: PIN_AB13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[14]	=>  Location: PIN_T3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[15]	=>  Location: PIN_AA12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[16]	=>  Location: PIN_R2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[17]	=>  Location: PIN_AB12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[18]	=>  Location: PIN_AC12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[19]	=>  Location: PIN_AC11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[20]	=>  Location: PIN_G14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[21]	=>  Location: PIN_R5,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[22]	=>  Location: PIN_E14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[23]	=>  Location: PIN_U4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[24]	=>  Location: PIN_AE13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[25]	=>  Location: PIN_T4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[26]	=>  Location: PIN_R3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[27]	=>  Location: PIN_AB10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[28]	=>  Location: PIN_R7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[29]	=>  Location: PIN_R4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[30]	=>  Location: PIN_AF13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// my_rf.wdat[31]	=>  Location: PIN_Y13,	 I/O Standard: 2.5 V,	 Current Strength: Default


wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
wire \registerArray[25][0]~q ;
wire \registerArray[26][0]~q ;
wire \registerArray[18][0]~q ;
wire \Mux63~2_combout ;
wire \registerArray[24][0]~q ;
wire \registerArray[16][0]~q ;
wire \Mux63~4_combout ;
wire \registerArray[23][0]~q ;
wire \registerArray[19][0]~q ;
wire \Mux63~7_combout ;
wire \Mux63~8_combout ;
wire \registerArray[6][0]~q ;
wire \registerArray[5][0]~q ;
wire \registerArray[4][0]~q ;
wire \Mux63~12_combout ;
wire \registerArray[7][0]~q ;
wire \Mux63~13_combout ;
wire \registerArray[3][0]~q ;
wire \registerArray[1][0]~q ;
wire \Mux63~14_combout ;
wire \registerArray[2][0]~q ;
wire \Mux63~15_combout ;
wire \Mux63~16_combout ;
wire \registerArray[21][1]~q ;
wire \registerArray[25][1]~q ;
wire \registerArray[17][1]~q ;
wire \Mux62~0_combout ;
wire \registerArray[29][1]~q ;
wire \Mux62~1_combout ;
wire \registerArray[18][1]~q ;
wire \registerArray[27][1]~q ;
wire \registerArray[19][1]~q ;
wire \Mux62~7_combout ;
wire \registerArray[9][1]~q ;
wire \registerArray[10][1]~q ;
wire \registerArray[8][1]~q ;
wire \Mux62~12_combout ;
wire \registerArray[11][1]~q ;
wire \Mux62~13_combout ;
wire \registerArray[3][1]~q ;
wire \registerArray[1][1]~q ;
wire \Mux62~14_combout ;
wire \registerArray[2][1]~q ;
wire \Mux62~15_combout ;
wire \Mux62~16_combout ;
wire \registerArray[22][2]~q ;
wire \registerArray[26][2]~q ;
wire \registerArray[18][2]~q ;
wire \Mux61~2_combout ;
wire \registerArray[30][2]~q ;
wire \Mux61~3_combout ;
wire \Mux61~4_combout ;
wire \Mux61~5_combout ;
wire \Mux61~6_combout ;
wire \registerArray[10][2]~q ;
wire \registerArray[8][2]~q ;
wire \Mux61~10_combout ;
wire \Mux61~11_combout ;
wire \registerArray[4][2]~q ;
wire \registerArray[7][2]~q ;
wire \registerArray[1][2]~q ;
wire \registerArray[13][2]~q ;
wire \registerArray[12][2]~q ;
wire \Mux61~17_combout ;
wire \registerArray[17][3]~q ;
wire \registerArray[22][3]~q ;
wire \registerArray[18][3]~q ;
wire \Mux60~2_combout ;
wire \Mux60~3_combout ;
wire \registerArray[20][3]~q ;
wire \registerArray[16][3]~q ;
wire \Mux60~4_combout ;
wire \Mux60~5_combout ;
wire \Mux60~6_combout ;
wire \Mux60~10_combout ;
wire \registerArray[8][3]~q ;
wire \registerArray[11][3]~q ;
wire \registerArray[1][3]~q ;
wire \registerArray[22][4]~q ;
wire \registerArray[26][4]~q ;
wire \registerArray[18][4]~q ;
wire \Mux59~2_combout ;
wire \registerArray[30][4]~q ;
wire \Mux59~3_combout ;
wire \Mux59~7_combout ;
wire \registerArray[6][4]~q ;
wire \registerArray[5][4]~q ;
wire \registerArray[4][4]~q ;
wire \Mux59~12_combout ;
wire \registerArray[7][4]~q ;
wire \Mux59~13_combout ;
wire \Mux59~14_combout ;
wire \Mux59~15_combout ;
wire \Mux59~16_combout ;
wire \registerArray[21][5]~q ;
wire \registerArray[18][5]~q ;
wire \registerArray[5][5]~q ;
wire \registerArray[4][5]~q ;
wire \Mux58~10_combout ;
wire \Mux58~11_combout ;
wire \registerArray[9][5]~q ;
wire \Mux58~12_combout ;
wire \Mux58~13_combout ;
wire \Mux58~14_combout ;
wire \Mux57~0_combout ;
wire \Mux57~1_combout ;
wire \Mux57~2_combout ;
wire \Mux57~3_combout ;
wire \registerArray[31][6]~q ;
wire \registerArray[5][6]~q ;
wire \registerArray[4][6]~q ;
wire \Mux57~12_combout ;
wire \registerArray[3][6]~q ;
wire \registerArray[1][6]~q ;
wire \Mux57~14_combout ;
wire \registerArray[2][6]~q ;
wire \Mux57~15_combout ;
wire \Mux57~17_combout ;
wire \Mux57~18_combout ;
wire \registerArray[25][7]~q ;
wire \registerArray[17][7]~q ;
wire \Mux56~0_combout ;
wire \Mux56~1_combout ;
wire \registerArray[28][7]~q ;
wire \Mux56~7_combout ;
wire \registerArray[4][7]~q ;
wire \registerArray[10][7]~q ;
wire \registerArray[8][7]~q ;
wire \Mux56~12_combout ;
wire \Mux56~13_combout ;
wire \registerArray[14][7]~q ;
wire \registerArray[13][7]~q ;
wire \registerArray[12][7]~q ;
wire \Mux56~17_combout ;
wire \registerArray[15][7]~q ;
wire \Mux56~18_combout ;
wire \Mux55~2_combout ;
wire \Mux55~4_combout ;
wire \registerArray[27][8]~q ;
wire \registerArray[23][8]~q ;
wire \Mux55~7_combout ;
wire \Mux55~8_combout ;
wire \registerArray[8][8]~q ;
wire \registerArray[4][8]~q ;
wire \Mux55~14_combout ;
wire \Mux54~0_combout ;
wire \registerArray[19][9]~q ;
wire \registerArray[5][9]~q ;
wire \registerArray[4][9]~q ;
wire \Mux54~10_combout ;
wire \registerArray[9][9]~q ;
wire \registerArray[10][9]~q ;
wire \registerArray[8][9]~q ;
wire \Mux54~12_combout ;
wire \registerArray[11][9]~q ;
wire \Mux54~13_combout ;
wire \Mux54~14_combout ;
wire \registerArray[14][9]~q ;
wire \registerArray[13][9]~q ;
wire \registerArray[12][9]~q ;
wire \Mux54~17_combout ;
wire \registerArray[15][9]~q ;
wire \Mux54~18_combout ;
wire \registerArray[25][10]~q ;
wire \registerArray[21][10]~q ;
wire \registerArray[17][10]~q ;
wire \Mux53~0_combout ;
wire \registerArray[29][10]~q ;
wire \Mux53~1_combout ;
wire \registerArray[22][10]~q ;
wire \registerArray[26][10]~q ;
wire \registerArray[18][10]~q ;
wire \Mux53~2_combout ;
wire \registerArray[30][10]~q ;
wire \Mux53~3_combout ;
wire \registerArray[10][10]~q ;
wire \registerArray[8][10]~q ;
wire \Mux53~10_combout ;
wire \Mux53~11_combout ;
wire \registerArray[21][11]~q ;
wire \registerArray[25][11]~q ;
wire \Mux52~0_combout ;
wire \Mux52~1_combout ;
wire \registerArray[24][11]~q ;
wire \Mux52~4_combout ;
wire \Mux52~5_combout ;
wire \registerArray[10][11]~q ;
wire \registerArray[8][11]~q ;
wire \Mux52~12_combout ;
wire \registerArray[13][11]~q ;
wire \registerArray[12][11]~q ;
wire \Mux52~17_combout ;
wire \Mux52~18_combout ;
wire \registerArray[21][12]~q ;
wire \Mux51~0_combout ;
wire \registerArray[22][12]~q ;
wire \registerArray[26][12]~q ;
wire \registerArray[18][12]~q ;
wire \Mux51~2_combout ;
wire \registerArray[30][12]~q ;
wire \Mux51~3_combout ;
wire \registerArray[23][12]~q ;
wire \Mux51~7_combout ;
wire \Mux51~8_combout ;
wire \registerArray[10][12]~q ;
wire \registerArray[8][12]~q ;
wire \Mux51~10_combout ;
wire \registerArray[7][12]~q ;
wire \Mux51~14_combout ;
wire \Mux51~15_combout ;
wire \registerArray[25][13]~q ;
wire \registerArray[17][13]~q ;
wire \Mux50~0_combout ;
wire \Mux50~1_combout ;
wire \Mux50~2_combout ;
wire \registerArray[24][13]~q ;
wire \Mux50~4_combout ;
wire \Mux50~5_combout ;
wire \registerArray[9][13]~q ;
wire \registerArray[10][13]~q ;
wire \registerArray[8][13]~q ;
wire \Mux50~12_combout ;
wire \registerArray[11][13]~q ;
wire \Mux50~13_combout ;
wire \registerArray[3][13]~q ;
wire \registerArray[1][13]~q ;
wire \Mux50~14_combout ;
wire \registerArray[2][13]~q ;
wire \Mux50~15_combout ;
wire \Mux50~16_combout ;
wire \registerArray[30][14]~q ;
wire \registerArray[28][14]~q ;
wire \registerArray[23][14]~q ;
wire \registerArray[19][14]~q ;
wire \Mux49~7_combout ;
wire \Mux49~10_combout ;
wire \registerArray[5][14]~q ;
wire \registerArray[4][14]~q ;
wire \Mux49~12_combout ;
wire \Mux49~13_combout ;
wire \Mux49~14_combout ;
wire \Mux49~15_combout ;
wire \Mux49~16_combout ;
wire \registerArray[12][14]~q ;
wire \Mux48~2_combout ;
wire \registerArray[28][15]~q ;
wire \registerArray[31][15]~q ;
wire \registerArray[9][15]~q ;
wire \registerArray[10][15]~q ;
wire \registerArray[8][15]~q ;
wire \Mux48~12_combout ;
wire \registerArray[11][15]~q ;
wire \Mux48~13_combout ;
wire \registerArray[13][15]~q ;
wire \registerArray[12][15]~q ;
wire \Mux48~17_combout ;
wire \Mux48~18_combout ;
wire \Mux47~2_combout ;
wire \registerArray[24][16]~q ;
wire \registerArray[16][16]~q ;
wire \Mux47~4_combout ;
wire \Mux47~5_combout ;
wire \registerArray[27][16]~q ;
wire \registerArray[23][16]~q ;
wire \registerArray[19][16]~q ;
wire \Mux47~7_combout ;
wire \registerArray[31][16]~q ;
wire \Mux47~8_combout ;
wire \Mux47~10_combout ;
wire \registerArray[6][16]~q ;
wire \registerArray[5][16]~q ;
wire \registerArray[4][16]~q ;
wire \Mux47~12_combout ;
wire \registerArray[7][16]~q ;
wire \Mux47~13_combout ;
wire \Mux47~14_combout ;
wire \Mux47~15_combout ;
wire \Mux47~16_combout ;
wire \registerArray[13][16]~q ;
wire \registerArray[12][16]~q ;
wire \Mux47~17_combout ;
wire \registerArray[25][17]~q ;
wire \registerArray[17][17]~q ;
wire \Mux46~0_combout ;
wire \Mux46~4_combout ;
wire \Mux46~5_combout ;
wire \registerArray[27][17]~q ;
wire \registerArray[19][17]~q ;
wire \Mux46~7_combout ;
wire \Mux46~8_combout ;
wire \registerArray[5][17]~q ;
wire \registerArray[4][17]~q ;
wire \Mux46~10_combout ;
wire \registerArray[9][17]~q ;
wire \registerArray[10][17]~q ;
wire \registerArray[8][17]~q ;
wire \Mux46~12_combout ;
wire \registerArray[11][17]~q ;
wire \Mux46~13_combout ;
wire \registerArray[3][17]~q ;
wire \Mux46~14_combout ;
wire \Mux46~15_combout ;
wire \Mux46~16_combout ;
wire \registerArray[13][17]~q ;
wire \registerArray[12][17]~q ;
wire \Mux46~17_combout ;
wire \registerArray[24][18]~q ;
wire \registerArray[16][18]~q ;
wire \Mux45~4_combout ;
wire \registerArray[10][18]~q ;
wire \registerArray[8][18]~q ;
wire \Mux45~10_combout ;
wire \registerArray[4][18]~q ;
wire \registerArray[7][18]~q ;
wire \registerArray[26][19]~q ;
wire \registerArray[22][19]~q ;
wire \registerArray[18][19]~q ;
wire \Mux44~2_combout ;
wire \registerArray[30][19]~q ;
wire \Mux44~3_combout ;
wire \registerArray[24][19]~q ;
wire \Mux44~4_combout ;
wire \Mux44~5_combout ;
wire \Mux44~6_combout ;
wire \registerArray[27][19]~q ;
wire \registerArray[19][19]~q ;
wire \Mux44~7_combout ;
wire \registerArray[8][19]~q ;
wire \registerArray[11][19]~q ;
wire \registerArray[1][19]~q ;
wire \registerArray[17][20]~q ;
wire \registerArray[26][20]~q ;
wire \registerArray[18][20]~q ;
wire \Mux43~2_combout ;
wire \Mux43~3_combout ;
wire \registerArray[20][20]~q ;
wire \Mux43~4_combout ;
wire \Mux43~5_combout ;
wire \Mux43~6_combout ;
wire \registerArray[3][20]~q ;
wire \registerArray[1][20]~q ;
wire \Mux43~14_combout ;
wire \Mux43~15_combout ;
wire \registerArray[13][20]~q ;
wire \registerArray[12][20]~q ;
wire \Mux43~17_combout ;
wire \Mux43~18_combout ;
wire \registerArray[21][21]~q ;
wire \Mux42~0_combout ;
wire \Mux42~1_combout ;
wire \registerArray[24][21]~q ;
wire \Mux42~4_combout ;
wire \Mux42~5_combout ;
wire \registerArray[10][21]~q ;
wire \registerArray[8][21]~q ;
wire \Mux42~12_combout ;
wire \Mux42~14_combout ;
wire \registerArray[13][21]~q ;
wire \registerArray[12][21]~q ;
wire \Mux42~17_combout ;
wire \registerArray[22][22]~q ;
wire \registerArray[26][22]~q ;
wire \registerArray[18][22]~q ;
wire \Mux41~2_combout ;
wire \registerArray[30][22]~q ;
wire \Mux41~3_combout ;
wire \registerArray[20][22]~q ;
wire \registerArray[24][22]~q ;
wire \registerArray[16][22]~q ;
wire \Mux41~4_combout ;
wire \registerArray[28][22]~q ;
wire \Mux41~5_combout ;
wire \Mux41~6_combout ;
wire \registerArray[19][22]~q ;
wire \registerArray[3][22]~q ;
wire \registerArray[1][22]~q ;
wire \Mux41~14_combout ;
wire \registerArray[13][22]~q ;
wire \registerArray[12][22]~q ;
wire \Mux41~17_combout ;
wire \registerArray[25][23]~q ;
wire \registerArray[17][23]~q ;
wire \Mux40~0_combout ;
wire \registerArray[22][23]~q ;
wire \registerArray[18][23]~q ;
wire \Mux40~2_combout ;
wire \Mux40~3_combout ;
wire \registerArray[24][23]~q ;
wire \registerArray[20][23]~q ;
wire \registerArray[16][23]~q ;
wire \Mux40~4_combout ;
wire \registerArray[28][23]~q ;
wire \Mux40~5_combout ;
wire \Mux40~6_combout ;
wire \Mux40~12_combout ;
wire \Mux40~13_combout ;
wire \registerArray[3][23]~q ;
wire \registerArray[1][23]~q ;
wire \Mux40~14_combout ;
wire \registerArray[2][23]~q ;
wire \Mux40~15_combout ;
wire \Mux40~16_combout ;
wire \Mux39~0_combout ;
wire \registerArray[22][24]~q ;
wire \registerArray[26][24]~q ;
wire \registerArray[18][24]~q ;
wire \Mux39~2_combout ;
wire \registerArray[30][24]~q ;
wire \Mux39~3_combout ;
wire \registerArray[28][24]~q ;
wire \registerArray[23][24]~q ;
wire \registerArray[19][24]~q ;
wire \Mux39~7_combout ;
wire \Mux39~8_combout ;
wire \registerArray[8][24]~q ;
wire \Mux39~14_combout ;
wire \Mux39~15_combout ;
wire \registerArray[13][24]~q ;
wire \registerArray[12][24]~q ;
wire \Mux39~17_combout ;
wire \Mux39~18_combout ;
wire \registerArray[20][25]~q ;
wire \registerArray[16][25]~q ;
wire \Mux38~4_combout ;
wire \Mux38~5_combout ;
wire \Mux38~7_combout ;
wire \Mux38~8_combout ;
wire \registerArray[4][25]~q ;
wire \registerArray[11][25]~q ;
wire \registerArray[25][26]~q ;
wire \registerArray[22][26]~q ;
wire \registerArray[26][26]~q ;
wire \registerArray[18][26]~q ;
wire \Mux37~2_combout ;
wire \registerArray[30][26]~q ;
wire \Mux37~3_combout ;
wire \registerArray[24][26]~q ;
wire \registerArray[16][26]~q ;
wire \Mux37~4_combout ;
wire \Mux37~5_combout ;
wire \Mux37~6_combout ;
wire \registerArray[23][26]~q ;
wire \registerArray[19][26]~q ;
wire \Mux37~7_combout ;
wire \registerArray[9][26]~q ;
wire \registerArray[10][26]~q ;
wire \registerArray[8][26]~q ;
wire \Mux37~10_combout ;
wire \registerArray[11][26]~q ;
wire \Mux37~11_combout ;
wire \registerArray[4][26]~q ;
wire \registerArray[12][26]~q ;
wire \registerArray[21][27]~q ;
wire \registerArray[26][27]~q ;
wire \registerArray[22][27]~q ;
wire \registerArray[18][27]~q ;
wire \Mux36~2_combout ;
wire \registerArray[30][27]~q ;
wire \Mux36~3_combout ;
wire \registerArray[28][27]~q ;
wire \Mux36~7_combout ;
wire \Mux36~8_combout ;
wire \registerArray[8][27]~q ;
wire \registerArray[11][27]~q ;
wire \Mux36~17_combout ;
wire \Mux35~0_combout ;
wire \Mux35~2_combout ;
wire \Mux35~3_combout ;
wire \registerArray[27][28]~q ;
wire \registerArray[23][28]~q ;
wire \registerArray[19][28]~q ;
wire \Mux35~7_combout ;
wire \registerArray[31][28]~q ;
wire \Mux35~8_combout ;
wire \registerArray[13][28]~q ;
wire \registerArray[12][28]~q ;
wire \Mux35~17_combout ;
wire \Mux34~0_combout ;
wire \Mux34~1_combout ;
wire \registerArray[22][29]~q ;
wire \registerArray[18][29]~q ;
wire \Mux34~2_combout ;
wire \registerArray[20][29]~q ;
wire \Mux34~4_combout ;
wire \Mux34~5_combout ;
wire \registerArray[4][29]~q ;
wire \registerArray[12][29]~q ;
wire \registerArray[15][29]~q ;
wire \registerArray[21][30]~q ;
wire \registerArray[17][30]~q ;
wire \Mux33~0_combout ;
wire \Mux33~1_combout ;
wire \registerArray[18][30]~q ;
wire \registerArray[24][30]~q ;
wire \registerArray[16][30]~q ;
wire \Mux33~4_combout ;
wire \registerArray[11][30]~q ;
wire \registerArray[5][30]~q ;
wire \registerArray[4][30]~q ;
wire \Mux33~12_combout ;
wire \Mux33~13_combout ;
wire \registerArray[3][30]~q ;
wire \registerArray[1][30]~q ;
wire \Mux33~14_combout ;
wire \registerArray[2][30]~q ;
wire \Mux33~15_combout ;
wire \Mux33~16_combout ;
wire \registerArray[21][31]~q ;
wire \registerArray[26][31]~q ;
wire \registerArray[22][31]~q ;
wire \registerArray[18][31]~q ;
wire \Mux32~2_combout ;
wire \registerArray[30][31]~q ;
wire \Mux32~3_combout ;
wire \Mux32~4_combout ;
wire \Mux32~5_combout ;
wire \Mux32~6_combout ;
wire \registerArray[27][31]~q ;
wire \registerArray[19][31]~q ;
wire \Mux32~7_combout ;
wire \Mux32~10_combout ;
wire \Mux32~11_combout ;
wire \registerArray[9][31]~q ;
wire \registerArray[10][31]~q ;
wire \registerArray[8][31]~q ;
wire \Mux32~12_combout ;
wire \registerArray[11][31]~q ;
wire \Mux32~13_combout ;
wire \registerArray[1][31]~q ;
wire \registerArray[15][31]~q ;
wire \Mux31~0_combout ;
wire \Mux31~1_combout ;
wire \Mux31~2_combout ;
wire \Mux31~3_combout ;
wire \Mux31~4_combout ;
wire \Mux31~7_combout ;
wire \Mux31~10_combout ;
wire \Mux31~12_combout ;
wire \Mux31~13_combout ;
wire \Mux31~14_combout ;
wire \Mux31~15_combout ;
wire \Mux31~16_combout ;
wire \Mux31~17_combout ;
wire \Mux30~0_combout ;
wire \Mux30~1_combout ;
wire \Mux30~2_combout ;
wire \Mux30~4_combout ;
wire \Mux30~5_combout ;
wire \Mux30~7_combout ;
wire \Mux30~12_combout ;
wire \Mux30~13_combout ;
wire \Mux30~14_combout ;
wire \Mux30~15_combout ;
wire \Mux30~16_combout ;
wire \Mux29~0_combout ;
wire \Mux29~2_combout ;
wire \Mux29~3_combout ;
wire \Mux29~7_combout ;
wire \Mux29~8_combout ;
wire \Mux29~10_combout ;
wire \Mux29~12_combout ;
wire \Mux29~13_combout ;
wire \Mux29~14_combout ;
wire \Mux29~15_combout ;
wire \Mux29~16_combout ;
wire \Mux29~17_combout ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \Mux28~2_combout ;
wire \Mux28~4_combout ;
wire \Mux28~7_combout ;
wire \Mux28~12_combout ;
wire \Mux28~13_combout ;
wire \Mux28~14_combout ;
wire \Mux28~17_combout ;
wire \Mux27~2_combout ;
wire \Mux27~3_combout ;
wire \Mux27~12_combout ;
wire \Mux27~13_combout ;
wire \Mux27~17_combout ;
wire \Mux27~18_combout ;
wire \Mux26~2_combout ;
wire \Mux26~10_combout ;
wire \Mux25~7_combout ;
wire \Mux25~8_combout ;
wire \Mux25~12_combout ;
wire \Mux25~13_combout ;
wire \Mux25~14_combout ;
wire \Mux25~15_combout ;
wire \Mux25~16_combout ;
wire \Mux24~0_combout ;
wire \Mux24~2_combout ;
wire \Mux24~3_combout ;
wire \Mux24~4_combout ;
wire \Mux24~5_combout ;
wire \Mux24~6_combout ;
wire \Mux24~10_combout ;
wire \Mux24~12_combout ;
wire \Mux24~17_combout ;
wire \Mux24~18_combout ;
wire \Mux23~10_combout ;
wire \Mux23~12_combout ;
wire \Mux23~17_combout ;
wire \Mux23~18_combout ;
wire \Mux22~7_combout ;
wire \Mux22~10_combout ;
wire \Mux22~12_combout ;
wire \Mux22~13_combout ;
wire \Mux22~17_combout ;
wire \Mux22~18_combout ;
wire \Mux21~0_combout ;
wire \Mux21~1_combout ;
wire \Mux21~2_combout ;
wire \Mux21~3_combout ;
wire \Mux21~10_combout ;
wire \Mux21~12_combout ;
wire \Mux20~7_combout ;
wire \Mux20~10_combout ;
wire \Mux20~12_combout ;
wire \Mux20~13_combout ;
wire \Mux20~14_combout ;
wire \Mux20~15_combout ;
wire \Mux20~16_combout ;
wire \Mux20~17_combout ;
wire \Mux19~2_combout ;
wire \Mux19~3_combout ;
wire \Mux19~4_combout ;
wire \Mux19~5_combout ;
wire \Mux19~6_combout ;
wire \Mux19~10_combout ;
wire \Mux19~11_combout ;
wire \Mux19~12_combout ;
wire \Mux19~13_combout ;
wire \Mux18~0_combout ;
wire \Mux18~10_combout ;
wire \Mux18~12_combout ;
wire \Mux18~13_combout ;
wire \Mux18~14_combout ;
wire \Mux18~15_combout ;
wire \Mux18~16_combout ;
wire \Mux17~2_combout ;
wire \Mux17~3_combout ;
wire \Mux17~4_combout ;
wire \Mux17~5_combout ;
wire \Mux17~6_combout ;
wire \Mux17~7_combout ;
wire \Mux17~12_combout ;
wire \Mux17~17_combout ;
wire \Mux16~4_combout ;
wire \Mux16~5_combout ;
wire \Mux16~7_combout ;
wire \Mux16~8_combout ;
wire \Mux16~12_combout ;
wire \Mux16~13_combout ;
wire \Mux16~14_combout ;
wire \Mux16~15_combout ;
wire \Mux16~16_combout ;
wire \Mux16~17_combout ;
wire \Mux15~4_combout ;
wire \Mux15~7_combout ;
wire \Mux15~8_combout ;
wire \Mux15~12_combout ;
wire \Mux15~13_combout ;
wire \Mux15~17_combout ;
wire \Mux15~18_combout ;
wire \Mux14~0_combout ;
wire \Mux14~1_combout ;
wire \Mux14~7_combout ;
wire \Mux14~10_combout ;
wire \Mux14~11_combout ;
wire \Mux14~12_combout ;
wire \Mux14~13_combout ;
wire \Mux14~17_combout ;
wire \Mux13~0_combout ;
wire \Mux13~1_combout ;
wire \Mux13~4_combout ;
wire \Mux13~10_combout ;
wire \Mux13~12_combout ;
wire \Mux13~13_combout ;
wire \Mux13~14_combout ;
wire \Mux13~15_combout ;
wire \Mux13~16_combout ;
wire \Mux13~17_combout ;
wire \Mux12~0_combout ;
wire \Mux12~2_combout ;
wire \Mux12~3_combout ;
wire \Mux12~7_combout ;
wire \Mux12~8_combout ;
wire \Mux12~12_combout ;
wire \Mux12~13_combout ;
wire \Mux12~14_combout ;
wire \Mux12~17_combout ;
wire \Mux12~18_combout ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \Mux11~2_combout ;
wire \Mux11~14_combout ;
wire \Mux11~17_combout ;
wire \Mux10~7_combout ;
wire \Mux10~8_combout ;
wire \Mux10~10_combout ;
wire \Mux10~12_combout ;
wire \Mux10~13_combout ;
wire \Mux10~17_combout ;
wire \Mux9~2_combout ;
wire \Mux9~3_combout ;
wire \Mux9~4_combout ;
wire \Mux9~5_combout ;
wire \Mux9~6_combout ;
wire \Mux9~7_combout ;
wire \Mux9~12_combout ;
wire \Mux9~14_combout ;
wire \Mux9~15_combout ;
wire \Mux9~17_combout ;
wire \Mux9~18_combout ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \Mux8~2_combout ;
wire \Mux8~4_combout ;
wire \Mux8~5_combout ;
wire \Mux8~10_combout ;
wire \Mux8~11_combout ;
wire \Mux8~14_combout ;
wire \Mux8~15_combout ;
wire \Mux8~17_combout ;
wire \Mux7~2_combout ;
wire \Mux7~3_combout ;
wire \Mux7~4_combout ;
wire \Mux7~5_combout ;
wire \Mux7~6_combout ;
wire \Mux7~7_combout ;
wire \Mux7~10_combout ;
wire \Mux7~12_combout ;
wire \Mux7~17_combout ;
wire \Mux6~2_combout ;
wire \Mux6~4_combout ;
wire \Mux6~10_combout ;
wire \Mux6~12_combout ;
wire \Mux6~13_combout ;
wire \Mux6~17_combout ;
wire \Mux6~18_combout ;
wire \Mux5~0_combout ;
wire \Mux5~1_combout ;
wire \Mux5~2_combout ;
wire \Mux5~3_combout ;
wire \Mux5~4_combout ;
wire \Mux5~7_combout ;
wire \Mux5~10_combout ;
wire \Mux5~11_combout ;
wire \Mux5~12_combout ;
wire \Mux5~17_combout ;
wire \Mux4~2_combout ;
wire \Mux4~3_combout ;
wire \Mux4~4_combout ;
wire \Mux4~5_combout ;
wire \Mux4~6_combout ;
wire \Mux4~12_combout ;
wire \Mux4~13_combout ;
wire \Mux3~7_combout ;
wire \Mux3~8_combout ;
wire \Mux3~10_combout ;
wire \Mux3~12_combout ;
wire \Mux3~13_combout ;
wire \Mux3~14_combout ;
wire \Mux3~17_combout ;
wire \Mux3~18_combout ;
wire \Mux2~2_combout ;
wire \Mux2~3_combout ;
wire \Mux2~7_combout ;
wire \Mux2~8_combout ;
wire \Mux2~10_combout ;
wire \Mux2~12_combout ;
wire \Mux2~13_combout ;
wire \Mux2~17_combout ;
wire \Mux2~18_combout ;
wire \Mux1~0_combout ;
wire \Mux1~2_combout ;
wire \Mux1~3_combout ;
wire \Mux1~4_combout ;
wire \Mux1~5_combout ;
wire \Mux1~6_combout ;
wire \Mux1~10_combout ;
wire \Mux1~11_combout ;
wire \Mux1~12_combout ;
wire \Mux1~14_combout ;
wire \Mux1~15_combout ;
wire \Mux1~17_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \Mux0~7_combout ;
wire \Mux0~12_combout ;
wire \Mux0~13_combout ;
wire \Mux0~14_combout ;
wire \Mux0~17_combout ;
wire \Mux0~18_combout ;
wire \clk~input_o ;
wire \clk~inputclkctrl_outclk ;
wire \my_rf.rsel2[4]~input_o ;
wire \my_rf.rsel2[3]~input_o ;
wire \my_rf.rsel2[0]~input_o ;
wire \my_rf.wdat[0]~input_o ;
wire \n_rst~input_o ;
wire \n_rst~inputclkctrl_outclk ;
wire \my_rf.wsel[3]~input_o ;
wire \my_rf.wsel[1]~input_o ;
wire \my_rf.wsel[0]~input_o ;
wire \Decoder0~8_combout ;
wire \my_rf.wsel[2]~input_o ;
wire \my_rf.wsel[4]~input_o ;
wire \Decoder0~25_combout ;
wire \registerArray[10][0]~q ;
wire \my_rf.WEN~input_o ;
wire \Decoder0~14_combout ;
wire \Decoder0~26_combout ;
wire \registerArray[8][0]~q ;
wire \Mux63~10_combout ;
wire \Decoder0~0_combout ;
wire \Decoder0~24_combout ;
wire \registerArray[9][0]~q ;
wire \Mux63~11_combout ;
wire \my_rf.rsel2[1]~input_o ;
wire \Decoder0~35_combout ;
wire \registerArray[14][0]~q ;
wire \Decoder0~12_combout ;
wire \Decoder0~37_combout ;
wire \registerArray[12][0]~q ;
wire \Decoder0~2_combout ;
wire \Decoder0~36_combout ;
wire \registerArray[13][0]~q ;
wire \Mux63~17_combout ;
wire \Mux63~18_combout ;
wire \Mux63~19_combout ;
wire \my_rf.rsel2[2]~input_o ;
wire \Decoder0~6_combout ;
wire \Decoder0~7_combout ;
wire \registerArray[22][0]~q ;
wire \Decoder0~11_combout ;
wire \registerArray[30][0]~q ;
wire \Mux63~3_combout ;
wire \Decoder0~13_combout ;
wire \registerArray[20][0]~q ;
wire \Decoder0~18_combout ;
wire \registerArray[28][0]~q ;
wire \Mux63~5_combout ;
wire \Mux63~6_combout ;
wire \Decoder0~5_combout ;
wire \registerArray[29][0]~q ;
wire \Decoder0~3_combout ;
wire \registerArray[21][0]~q ;
wire \Decoder0~4_combout ;
wire \registerArray[17][0]~q ;
wire \Mux63~0_combout ;
wire \Mux63~1_combout ;
wire \Mux63~9_combout ;
wire \Mux63~20_combout ;
wire \my_rf.wdat[1]~input_o ;
wire \registerArray[14][1]~q ;
wire \registerArray[13][1]~q ;
wire \Mux62~17_combout ;
wire \Mux62~18_combout ;
wire \Decoder0~28_combout ;
wire \registerArray[6][1]~q ;
wire \Decoder0~29_combout ;
wire \registerArray[5][1]~q ;
wire \Mux62~10_combout ;
wire \Mux62~11_combout ;
wire \Mux62~19_combout ;
wire \Decoder0~19_combout ;
wire \Decoder0~21_combout ;
wire \registerArray[23][1]~q ;
wire \Decoder0~23_combout ;
wire \registerArray[31][1]~q ;
wire \Mux62~8_combout ;
wire \registerArray[20][1]~q ;
wire \Decoder0~16_combout ;
wire \Decoder0~17_combout ;
wire \registerArray[16][1]~q ;
wire \Mux62~4_combout ;
wire \Decoder0~15_combout ;
wire \registerArray[24][1]~q ;
wire \registerArray[28][1]~q ;
wire \Mux62~5_combout ;
wire \Decoder0~9_combout ;
wire \registerArray[26][1]~q ;
wire \registerArray[22][1]~q ;
wire \Mux62~2_combout ;
wire \Mux62~3_combout ;
wire \Mux62~6_combout ;
wire \Mux62~9_combout ;
wire \Mux62~20_combout ;
wire \my_rf.wdat[2]~input_o ;
wire \registerArray[14][2]~q ;
wire \Decoder0~38_combout ;
wire \registerArray[15][2]~q ;
wire \Mux61~18_combout ;
wire \registerArray[6][2]~q ;
wire \registerArray[5][2]~q ;
wire \Mux61~12_combout ;
wire \Mux61~13_combout ;
wire \Decoder0~34_combout ;
wire \registerArray[2][2]~q ;
wire \Decoder0~32_combout ;
wire \registerArray[3][2]~q ;
wire \Mux61~14_combout ;
wire \Mux61~15_combout ;
wire \Mux61~16_combout ;
wire \Mux61~19_combout ;
wire \registerArray[31][2]~q ;
wire \Decoder0~20_combout ;
wire \registerArray[27][2]~q ;
wire \registerArray[23][2]~q ;
wire \Decoder0~22_combout ;
wire \registerArray[19][2]~q ;
wire \Mux61~7_combout ;
wire \Mux61~8_combout ;
wire \registerArray[29][2]~q ;
wire \registerArray[21][2]~q ;
wire \registerArray[17][2]~q ;
wire \Mux61~0_combout ;
wire \Mux61~1_combout ;
wire \Mux61~9_combout ;
wire \Mux61~20_combout ;
wire \my_rf.wdat[3]~input_o ;
wire \Decoder0~31_combout ;
wire \registerArray[7][3]~q ;
wire \registerArray[6][3]~q ;
wire \Mux60~11_combout ;
wire \registerArray[9][3]~q ;
wire \registerArray[10][3]~q ;
wire \Mux60~12_combout ;
wire \Mux60~13_combout ;
wire \registerArray[2][3]~q ;
wire \registerArray[3][3]~q ;
wire \Mux60~14_combout ;
wire \Mux60~15_combout ;
wire \Mux60~16_combout ;
wire \registerArray[14][3]~q ;
wire \registerArray[12][3]~q ;
wire \registerArray[13][3]~q ;
wire \Mux60~17_combout ;
wire \Mux60~18_combout ;
wire \Mux60~19_combout ;
wire \registerArray[29][3]~q ;
wire \registerArray[21][3]~q ;
wire \Decoder0~1_combout ;
wire \registerArray[25][3]~q ;
wire \Mux60~0_combout ;
wire \Mux60~1_combout ;
wire \registerArray[23][3]~q ;
wire \registerArray[27][3]~q ;
wire \registerArray[19][3]~q ;
wire \Mux60~7_combout ;
wire \Mux60~8_combout ;
wire \Mux60~9_combout ;
wire \Mux60~20_combout ;
wire \my_rf.wdat[4]~input_o ;
wire \registerArray[21][4]~q ;
wire \registerArray[17][4]~q ;
wire \Mux59~0_combout ;
wire \registerArray[25][4]~q ;
wire \Mux59~1_combout ;
wire \registerArray[27][4]~q ;
wire \registerArray[31][4]~q ;
wire \Mux59~8_combout ;
wire \registerArray[28][4]~q ;
wire \registerArray[20][4]~q ;
wire \registerArray[24][4]~q ;
wire \registerArray[16][4]~q ;
wire \Mux59~4_combout ;
wire \Mux59~5_combout ;
wire \Mux59~6_combout ;
wire \Mux59~9_combout ;
wire \registerArray[10][4]~q ;
wire \Mux59~10_combout ;
wire \registerArray[9][4]~q ;
wire \Mux59~11_combout ;
wire \registerArray[12][4]~q ;
wire \registerArray[13][4]~q ;
wire \Mux59~17_combout ;
wire \registerArray[14][4]~q ;
wire \registerArray[15][4]~q ;
wire \Mux59~18_combout ;
wire \Mux59~19_combout ;
wire \Mux59~20_combout ;
wire \my_rf.wdat[5]~input_o ;
wire \registerArray[2][5]~q ;
wire \Mux58~15_combout ;
wire \Mux58~16_combout ;
wire \registerArray[14][5]~q ;
wire \registerArray[12][5]~q ;
wire \registerArray[13][5]~q ;
wire \Mux58~17_combout ;
wire \Mux58~18_combout ;
wire \Mux58~19_combout ;
wire \registerArray[25][5]~q ;
wire \Mux58~0_combout ;
wire \registerArray[29][5]~q ;
wire \Mux58~1_combout ;
wire \registerArray[27][5]~q ;
wire \Mux58~7_combout ;
wire \registerArray[23][5]~q ;
wire \Mux58~8_combout ;
wire \registerArray[30][5]~q ;
wire \registerArray[26][5]~q ;
wire \registerArray[22][5]~q ;
wire \Mux58~2_combout ;
wire \Mux58~3_combout ;
wire \registerArray[20][5]~q ;
wire \registerArray[16][5]~q ;
wire \Mux58~4_combout ;
wire \registerArray[24][5]~q ;
wire \Mux58~5_combout ;
wire \Mux58~6_combout ;
wire \Mux58~9_combout ;
wire \Mux58~20_combout ;
wire \my_rf.wdat[6]~input_o ;
wire \registerArray[9][6]~q ;
wire \registerArray[10][6]~q ;
wire \registerArray[8][6]~q ;
wire \Mux57~10_combout ;
wire \Mux57~11_combout ;
wire \registerArray[6][6]~q ;
wire \registerArray[7][6]~q ;
wire \Mux57~13_combout ;
wire \Mux57~16_combout ;
wire \Mux57~19_combout ;
wire \registerArray[23][6]~q ;
wire \registerArray[19][6]~q ;
wire \Mux57~7_combout ;
wire \registerArray[27][6]~q ;
wire \Mux57~8_combout ;
wire \registerArray[20][6]~q ;
wire \registerArray[24][6]~q ;
wire \Mux57~4_combout ;
wire \Mux57~5_combout ;
wire \Mux57~6_combout ;
wire \Mux57~9_combout ;
wire \Mux57~20_combout ;
wire \my_rf.wdat[7]~input_o ;
wire \registerArray[30][7]~q ;
wire \registerArray[26][7]~q ;
wire \registerArray[22][7]~q ;
wire \Decoder0~10_combout ;
wire \registerArray[18][7]~q ;
wire \Mux56~2_combout ;
wire \Mux56~3_combout ;
wire \registerArray[20][7]~q ;
wire \registerArray[16][7]~q ;
wire \Mux56~4_combout ;
wire \registerArray[24][7]~q ;
wire \Mux56~5_combout ;
wire \Mux56~6_combout ;
wire \registerArray[23][7]~q ;
wire \registerArray[31][7]~q ;
wire \Mux56~8_combout ;
wire \Mux56~9_combout ;
wire \registerArray[3][7]~q ;
wire \Decoder0~33_combout ;
wire \registerArray[1][7]~q ;
wire \Mux56~14_combout ;
wire \registerArray[2][7]~q ;
wire \Mux56~15_combout ;
wire \Mux56~16_combout ;
wire \registerArray[6][7]~q ;
wire \registerArray[5][7]~q ;
wire \Mux56~10_combout ;
wire \Mux56~11_combout ;
wire \Mux56~19_combout ;
wire \Mux56~20_combout ;
wire \my_rf.wdat[8]~input_o ;
wire \registerArray[13][8]~q ;
wire \registerArray[12][8]~q ;
wire \Mux55~17_combout ;
wire \registerArray[14][8]~q ;
wire \registerArray[15][8]~q ;
wire \Mux55~18_combout ;
wire \registerArray[2][8]~q ;
wire \Mux55~15_combout ;
wire \registerArray[5][8]~q ;
wire \Mux55~12_combout ;
wire \registerArray[6][8]~q ;
wire \registerArray[7][8]~q ;
wire \Mux55~13_combout ;
wire \Mux55~16_combout ;
wire \registerArray[9][8]~q ;
wire \registerArray[10][8]~q ;
wire \Mux55~10_combout ;
wire \Mux55~11_combout ;
wire \Mux55~19_combout ;
wire \registerArray[21][8]~q ;
wire \registerArray[17][8]~q ;
wire \Mux55~0_combout ;
wire \registerArray[25][8]~q ;
wire \registerArray[29][8]~q ;
wire \Mux55~1_combout ;
wire \registerArray[20][8]~q ;
wire \registerArray[28][8]~q ;
wire \Mux55~5_combout ;
wire \registerArray[22][8]~q ;
wire \registerArray[30][8]~q ;
wire \Mux55~3_combout ;
wire \Mux55~6_combout ;
wire \Mux55~9_combout ;
wire \Mux55~20_combout ;
wire \my_rf.wdat[9]~input_o ;
wire \registerArray[2][9]~q ;
wire \Mux54~15_combout ;
wire \Mux54~16_combout ;
wire \registerArray[6][9]~q ;
wire \registerArray[7][9]~q ;
wire \Mux54~11_combout ;
wire \Mux54~19_combout ;
wire \registerArray[23][9]~q ;
wire \registerArray[27][9]~q ;
wire \Mux54~7_combout ;
wire \Mux54~8_combout ;
wire \registerArray[20][9]~q ;
wire \Mux54~4_combout ;
wire \registerArray[24][9]~q ;
wire \Mux54~5_combout ;
wire \registerArray[26][9]~q ;
wire \registerArray[22][9]~q ;
wire \registerArray[18][9]~q ;
wire \Mux54~2_combout ;
wire \Mux54~3_combout ;
wire \Mux54~6_combout ;
wire \registerArray[29][9]~q ;
wire \registerArray[21][9]~q ;
wire \Mux54~1_combout ;
wire \Mux54~9_combout ;
wire \Mux54~20_combout ;
wire \my_rf.wdat[10]~input_o ;
wire \registerArray[5][10]~q ;
wire \Decoder0~30_combout ;
wire \registerArray[4][10]~q ;
wire \Mux53~12_combout ;
wire \registerArray[6][10]~q ;
wire \registerArray[7][10]~q ;
wire \Mux53~13_combout ;
wire \registerArray[2][10]~q ;
wire \registerArray[3][10]~q ;
wire \registerArray[1][10]~q ;
wire \Mux53~14_combout ;
wire \Mux53~15_combout ;
wire \Mux53~16_combout ;
wire \registerArray[15][10]~q ;
wire \registerArray[14][10]~q ;
wire \registerArray[13][10]~q ;
wire \Mux53~17_combout ;
wire \Mux53~18_combout ;
wire \Mux53~19_combout ;
wire \registerArray[31][10]~q ;
wire \registerArray[27][10]~q ;
wire \registerArray[23][10]~q ;
wire \registerArray[19][10]~q ;
wire \Mux53~7_combout ;
wire \Mux53~8_combout ;
wire \registerArray[20][10]~q ;
wire \registerArray[16][10]~q ;
wire \registerArray[24][10]~q ;
wire \Mux53~4_combout ;
wire \Mux53~5_combout ;
wire \Mux53~6_combout ;
wire \Mux53~9_combout ;
wire \Mux53~20_combout ;
wire \my_rf.wdat[11]~input_o ;
wire \registerArray[26][11]~q ;
wire \registerArray[22][11]~q ;
wire \Mux52~2_combout ;
wire \Mux52~3_combout ;
wire \Mux52~6_combout ;
wire \registerArray[23][11]~q ;
wire \registerArray[19][11]~q ;
wire \registerArray[27][11]~q ;
wire \Mux52~7_combout ;
wire \Mux52~8_combout ;
wire \Mux52~9_combout ;
wire \registerArray[2][11]~q ;
wire \registerArray[3][11]~q ;
wire \registerArray[1][11]~q ;
wire \Mux52~14_combout ;
wire \Mux52~15_combout ;
wire \Decoder0~27_combout ;
wire \registerArray[11][11]~q ;
wire \registerArray[9][11]~q ;
wire \Mux52~13_combout ;
wire \Mux52~16_combout ;
wire \registerArray[5][11]~q ;
wire \registerArray[4][11]~q ;
wire \Mux52~10_combout ;
wire \registerArray[6][11]~q ;
wire \registerArray[7][11]~q ;
wire \Mux52~11_combout ;
wire \Mux52~19_combout ;
wire \Mux52~20_combout ;
wire \my_rf.wdat[12]~input_o ;
wire \registerArray[25][12]~q ;
wire \registerArray[29][12]~q ;
wire \Mux51~1_combout ;
wire \registerArray[28][12]~q ;
wire \registerArray[20][12]~q ;
wire \registerArray[24][12]~q ;
wire \registerArray[16][12]~q ;
wire \Mux51~4_combout ;
wire \Mux51~5_combout ;
wire \Mux51~6_combout ;
wire \Mux51~9_combout ;
wire \registerArray[11][12]~q ;
wire \registerArray[9][12]~q ;
wire \Mux51~11_combout ;
wire \registerArray[15][12]~q ;
wire \registerArray[14][12]~q ;
wire \registerArray[13][12]~q ;
wire \registerArray[12][12]~q ;
wire \Mux51~17_combout ;
wire \Mux51~18_combout ;
wire \registerArray[5][12]~q ;
wire \registerArray[4][12]~q ;
wire \Mux51~12_combout ;
wire \registerArray[6][12]~q ;
wire \Mux51~13_combout ;
wire \Mux51~16_combout ;
wire \Mux51~19_combout ;
wire \Mux51~20_combout ;
wire \my_rf.wdat[13]~input_o ;
wire \registerArray[4][13]~q ;
wire \registerArray[5][13]~q ;
wire \Mux50~10_combout ;
wire \registerArray[6][13]~q ;
wire \Mux50~11_combout ;
wire \registerArray[13][13]~q ;
wire \registerArray[12][13]~q ;
wire \Mux50~17_combout ;
wire \registerArray[14][13]~q ;
wire \registerArray[15][13]~q ;
wire \Mux50~18_combout ;
wire \Mux50~19_combout ;
wire \registerArray[23][13]~q ;
wire \registerArray[27][13]~q ;
wire \Mux50~7_combout ;
wire \Mux50~8_combout ;
wire \registerArray[26][13]~q ;
wire \registerArray[30][13]~q ;
wire \Mux50~3_combout ;
wire \Mux50~6_combout ;
wire \Mux50~9_combout ;
wire \Mux50~20_combout ;
wire \my_rf.wdat[14]~input_o ;
wire \registerArray[14][14]~q ;
wire \registerArray[13][14]~q ;
wire \Mux49~17_combout ;
wire \Mux49~18_combout ;
wire \registerArray[9][14]~q ;
wire \registerArray[11][14]~q ;
wire \Mux49~11_combout ;
wire \Mux49~19_combout ;
wire \registerArray[20][14]~q ;
wire \registerArray[24][14]~q ;
wire \registerArray[16][14]~q ;
wire \Mux49~4_combout ;
wire \Mux49~5_combout ;
wire \registerArray[22][14]~q ;
wire \registerArray[18][14]~q ;
wire \registerArray[26][14]~q ;
wire \Mux49~2_combout ;
wire \Mux49~3_combout ;
wire \Mux49~6_combout ;
wire \registerArray[27][14]~q ;
wire \registerArray[31][14]~q ;
wire \Mux49~8_combout ;
wire \registerArray[29][14]~q ;
wire \registerArray[21][14]~q ;
wire \Mux49~0_combout ;
wire \registerArray[25][14]~q ;
wire \Mux49~1_combout ;
wire \Mux49~9_combout ;
wire \Mux49~20_combout ;
wire \my_rf.wdat[15]~input_o ;
wire \registerArray[7][15]~q ;
wire \registerArray[6][15]~q ;
wire \registerArray[5][15]~q ;
wire \Mux48~10_combout ;
wire \Mux48~11_combout ;
wire \registerArray[3][15]~q ;
wire \registerArray[1][15]~q ;
wire \Mux48~14_combout ;
wire \registerArray[2][15]~q ;
wire \Mux48~15_combout ;
wire \Mux48~16_combout ;
wire \Mux48~19_combout ;
wire \registerArray[20][15]~q ;
wire \registerArray[16][15]~q ;
wire \Mux48~4_combout ;
wire \registerArray[24][15]~q ;
wire \Mux48~5_combout ;
wire \registerArray[30][15]~q ;
wire \registerArray[26][15]~q ;
wire \Mux48~3_combout ;
wire \Mux48~6_combout ;
wire \registerArray[27][15]~q ;
wire \registerArray[19][15]~q ;
wire \Mux48~7_combout ;
wire \registerArray[23][15]~q ;
wire \Mux48~8_combout ;
wire \registerArray[29][15]~q ;
wire \registerArray[17][15]~q ;
wire \registerArray[25][15]~q ;
wire \Mux48~0_combout ;
wire \registerArray[21][15]~q ;
wire \Mux48~1_combout ;
wire \Mux48~9_combout ;
wire \Mux48~20_combout ;
wire \my_rf.wdat[16]~input_o ;
wire \registerArray[11][16]~q ;
wire \registerArray[9][16]~q ;
wire \Mux47~11_combout ;
wire \registerArray[14][16]~q ;
wire \registerArray[15][16]~q ;
wire \Mux47~18_combout ;
wire \Mux47~19_combout ;
wire \registerArray[25][16]~q ;
wire \registerArray[21][16]~q ;
wire \registerArray[17][16]~q ;
wire \Mux47~0_combout ;
wire \Mux47~1_combout ;
wire \registerArray[22][16]~q ;
wire \registerArray[30][16]~q ;
wire \Mux47~3_combout ;
wire \Mux47~6_combout ;
wire \Mux47~9_combout ;
wire \Mux47~20_combout ;
wire \my_rf.wdat[17]~input_o ;
wire \registerArray[7][17]~q ;
wire \registerArray[6][17]~q ;
wire \Mux46~11_combout ;
wire \registerArray[14][17]~q ;
wire \registerArray[15][17]~q ;
wire \Mux46~18_combout ;
wire \Mux46~19_combout ;
wire \registerArray[21][17]~q ;
wire \registerArray[29][17]~q ;
wire \Mux46~1_combout ;
wire \registerArray[26][17]~q ;
wire \registerArray[18][17]~q ;
wire \registerArray[22][17]~q ;
wire \Mux46~2_combout ;
wire \Mux46~3_combout ;
wire \Mux46~6_combout ;
wire \Mux46~9_combout ;
wire \Mux46~20_combout ;
wire \my_rf.wdat[18]~input_o ;
wire \registerArray[6][18]~q ;
wire \registerArray[5][18]~q ;
wire \Mux45~12_combout ;
wire \Mux45~13_combout ;
wire \registerArray[2][18]~q ;
wire \registerArray[3][18]~q ;
wire \registerArray[1][18]~q ;
wire \Mux45~14_combout ;
wire \Mux45~15_combout ;
wire \Mux45~16_combout ;
wire \registerArray[13][18]~q ;
wire \registerArray[12][18]~q ;
wire \Mux45~17_combout ;
wire \registerArray[14][18]~q ;
wire \registerArray[15][18]~q ;
wire \Mux45~18_combout ;
wire \registerArray[9][18]~q ;
wire \registerArray[11][18]~q ;
wire \Mux45~11_combout ;
wire \Mux45~19_combout ;
wire \registerArray[29][18]~q ;
wire \registerArray[21][18]~q ;
wire \registerArray[17][18]~q ;
wire \Mux45~0_combout ;
wire \registerArray[25][18]~q ;
wire \Mux45~1_combout ;
wire \registerArray[20][18]~q ;
wire \registerArray[28][18]~q ;
wire \Mux45~5_combout ;
wire \registerArray[26][18]~q ;
wire \registerArray[18][18]~q ;
wire \Mux45~2_combout ;
wire \registerArray[22][18]~q ;
wire \registerArray[30][18]~q ;
wire \Mux45~3_combout ;
wire \Mux45~6_combout ;
wire \registerArray[19][18]~q ;
wire \registerArray[23][18]~q ;
wire \Mux45~7_combout ;
wire \registerArray[27][18]~q ;
wire \Mux45~8_combout ;
wire \Mux45~9_combout ;
wire \Mux45~20_combout ;
wire \my_rf.wdat[19]~input_o ;
wire \registerArray[9][19]~q ;
wire \registerArray[10][19]~q ;
wire \Mux44~12_combout ;
wire \Mux44~13_combout ;
wire \registerArray[2][19]~q ;
wire \registerArray[3][19]~q ;
wire \Mux44~14_combout ;
wire \Mux44~15_combout ;
wire \Mux44~16_combout ;
wire \registerArray[15][19]~q ;
wire \registerArray[14][19]~q ;
wire \registerArray[13][19]~q ;
wire \registerArray[12][19]~q ;
wire \Mux44~17_combout ;
wire \Mux44~18_combout ;
wire \registerArray[7][19]~q ;
wire \registerArray[6][19]~q ;
wire \registerArray[5][19]~q ;
wire \Mux44~10_combout ;
wire \Mux44~11_combout ;
wire \Mux44~19_combout ;
wire \registerArray[31][19]~q ;
wire \registerArray[23][19]~q ;
wire \Mux44~8_combout ;
wire \registerArray[21][19]~q ;
wire \registerArray[25][19]~q ;
wire \registerArray[17][19]~q ;
wire \Mux44~0_combout ;
wire \Mux44~1_combout ;
wire \Mux44~9_combout ;
wire \Mux44~20_combout ;
wire \my_rf.wdat[20]~input_o ;
wire \registerArray[9][20]~q ;
wire \registerArray[10][20]~q ;
wire \Mux43~10_combout ;
wire \Mux43~11_combout ;
wire \registerArray[5][20]~q ;
wire \registerArray[4][20]~q ;
wire \Mux43~12_combout ;
wire \registerArray[6][20]~q ;
wire \Mux43~13_combout ;
wire \Mux43~16_combout ;
wire \Mux43~19_combout ;
wire \registerArray[23][20]~q ;
wire \registerArray[19][20]~q ;
wire \Mux43~7_combout ;
wire \registerArray[27][20]~q ;
wire \registerArray[31][20]~q ;
wire \Mux43~8_combout ;
wire \registerArray[21][20]~q ;
wire \Mux43~0_combout ;
wire \registerArray[25][20]~q ;
wire \registerArray[29][20]~q ;
wire \Mux43~1_combout ;
wire \Mux43~9_combout ;
wire \Mux43~20_combout ;
wire \my_rf.wdat[21]~input_o ;
wire \registerArray[31][21]~q ;
wire \registerArray[23][21]~q ;
wire \registerArray[27][21]~q ;
wire \registerArray[19][21]~q ;
wire \Mux42~7_combout ;
wire \Mux42~8_combout ;
wire \registerArray[18][21]~q ;
wire \registerArray[22][21]~q ;
wire \Mux42~2_combout ;
wire \registerArray[26][21]~q ;
wire \Mux42~3_combout ;
wire \Mux42~6_combout ;
wire \Mux42~9_combout ;
wire \registerArray[14][21]~q ;
wire \registerArray[15][21]~q ;
wire \Mux42~18_combout ;
wire \registerArray[6][21]~q ;
wire \registerArray[5][21]~q ;
wire \registerArray[4][21]~q ;
wire \Mux42~10_combout ;
wire \Mux42~11_combout ;
wire \registerArray[9][21]~q ;
wire \registerArray[11][21]~q ;
wire \Mux42~13_combout ;
wire \registerArray[2][21]~q ;
wire \Mux42~15_combout ;
wire \Mux42~16_combout ;
wire \Mux42~19_combout ;
wire \Mux42~20_combout ;
wire \my_rf.wdat[22]~input_o ;
wire \registerArray[27][22]~q ;
wire \registerArray[23][22]~q ;
wire \Mux41~7_combout ;
wire \Mux41~8_combout ;
wire \registerArray[25][22]~q ;
wire \registerArray[21][22]~q ;
wire \Mux41~0_combout ;
wire \Mux41~1_combout ;
wire \Mux41~9_combout ;
wire \registerArray[10][22]~q ;
wire \registerArray[8][22]~q ;
wire \Mux41~10_combout ;
wire \registerArray[9][22]~q ;
wire \Mux41~11_combout ;
wire \registerArray[2][22]~q ;
wire \Mux41~15_combout ;
wire \registerArray[7][22]~q ;
wire \registerArray[6][22]~q ;
wire \registerArray[4][22]~q ;
wire \registerArray[5][22]~q ;
wire \Mux41~12_combout ;
wire \Mux41~13_combout ;
wire \Mux41~16_combout ;
wire \registerArray[14][22]~q ;
wire \registerArray[15][22]~q ;
wire \Mux41~18_combout ;
wire \Mux41~19_combout ;
wire \Mux41~20_combout ;
wire \my_rf.wdat[23]~input_o ;
wire \registerArray[31][23]~q ;
wire \registerArray[23][23]~q ;
wire \registerArray[27][23]~q ;
wire \registerArray[19][23]~q ;
wire \Mux40~7_combout ;
wire \Mux40~8_combout ;
wire \registerArray[29][23]~q ;
wire \registerArray[21][23]~q ;
wire \Mux40~1_combout ;
wire \Mux40~9_combout ;
wire \registerArray[12][23]~q ;
wire \registerArray[13][23]~q ;
wire \Mux40~17_combout ;
wire \registerArray[14][23]~q ;
wire \registerArray[15][23]~q ;
wire \Mux40~18_combout ;
wire \registerArray[7][23]~q ;
wire \registerArray[6][23]~q ;
wire \registerArray[5][23]~q ;
wire \registerArray[4][23]~q ;
wire \Mux40~10_combout ;
wire \Mux40~11_combout ;
wire \Mux40~19_combout ;
wire \Mux40~20_combout ;
wire \my_rf.wdat[24]~input_o ;
wire \registerArray[6][24]~q ;
wire \registerArray[5][24]~q ;
wire \registerArray[4][24]~q ;
wire \Mux39~12_combout ;
wire \Mux39~13_combout ;
wire \Mux39~16_combout ;
wire \registerArray[10][24]~q ;
wire \Mux39~10_combout ;
wire \registerArray[9][24]~q ;
wire \registerArray[11][24]~q ;
wire \Mux39~11_combout ;
wire \Mux39~19_combout ;
wire \registerArray[29][24]~q ;
wire \registerArray[25][24]~q ;
wire \Mux39~1_combout ;
wire \registerArray[24][24]~q ;
wire \registerArray[16][24]~q ;
wire \Mux39~4_combout ;
wire \registerArray[20][24]~q ;
wire \Mux39~5_combout ;
wire \Mux39~6_combout ;
wire \Mux39~9_combout ;
wire \Mux39~20_combout ;
wire \my_rf.wdat[25]~input_o ;
wire \registerArray[13][25]~q ;
wire \registerArray[12][25]~q ;
wire \Mux38~17_combout ;
wire \registerArray[14][25]~q ;
wire \registerArray[15][25]~q ;
wire \Mux38~18_combout ;
wire \registerArray[1][25]~q ;
wire \registerArray[3][25]~q ;
wire \Mux38~14_combout ;
wire \registerArray[2][25]~q ;
wire \Mux38~15_combout ;
wire \registerArray[8][25]~q ;
wire \registerArray[10][25]~q ;
wire \Mux38~12_combout ;
wire \registerArray[9][25]~q ;
wire \Mux38~13_combout ;
wire \Mux38~16_combout ;
wire \registerArray[5][25]~q ;
wire \Mux38~10_combout ;
wire \registerArray[6][25]~q ;
wire \Mux38~11_combout ;
wire \Mux38~19_combout ;
wire \registerArray[25][25]~q ;
wire \registerArray[17][25]~q ;
wire \Mux38~0_combout ;
wire \registerArray[29][25]~q ;
wire \Mux38~1_combout ;
wire \registerArray[26][25]~q ;
wire \registerArray[18][25]~q ;
wire \registerArray[22][25]~q ;
wire \Mux38~2_combout ;
wire \Mux38~3_combout ;
wire \Mux38~6_combout ;
wire \Mux38~9_combout ;
wire \Mux38~20_combout ;
wire \my_rf.wdat[26]~input_o ;
wire \registerArray[14][26]~q ;
wire \registerArray[13][26]~q ;
wire \Mux37~17_combout ;
wire \Mux37~18_combout ;
wire \registerArray[5][26]~q ;
wire \Mux37~12_combout ;
wire \registerArray[6][26]~q ;
wire \Mux37~13_combout ;
wire \registerArray[2][26]~q ;
wire \registerArray[3][26]~q ;
wire \registerArray[1][26]~q ;
wire \Mux37~14_combout ;
wire \Mux37~15_combout ;
wire \Mux37~16_combout ;
wire \Mux37~19_combout ;
wire \registerArray[29][26]~q ;
wire \registerArray[21][26]~q ;
wire \registerArray[17][26]~q ;
wire \Mux37~0_combout ;
wire \Mux37~1_combout ;
wire \registerArray[27][26]~q ;
wire \registerArray[31][26]~q ;
wire \Mux37~8_combout ;
wire \Mux37~9_combout ;
wire \Mux37~20_combout ;
wire \my_rf.wdat[27]~input_o ;
wire \registerArray[5][27]~q ;
wire \Mux36~10_combout ;
wire \registerArray[6][27]~q ;
wire \registerArray[7][27]~q ;
wire \Mux36~11_combout ;
wire \registerArray[10][27]~q ;
wire \Mux36~12_combout ;
wire \registerArray[9][27]~q ;
wire \Mux36~13_combout ;
wire \registerArray[2][27]~q ;
wire \registerArray[1][27]~q ;
wire \registerArray[3][27]~q ;
wire \Mux36~14_combout ;
wire \Mux36~15_combout ;
wire \Mux36~16_combout ;
wire \registerArray[15][27]~q ;
wire \registerArray[14][27]~q ;
wire \Mux36~18_combout ;
wire \Mux36~19_combout ;
wire \registerArray[29][27]~q ;
wire \registerArray[25][27]~q ;
wire \Mux36~0_combout ;
wire \Mux36~1_combout ;
wire \registerArray[24][27]~q ;
wire \registerArray[16][27]~q ;
wire \registerArray[20][27]~q ;
wire \Mux36~4_combout ;
wire \Mux36~5_combout ;
wire \Mux36~6_combout ;
wire \Mux36~9_combout ;
wire \Mux36~20_combout ;
wire \my_rf.wdat[28]~input_o ;
wire \registerArray[25][28]~q ;
wire \registerArray[29][28]~q ;
wire \Mux35~1_combout ;
wire \registerArray[28][28]~q ;
wire \registerArray[20][28]~q ;
wire \registerArray[24][28]~q ;
wire \registerArray[16][28]~q ;
wire \Mux35~4_combout ;
wire \Mux35~5_combout ;
wire \Mux35~6_combout ;
wire \Mux35~9_combout ;
wire \registerArray[14][28]~q ;
wire \registerArray[15][28]~q ;
wire \Mux35~18_combout ;
wire \registerArray[9][28]~q ;
wire \registerArray[8][28]~q ;
wire \registerArray[10][28]~q ;
wire \Mux35~10_combout ;
wire \Mux35~11_combout ;
wire \registerArray[7][28]~q ;
wire \registerArray[6][28]~q ;
wire \registerArray[5][28]~q ;
wire \registerArray[4][28]~q ;
wire \Mux35~12_combout ;
wire \Mux35~13_combout ;
wire \registerArray[2][28]~q ;
wire \registerArray[3][28]~q ;
wire \registerArray[1][28]~q ;
wire \Mux35~14_combout ;
wire \Mux35~15_combout ;
wire \Mux35~16_combout ;
wire \Mux35~19_combout ;
wire \Mux35~20_combout ;
wire \my_rf.wdat[29]~input_o ;
wire \registerArray[2][29]~q ;
wire \registerArray[1][29]~q ;
wire \registerArray[3][29]~q ;
wire \Mux34~14_combout ;
wire \Mux34~15_combout ;
wire \registerArray[11][29]~q ;
wire \registerArray[9][29]~q ;
wire \registerArray[8][29]~q ;
wire \registerArray[10][29]~q ;
wire \Mux34~12_combout ;
wire \Mux34~13_combout ;
wire \Mux34~16_combout ;
wire \registerArray[5][29]~q ;
wire \Mux34~10_combout ;
wire \registerArray[6][29]~q ;
wire \Mux34~11_combout ;
wire \registerArray[14][29]~q ;
wire \registerArray[13][29]~q ;
wire \Mux34~17_combout ;
wire \Mux34~18_combout ;
wire \Mux34~19_combout ;
wire \registerArray[31][29]~q ;
wire \registerArray[23][29]~q ;
wire \registerArray[27][29]~q ;
wire \registerArray[19][29]~q ;
wire \Mux34~7_combout ;
wire \Mux34~8_combout ;
wire \registerArray[30][29]~q ;
wire \registerArray[26][29]~q ;
wire \Mux34~3_combout ;
wire \Mux34~6_combout ;
wire \Mux34~9_combout ;
wire \Mux34~20_combout ;
wire \my_rf.wdat[30]~input_o ;
wire \registerArray[14][30]~q ;
wire \registerArray[12][30]~q ;
wire \registerArray[13][30]~q ;
wire \Mux33~17_combout ;
wire \Mux33~18_combout ;
wire \registerArray[8][30]~q ;
wire \registerArray[10][30]~q ;
wire \Mux33~10_combout ;
wire \registerArray[9][30]~q ;
wire \Mux33~11_combout ;
wire \Mux33~19_combout ;
wire \registerArray[20][30]~q ;
wire \registerArray[28][30]~q ;
wire \Mux33~5_combout ;
wire \registerArray[26][30]~q ;
wire \Mux33~2_combout ;
wire \registerArray[22][30]~q ;
wire \registerArray[30][30]~q ;
wire \Mux33~3_combout ;
wire \Mux33~6_combout ;
wire \registerArray[27][30]~q ;
wire \registerArray[23][30]~q ;
wire \Mux33~7_combout ;
wire \Mux33~8_combout ;
wire \Mux33~9_combout ;
wire \Mux33~20_combout ;
wire \my_rf.wdat[31]~input_o ;
wire \registerArray[25][31]~q ;
wire \registerArray[17][31]~q ;
wire \Mux32~0_combout ;
wire \registerArray[29][31]~q ;
wire \Mux32~1_combout ;
wire \registerArray[23][31]~q ;
wire \registerArray[31][31]~q ;
wire \Mux32~8_combout ;
wire \Mux32~9_combout ;
wire \registerArray[2][31]~q ;
wire \registerArray[3][31]~q ;
wire \Mux32~14_combout ;
wire \Mux32~15_combout ;
wire \Mux32~16_combout ;
wire \registerArray[14][31]~q ;
wire \registerArray[13][31]~q ;
wire \registerArray[12][31]~q ;
wire \Mux32~17_combout ;
wire \Mux32~18_combout ;
wire \Mux32~19_combout ;
wire \Mux32~20_combout ;
wire \my_rf.rsel1[4]~input_o ;
wire \registerArray[15][0]~q ;
wire \my_rf.rsel1[1]~input_o ;
wire \Mux31~18_combout ;
wire \my_rf.rsel1[3]~input_o ;
wire \my_rf.rsel1[0]~input_o ;
wire \registerArray[11][0]~q ;
wire \Mux31~11_combout ;
wire \Mux31~19_combout ;
wire \registerArray[31][0]~q ;
wire \registerArray[27][0]~q ;
wire \Mux31~8_combout ;
wire \my_rf.rsel1[2]~input_o ;
wire \Mux31~5_combout ;
wire \Mux31~6_combout ;
wire \Mux31~9_combout ;
wire \Mux31~20_combout ;
wire \Mux30~8_combout ;
wire \registerArray[30][1]~q ;
wire \Mux30~3_combout ;
wire \Mux30~6_combout ;
wire \Mux30~9_combout ;
wire \registerArray[7][1]~q ;
wire \registerArray[4][1]~q ;
wire \Mux30~10_combout ;
wire \Mux30~11_combout ;
wire \registerArray[15][1]~q ;
wire \registerArray[12][1]~q ;
wire \Mux30~17_combout ;
wire \Mux30~18_combout ;
wire \Mux30~19_combout ;
wire \Mux30~20_combout ;
wire \registerArray[11][2]~q ;
wire \registerArray[9][2]~q ;
wire \Mux29~11_combout ;
wire \Mux29~18_combout ;
wire \Mux29~19_combout ;
wire \registerArray[25][2]~q ;
wire \Mux29~1_combout ;
wire \registerArray[24][2]~q ;
wire \registerArray[16][2]~q ;
wire \Mux29~4_combout ;
wire \registerArray[28][2]~q ;
wire \registerArray[20][2]~q ;
wire \Mux29~5_combout ;
wire \Mux29~6_combout ;
wire \Mux29~9_combout ;
wire \Mux29~20_combout ;
wire \registerArray[31][3]~q ;
wire \Mux28~8_combout ;
wire \registerArray[30][3]~q ;
wire \registerArray[26][3]~q ;
wire \Mux28~3_combout ;
wire \registerArray[24][3]~q ;
wire \registerArray[28][3]~q ;
wire \Mux28~5_combout ;
wire \Mux28~6_combout ;
wire \Mux28~9_combout ;
wire \Mux28~15_combout ;
wire \Mux28~16_combout ;
wire \registerArray[15][3]~q ;
wire \Mux28~18_combout ;
wire \registerArray[4][3]~q ;
wire \registerArray[5][3]~q ;
wire \Mux28~10_combout ;
wire \Mux28~11_combout ;
wire \Mux28~19_combout ;
wire \Mux28~20_combout ;
wire \registerArray[8][4]~q ;
wire \Mux27~10_combout ;
wire \registerArray[11][4]~q ;
wire \Mux27~11_combout ;
wire \registerArray[3][4]~q ;
wire \registerArray[1][4]~q ;
wire \Mux27~14_combout ;
wire \registerArray[2][4]~q ;
wire \Mux27~15_combout ;
wire \Mux27~16_combout ;
wire \Mux27~19_combout ;
wire \registerArray[29][4]~q ;
wire \Mux27~0_combout ;
wire \Mux27~1_combout ;
wire \Mux27~4_combout ;
wire \Mux27~5_combout ;
wire \Mux27~6_combout ;
wire \registerArray[19][4]~q ;
wire \registerArray[23][4]~q ;
wire \Mux27~7_combout ;
wire \Mux27~8_combout ;
wire \Mux27~9_combout ;
wire \Mux27~20_combout ;
wire \registerArray[6][5]~q ;
wire \registerArray[7][5]~q ;
wire \Mux26~11_combout ;
wire \registerArray[8][5]~q ;
wire \registerArray[10][5]~q ;
wire \Mux26~12_combout ;
wire \registerArray[11][5]~q ;
wire \Mux26~13_combout ;
wire \registerArray[3][5]~q ;
wire \registerArray[1][5]~q ;
wire \Mux26~14_combout ;
wire \Mux26~15_combout ;
wire \Mux26~16_combout ;
wire \Mux26~17_combout ;
wire \registerArray[15][5]~q ;
wire \Mux26~18_combout ;
wire \Mux26~19_combout ;
wire \registerArray[17][5]~q ;
wire \Mux26~0_combout ;
wire \Mux26~1_combout ;
wire \registerArray[28][5]~q ;
wire \Mux26~4_combout ;
wire \Mux26~5_combout ;
wire \Mux26~3_combout ;
wire \Mux26~6_combout ;
wire \registerArray[31][5]~q ;
wire \registerArray[19][5]~q ;
wire \Mux26~7_combout ;
wire \Mux26~8_combout ;
wire \Mux26~9_combout ;
wire \Mux26~20_combout ;
wire \registerArray[11][6]~q ;
wire \Mux25~10_combout ;
wire \Mux25~11_combout ;
wire \registerArray[12][6]~q ;
wire \registerArray[13][6]~q ;
wire \Mux25~17_combout ;
wire \registerArray[15][6]~q ;
wire \registerArray[14][6]~q ;
wire \Mux25~18_combout ;
wire \Mux25~19_combout ;
wire \registerArray[25][6]~q ;
wire \registerArray[29][6]~q ;
wire \registerArray[17][6]~q ;
wire \registerArray[21][6]~q ;
wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \registerArray[22][6]~q ;
wire \registerArray[30][6]~q ;
wire \registerArray[18][6]~q ;
wire \registerArray[26][6]~q ;
wire \Mux25~2_combout ;
wire \Mux25~3_combout ;
wire \registerArray[16][6]~q ;
wire \Mux25~4_combout ;
wire \registerArray[28][6]~q ;
wire \Mux25~5_combout ;
wire \Mux25~6_combout ;
wire \Mux25~9_combout ;
wire \Mux25~20_combout ;
wire \registerArray[29][7]~q ;
wire \registerArray[21][7]~q ;
wire \Mux24~1_combout ;
wire \registerArray[27][7]~q ;
wire \registerArray[19][7]~q ;
wire \Mux24~7_combout ;
wire \Mux24~8_combout ;
wire \Mux24~9_combout ;
wire \registerArray[7][7]~q ;
wire \Mux24~11_combout ;
wire \Mux24~14_combout ;
wire \Mux24~15_combout ;
wire \registerArray[11][7]~q ;
wire \registerArray[9][7]~q ;
wire \Mux24~13_combout ;
wire \Mux24~16_combout ;
wire \Mux24~19_combout ;
wire \Mux24~20_combout ;
wire \registerArray[31][8]~q ;
wire \registerArray[19][8]~q ;
wire \Mux23~7_combout ;
wire \Mux23~8_combout ;
wire \Mux23~0_combout ;
wire \Mux23~1_combout ;
wire \registerArray[16][8]~q ;
wire \registerArray[24][8]~q ;
wire \Mux23~4_combout ;
wire \Mux23~5_combout ;
wire \registerArray[18][8]~q ;
wire \registerArray[26][8]~q ;
wire \Mux23~2_combout ;
wire \Mux23~3_combout ;
wire \Mux23~6_combout ;
wire \Mux23~9_combout ;
wire \registerArray[11][8]~q ;
wire \Mux23~11_combout ;
wire \Mux23~13_combout ;
wire \registerArray[3][8]~q ;
wire \registerArray[1][8]~q ;
wire \Mux23~14_combout ;
wire \Mux23~15_combout ;
wire \Mux23~16_combout ;
wire \Mux23~19_combout ;
wire \Mux23~20_combout ;
wire \registerArray[3][9]~q ;
wire \registerArray[1][9]~q ;
wire \Mux22~14_combout ;
wire \Mux22~15_combout ;
wire \Mux22~16_combout ;
wire \Mux22~11_combout ;
wire \Mux22~19_combout ;
wire \registerArray[31][9]~q ;
wire \Mux22~8_combout ;
wire \registerArray[25][9]~q ;
wire \registerArray[17][9]~q ;
wire \Mux22~0_combout ;
wire \Mux22~1_combout ;
wire \registerArray[30][9]~q ;
wire \Mux22~2_combout ;
wire \Mux22~3_combout ;
wire \registerArray[16][9]~q ;
wire \Mux22~4_combout ;
wire \registerArray[28][9]~q ;
wire \Mux22~5_combout ;
wire \Mux22~6_combout ;
wire \Mux22~9_combout ;
wire \Mux22~20_combout ;
wire \registerArray[12][10]~q ;
wire \Mux21~17_combout ;
wire \Mux21~18_combout ;
wire \Mux21~14_combout ;
wire \Mux21~15_combout ;
wire \Mux21~13_combout ;
wire \Mux21~16_combout ;
wire \registerArray[9][10]~q ;
wire \registerArray[11][10]~q ;
wire \Mux21~11_combout ;
wire \Mux21~19_combout ;
wire \Mux21~7_combout ;
wire \Mux21~8_combout ;
wire \registerArray[28][10]~q ;
wire \Mux21~4_combout ;
wire \Mux21~5_combout ;
wire \Mux21~6_combout ;
wire \Mux21~9_combout ;
wire \Mux21~20_combout ;
wire \registerArray[15][11]~q ;
wire \registerArray[14][11]~q ;
wire \Mux20~18_combout ;
wire \Mux20~11_combout ;
wire \Mux20~19_combout ;
wire \registerArray[29][11]~q ;
wire \registerArray[17][11]~q ;
wire \Mux20~0_combout ;
wire \Mux20~1_combout ;
wire \registerArray[18][11]~q ;
wire \Mux20~2_combout ;
wire \registerArray[30][11]~q ;
wire \Mux20~3_combout ;
wire \registerArray[28][11]~q ;
wire \registerArray[16][11]~q ;
wire \registerArray[20][11]~q ;
wire \Mux20~4_combout ;
wire \Mux20~5_combout ;
wire \Mux20~6_combout ;
wire \registerArray[31][11]~q ;
wire \Mux20~8_combout ;
wire \Mux20~9_combout ;
wire \Mux20~20_combout ;
wire \registerArray[17][12]~q ;
wire \Mux19~0_combout ;
wire \Mux19~1_combout ;
wire \registerArray[27][12]~q ;
wire \registerArray[31][12]~q ;
wire \registerArray[19][12]~q ;
wire \Mux19~7_combout ;
wire \Mux19~8_combout ;
wire \Mux19~9_combout ;
wire \registerArray[2][12]~q ;
wire \registerArray[1][12]~q ;
wire \registerArray[3][12]~q ;
wire \Mux19~14_combout ;
wire \Mux19~15_combout ;
wire \Mux19~16_combout ;
wire \Mux19~17_combout ;
wire \Mux19~18_combout ;
wire \Mux19~19_combout ;
wire \Mux19~20_combout ;
wire \registerArray[7][13]~q ;
wire \Mux18~11_combout ;
wire \Mux18~17_combout ;
wire \Mux18~18_combout ;
wire \Mux18~19_combout ;
wire \registerArray[28][13]~q ;
wire \registerArray[16][13]~q ;
wire \registerArray[20][13]~q ;
wire \Mux18~4_combout ;
wire \Mux18~5_combout ;
wire \registerArray[18][13]~q ;
wire \registerArray[22][13]~q ;
wire \Mux18~2_combout ;
wire \Mux18~3_combout ;
wire \Mux18~6_combout ;
wire \registerArray[29][13]~q ;
wire \registerArray[21][13]~q ;
wire \Mux18~1_combout ;
wire \registerArray[31][13]~q ;
wire \registerArray[19][13]~q ;
wire \Mux18~7_combout ;
wire \Mux18~8_combout ;
wire \Mux18~9_combout ;
wire \Mux18~20_combout ;
wire \registerArray[15][14]~q ;
wire \Mux17~18_combout ;
wire \registerArray[8][14]~q ;
wire \registerArray[10][14]~q ;
wire \Mux17~10_combout ;
wire \Mux17~11_combout ;
wire \registerArray[2][14]~q ;
wire \registerArray[3][14]~q ;
wire \registerArray[1][14]~q ;
wire \Mux17~14_combout ;
wire \Mux17~15_combout ;
wire \registerArray[6][14]~q ;
wire \registerArray[7][14]~q ;
wire \Mux17~13_combout ;
wire \Mux17~16_combout ;
wire \Mux17~19_combout ;
wire \Mux17~8_combout ;
wire \registerArray[17][14]~q ;
wire \Mux17~0_combout ;
wire \Mux17~1_combout ;
wire \Mux17~9_combout ;
wire \Mux17~20_combout ;
wire \registerArray[18][15]~q ;
wire \registerArray[22][15]~q ;
wire \Mux16~2_combout ;
wire \Mux16~3_combout ;
wire \Mux16~6_combout ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \Mux16~9_combout ;
wire \registerArray[4][15]~q ;
wire \Mux16~10_combout ;
wire \Mux16~11_combout ;
wire \registerArray[14][15]~q ;
wire \registerArray[15][15]~q ;
wire \Mux16~18_combout ;
wire \Mux16~19_combout ;
wire \Mux16~20_combout ;
wire \registerArray[29][16]~q ;
wire \Mux15~0_combout ;
wire \Mux15~1_combout ;
wire \registerArray[26][16]~q ;
wire \registerArray[18][16]~q ;
wire \Mux15~2_combout ;
wire \Mux15~3_combout ;
wire \registerArray[28][16]~q ;
wire \registerArray[20][16]~q ;
wire \Mux15~5_combout ;
wire \Mux15~6_combout ;
wire \Mux15~9_combout ;
wire \registerArray[2][16]~q ;
wire \registerArray[1][16]~q ;
wire \registerArray[3][16]~q ;
wire \Mux15~14_combout ;
wire \Mux15~15_combout ;
wire \Mux15~16_combout ;
wire \registerArray[8][16]~q ;
wire \registerArray[10][16]~q ;
wire \Mux15~10_combout ;
wire \Mux15~11_combout ;
wire \Mux15~19_combout ;
wire \Mux15~20_combout ;
wire \registerArray[1][17]~q ;
wire \Mux14~14_combout ;
wire \registerArray[2][17]~q ;
wire \Mux14~15_combout ;
wire \Mux14~16_combout ;
wire \Mux14~18_combout ;
wire \Mux14~19_combout ;
wire \registerArray[20][17]~q ;
wire \registerArray[16][17]~q ;
wire \Mux14~4_combout ;
wire \registerArray[28][17]~q ;
wire \registerArray[24][17]~q ;
wire \Mux14~5_combout ;
wire \registerArray[30][17]~q ;
wire \Mux14~2_combout ;
wire \Mux14~3_combout ;
wire \Mux14~6_combout ;
wire \registerArray[31][17]~q ;
wire \registerArray[23][17]~q ;
wire \Mux14~8_combout ;
wire \Mux14~9_combout ;
wire \Mux14~20_combout ;
wire \Mux13~11_combout ;
wire \Mux13~18_combout ;
wire \Mux13~19_combout ;
wire \Mux13~7_combout ;
wire \registerArray[31][18]~q ;
wire \Mux13~8_combout ;
wire \Mux13~2_combout ;
wire \Mux13~3_combout ;
wire \Mux13~5_combout ;
wire \Mux13~6_combout ;
wire \Mux13~9_combout ;
wire \Mux13~20_combout ;
wire \registerArray[4][19]~q ;
wire \Mux12~10_combout ;
wire \Mux12~11_combout ;
wire \Mux12~15_combout ;
wire \Mux12~16_combout ;
wire \Mux12~19_combout ;
wire \registerArray[29][19]~q ;
wire \Mux12~1_combout ;
wire \registerArray[28][19]~q ;
wire \registerArray[20][19]~q ;
wire \registerArray[16][19]~q ;
wire \Mux12~4_combout ;
wire \Mux12~5_combout ;
wire \Mux12~6_combout ;
wire \Mux12~9_combout ;
wire \Mux12~20_combout ;
wire \Mux11~7_combout ;
wire \Mux11~8_combout ;
wire \registerArray[28][20]~q ;
wire \registerArray[24][20]~q ;
wire \registerArray[16][20]~q ;
wire \Mux11~4_combout ;
wire \Mux11~5_combout ;
wire \registerArray[30][20]~q ;
wire \registerArray[22][20]~q ;
wire \Mux11~3_combout ;
wire \Mux11~6_combout ;
wire \Mux11~9_combout ;
wire \registerArray[15][20]~q ;
wire \registerArray[14][20]~q ;
wire \Mux11~18_combout ;
wire \registerArray[8][20]~q ;
wire \Mux11~10_combout ;
wire \registerArray[11][20]~q ;
wire \Mux11~11_combout ;
wire \registerArray[2][20]~q ;
wire \Mux11~15_combout ;
wire \Mux11~12_combout ;
wire \registerArray[7][20]~q ;
wire \Mux11~13_combout ;
wire \Mux11~16_combout ;
wire \Mux11~19_combout ;
wire \Mux11~20_combout ;
wire \registerArray[17][21]~q ;
wire \registerArray[25][21]~q ;
wire \Mux10~0_combout ;
wire \registerArray[29][21]~q ;
wire \Mux10~1_combout ;
wire \registerArray[20][21]~q ;
wire \registerArray[16][21]~q ;
wire \Mux10~4_combout ;
wire \registerArray[28][21]~q ;
wire \Mux10~5_combout ;
wire \Mux10~2_combout ;
wire \registerArray[30][21]~q ;
wire \Mux10~3_combout ;
wire \Mux10~6_combout ;
wire \Mux10~9_combout ;
wire \registerArray[7][21]~q ;
wire \Mux10~11_combout ;
wire \Mux10~18_combout ;
wire \registerArray[1][21]~q ;
wire \registerArray[3][21]~q ;
wire \Mux10~14_combout ;
wire \Mux10~15_combout ;
wire \Mux10~16_combout ;
wire \Mux10~19_combout ;
wire \Mux10~20_combout ;
wire \Mux9~13_combout ;
wire \Mux9~16_combout ;
wire \Mux9~10_combout ;
wire \registerArray[11][22]~q ;
wire \Mux9~11_combout ;
wire \Mux9~19_combout ;
wire \registerArray[31][22]~q ;
wire \Mux9~8_combout ;
wire \registerArray[17][22]~q ;
wire \Mux9~0_combout ;
wire \registerArray[29][22]~q ;
wire \Mux9~1_combout ;
wire \Mux9~9_combout ;
wire \Mux9~20_combout ;
wire \Mux8~18_combout ;
wire \registerArray[9][23]~q ;
wire \registerArray[11][23]~q ;
wire \registerArray[8][23]~q ;
wire \registerArray[10][23]~q ;
wire \Mux8~12_combout ;
wire \Mux8~13_combout ;
wire \Mux8~16_combout ;
wire \Mux8~19_combout ;
wire \registerArray[30][23]~q ;
wire \registerArray[26][23]~q ;
wire \Mux8~3_combout ;
wire \Mux8~6_combout ;
wire \Mux8~7_combout ;
wire \Mux8~8_combout ;
wire \Mux8~9_combout ;
wire \Mux8~20_combout ;
wire \registerArray[14][24]~q ;
wire \registerArray[15][24]~q ;
wire \Mux7~18_combout ;
wire \Mux7~11_combout ;
wire \registerArray[1][24]~q ;
wire \registerArray[3][24]~q ;
wire \Mux7~14_combout ;
wire \registerArray[2][24]~q ;
wire \Mux7~15_combout ;
wire \registerArray[7][24]~q ;
wire \Mux7~13_combout ;
wire \Mux7~16_combout ;
wire \Mux7~19_combout ;
wire \registerArray[21][24]~q ;
wire \registerArray[17][24]~q ;
wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \registerArray[27][24]~q ;
wire \registerArray[31][24]~q ;
wire \Mux7~8_combout ;
wire \Mux7~9_combout ;
wire \Mux7~20_combout ;
wire \registerArray[7][25]~q ;
wire \Mux6~11_combout ;
wire \Mux6~14_combout ;
wire \Mux6~15_combout ;
wire \Mux6~16_combout ;
wire \Mux6~19_combout ;
wire \registerArray[23][25]~q ;
wire \registerArray[31][25]~q ;
wire \registerArray[27][25]~q ;
wire \registerArray[19][25]~q ;
wire \Mux6~7_combout ;
wire \Mux6~8_combout ;
wire \Mux6~0_combout ;
wire \registerArray[21][25]~q ;
wire \Mux6~1_combout ;
wire \registerArray[30][25]~q ;
wire \Mux6~3_combout ;
wire \registerArray[28][25]~q ;
wire \registerArray[24][25]~q ;
wire \Mux6~5_combout ;
wire \Mux6~6_combout ;
wire \Mux6~9_combout ;
wire \Mux6~20_combout ;
wire \registerArray[15][26]~q ;
wire \Mux5~18_combout ;
wire \registerArray[7][26]~q ;
wire \Mux5~13_combout ;
wire \Mux5~14_combout ;
wire \Mux5~15_combout ;
wire \Mux5~16_combout ;
wire \Mux5~19_combout ;
wire \registerArray[28][26]~q ;
wire \registerArray[20][26]~q ;
wire \Mux5~5_combout ;
wire \Mux5~6_combout ;
wire \Mux5~8_combout ;
wire \Mux5~9_combout ;
wire \Mux5~20_combout ;
wire \registerArray[17][27]~q ;
wire \Mux4~0_combout ;
wire \Mux4~1_combout ;
wire \registerArray[23][27]~q ;
wire \registerArray[31][27]~q ;
wire \registerArray[19][27]~q ;
wire \registerArray[27][27]~q ;
wire \Mux4~7_combout ;
wire \Mux4~8_combout ;
wire \Mux4~9_combout ;
wire \registerArray[13][27]~q ;
wire \registerArray[12][27]~q ;
wire \Mux4~17_combout ;
wire \Mux4~18_combout ;
wire \Mux4~14_combout ;
wire \Mux4~15_combout ;
wire \Mux4~16_combout ;
wire \registerArray[4][27]~q ;
wire \Mux4~10_combout ;
wire \Mux4~11_combout ;
wire \Mux4~19_combout ;
wire \Mux4~20_combout ;
wire \registerArray[22][28]~q ;
wire \registerArray[30][28]~q ;
wire \registerArray[18][28]~q ;
wire \registerArray[26][28]~q ;
wire \Mux3~2_combout ;
wire \Mux3~3_combout ;
wire \Mux3~4_combout ;
wire \Mux3~5_combout ;
wire \Mux3~6_combout ;
wire \registerArray[17][28]~q ;
wire \registerArray[21][28]~q ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \Mux3~9_combout ;
wire \Mux3~15_combout ;
wire \Mux3~16_combout ;
wire \registerArray[11][28]~q ;
wire \Mux3~11_combout ;
wire \Mux3~19_combout ;
wire \Mux3~20_combout ;
wire \Mux2~14_combout ;
wire \Mux2~15_combout ;
wire \Mux2~16_combout ;
wire \registerArray[7][29]~q ;
wire \Mux2~11_combout ;
wire \Mux2~19_combout ;
wire \registerArray[25][29]~q ;
wire \registerArray[17][29]~q ;
wire \Mux2~0_combout ;
wire \registerArray[29][29]~q ;
wire \registerArray[21][29]~q ;
wire \Mux2~1_combout ;
wire \registerArray[16][29]~q ;
wire \Mux2~4_combout ;
wire \registerArray[28][29]~q ;
wire \registerArray[24][29]~q ;
wire \Mux2~5_combout ;
wire \Mux2~6_combout ;
wire \Mux2~9_combout ;
wire \Mux2~20_combout ;
wire \registerArray[15][30]~q ;
wire \Mux1~18_combout ;
wire \registerArray[6][30]~q ;
wire \registerArray[7][30]~q ;
wire \Mux1~13_combout ;
wire \Mux1~16_combout ;
wire \Mux1~19_combout ;
wire \registerArray[29][30]~q ;
wire \registerArray[25][30]~q ;
wire \Mux1~1_combout ;
wire \registerArray[31][30]~q ;
wire \registerArray[19][30]~q ;
wire \Mux1~7_combout ;
wire \Mux1~8_combout ;
wire \Mux1~9_combout ;
wire \Mux1~20_combout ;
wire \registerArray[20][31]~q ;
wire \registerArray[16][31]~q ;
wire \Mux0~4_combout ;
wire \registerArray[28][31]~q ;
wire \registerArray[24][31]~q ;
wire \Mux0~5_combout ;
wire \Mux0~6_combout ;
wire \Mux0~8_combout ;
wire \Mux0~9_combout ;
wire \Mux0~15_combout ;
wire \Mux0~16_combout ;
wire \registerArray[4][31]~q ;
wire \registerArray[5][31]~q ;
wire \Mux0~10_combout ;
wire \registerArray[7][31]~q ;
wire \registerArray[6][31]~q ;
wire \Mux0~11_combout ;
wire \Mux0~19_combout ;
wire \Mux0~20_combout ;


// Location: FF_X56_Y0_N24
dffeas \registerArray[25][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[0]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][0] .is_wysiwyg = "true";
defparam \registerArray[25][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y38_N1
dffeas \registerArray[26][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][0] .is_wysiwyg = "true";
defparam \registerArray[26][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y38_N19
dffeas \registerArray[18][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][0] .is_wysiwyg = "true";
defparam \registerArray[18][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N0
cycloneive_lcell_comb \Mux63~2 (
// Equation(s):
// \Mux63~2_combout  = (\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o ) # ((\registerArray[26][0]~q )))) # (!\my_rf.rsel2[3]~input_o  & (!\my_rf.rsel2[2]~input_o  & ((\registerArray[18][0]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[26][0]~q ),
	.datad(\registerArray[18][0]~q ),
	.cin(gnd),
	.combout(\Mux63~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~2 .lut_mask = 16'hB9A8;
defparam \Mux63~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y31_N25
dffeas \registerArray[24][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][0] .is_wysiwyg = "true";
defparam \registerArray[24][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y31_N27
dffeas \registerArray[16][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][0] .is_wysiwyg = "true";
defparam \registerArray[16][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N24
cycloneive_lcell_comb \Mux63~4 (
// Equation(s):
// \Mux63~4_combout  = (\my_rf.rsel2[3]~input_o  & (((\registerArray[24][0]~q ) # (\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[16][0]~q  & ((!\my_rf.rsel2[2]~input_o ))))

	.dataa(\registerArray[16][0]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][0]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux63~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~4 .lut_mask = 16'hCCE2;
defparam \Mux63~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y28_N1
dffeas \registerArray[23][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][0] .is_wysiwyg = "true";
defparam \registerArray[23][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N3
dffeas \registerArray[19][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][0] .is_wysiwyg = "true";
defparam \registerArray[19][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N0
cycloneive_lcell_comb \Mux63~7 (
// Equation(s):
// \Mux63~7_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[23][0]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[19][0]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[23][0]~q ),
	.datad(\registerArray[19][0]~q ),
	.cin(gnd),
	.combout(\Mux63~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~7 .lut_mask = 16'hB9A8;
defparam \Mux63~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N16
cycloneive_lcell_comb \Mux63~8 (
// Equation(s):
// \Mux63~8_combout  = (\Mux63~7_combout  & ((\registerArray[31][0]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux63~7_combout  & (((\registerArray[27][0]~q  & \my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[31][0]~q ),
	.datab(\Mux63~7_combout ),
	.datac(\registerArray[27][0]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux63~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~8 .lut_mask = 16'hB8CC;
defparam \Mux63~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y29_N9
dffeas \registerArray[6][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][0] .is_wysiwyg = "true";
defparam \registerArray[6][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y29_N9
dffeas \registerArray[5][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][0] .is_wysiwyg = "true";
defparam \registerArray[5][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y29_N11
dffeas \registerArray[4][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][0] .is_wysiwyg = "true";
defparam \registerArray[4][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N8
cycloneive_lcell_comb \Mux63~12 (
// Equation(s):
// \Mux63~12_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[5][0]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][0]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[4][0]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][0]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux63~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~12 .lut_mask = 16'hCCE2;
defparam \Mux63~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y29_N3
dffeas \registerArray[7][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][0] .is_wysiwyg = "true";
defparam \registerArray[7][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N8
cycloneive_lcell_comb \Mux63~13 (
// Equation(s):
// \Mux63~13_combout  = (\Mux63~12_combout  & (((\registerArray[7][0]~q )) # (!\my_rf.rsel2[1]~input_o ))) # (!\Mux63~12_combout  & (\my_rf.rsel2[1]~input_o  & (\registerArray[6][0]~q )))

	.dataa(\Mux63~12_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[6][0]~q ),
	.datad(\registerArray[7][0]~q ),
	.cin(gnd),
	.combout(\Mux63~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~13 .lut_mask = 16'hEA62;
defparam \Mux63~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y31_N17
dffeas \registerArray[3][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][0] .is_wysiwyg = "true";
defparam \registerArray[3][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N3
dffeas \registerArray[1][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][0] .is_wysiwyg = "true";
defparam \registerArray[1][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N16
cycloneive_lcell_comb \Mux63~14 (
// Equation(s):
// \Mux63~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][0]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][0]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][0]~q ),
	.datad(\registerArray[1][0]~q ),
	.cin(gnd),
	.combout(\Mux63~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~14 .lut_mask = 16'hC480;
defparam \Mux63~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N25
dffeas \registerArray[2][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][0] .is_wysiwyg = "true";
defparam \registerArray[2][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N24
cycloneive_lcell_comb \Mux63~15 (
// Equation(s):
// \Mux63~15_combout  = (\Mux63~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][0]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][0]~q ),
	.datad(\Mux63~14_combout ),
	.cin(gnd),
	.combout(\Mux63~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~15 .lut_mask = 16'hFF20;
defparam \Mux63~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N26
cycloneive_lcell_comb \Mux63~16 (
// Equation(s):
// \Mux63~16_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux63~13_combout ) # ((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (((!\my_rf.rsel2[3]~input_o  & \Mux63~15_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux63~13_combout ),
	.datac(\my_rf.rsel2[3]~input_o ),
	.datad(\Mux63~15_combout ),
	.cin(gnd),
	.combout(\Mux63~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~16 .lut_mask = 16'hADA8;
defparam \Mux63~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y0_N24
dffeas \registerArray[21][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[1]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][1] .is_wysiwyg = "true";
defparam \registerArray[21][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N17
dffeas \registerArray[25][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][1] .is_wysiwyg = "true";
defparam \registerArray[25][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N3
dffeas \registerArray[17][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][1] .is_wysiwyg = "true";
defparam \registerArray[17][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N16
cycloneive_lcell_comb \Mux62~0 (
// Equation(s):
// \Mux62~0_combout  = (\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o ) # ((\registerArray[25][1]~q )))) # (!\my_rf.rsel2[3]~input_o  & (!\my_rf.rsel2[2]~input_o  & ((\registerArray[17][1]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[25][1]~q ),
	.datad(\registerArray[17][1]~q ),
	.cin(gnd),
	.combout(\Mux62~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~0 .lut_mask = 16'hB9A8;
defparam \Mux62~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N25
dffeas \registerArray[29][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][1] .is_wysiwyg = "true";
defparam \registerArray[29][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N2
cycloneive_lcell_comb \Mux62~1 (
// Equation(s):
// \Mux62~1_combout  = (\Mux62~0_combout  & ((\registerArray[29][1]~q ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux62~0_combout  & (((\registerArray[21][1]~q  & \my_rf.rsel2[2]~input_o ))))

	.dataa(\Mux62~0_combout ),
	.datab(\registerArray[29][1]~q ),
	.datac(\registerArray[21][1]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux62~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~1 .lut_mask = 16'hD8AA;
defparam \Mux62~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N27
dffeas \registerArray[18][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][1] .is_wysiwyg = "true";
defparam \registerArray[18][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y28_N21
dffeas \registerArray[27][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][1] .is_wysiwyg = "true";
defparam \registerArray[27][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N7
dffeas \registerArray[19][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][1] .is_wysiwyg = "true";
defparam \registerArray[19][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N20
cycloneive_lcell_comb \Mux62~7 (
// Equation(s):
// \Mux62~7_combout  = (\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o ) # ((\registerArray[27][1]~q )))) # (!\my_rf.rsel2[3]~input_o  & (!\my_rf.rsel2[2]~input_o  & ((\registerArray[19][1]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[27][1]~q ),
	.datad(\registerArray[19][1]~q ),
	.cin(gnd),
	.combout(\Mux62~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~7 .lut_mask = 16'hB9A8;
defparam \Mux62~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y31_N13
dffeas \registerArray[9][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][1] .is_wysiwyg = "true";
defparam \registerArray[9][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y31_N13
dffeas \registerArray[10][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][1] .is_wysiwyg = "true";
defparam \registerArray[10][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y31_N7
dffeas \registerArray[8][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][1] .is_wysiwyg = "true";
defparam \registerArray[8][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N12
cycloneive_lcell_comb \Mux62~12 (
// Equation(s):
// \Mux62~12_combout  = (\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o ) # ((\registerArray[10][1]~q )))) # (!\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & ((\registerArray[8][1]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[10][1]~q ),
	.datad(\registerArray[8][1]~q ),
	.cin(gnd),
	.combout(\Mux62~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~12 .lut_mask = 16'hB9A8;
defparam \Mux62~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y31_N31
dffeas \registerArray[11][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][1] .is_wysiwyg = "true";
defparam \registerArray[11][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N12
cycloneive_lcell_comb \Mux62~13 (
// Equation(s):
// \Mux62~13_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux62~12_combout  & ((\registerArray[11][1]~q ))) # (!\Mux62~12_combout  & (\registerArray[9][1]~q )))) # (!\my_rf.rsel2[0]~input_o  & (\Mux62~12_combout ))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\Mux62~12_combout ),
	.datac(\registerArray[9][1]~q ),
	.datad(\registerArray[11][1]~q ),
	.cin(gnd),
	.combout(\Mux62~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~13 .lut_mask = 16'hEC64;
defparam \Mux62~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y31_N29
dffeas \registerArray[3][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][1] .is_wysiwyg = "true";
defparam \registerArray[3][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N7
dffeas \registerArray[1][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][1] .is_wysiwyg = "true";
defparam \registerArray[1][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N28
cycloneive_lcell_comb \Mux62~14 (
// Equation(s):
// \Mux62~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][1]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][1]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][1]~q ),
	.datad(\registerArray[1][1]~q ),
	.cin(gnd),
	.combout(\Mux62~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~14 .lut_mask = 16'hC480;
defparam \Mux62~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N9
dffeas \registerArray[2][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][1] .is_wysiwyg = "true";
defparam \registerArray[2][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N8
cycloneive_lcell_comb \Mux62~15 (
// Equation(s):
// \Mux62~15_combout  = (\Mux62~14_combout ) # ((!\my_rf.rsel2[0]~input_o  & (\my_rf.rsel2[1]~input_o  & \registerArray[2][1]~q )))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[2][1]~q ),
	.datad(\Mux62~14_combout ),
	.cin(gnd),
	.combout(\Mux62~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~15 .lut_mask = 16'hFF40;
defparam \Mux62~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N12
cycloneive_lcell_comb \Mux62~16 (
// Equation(s):
// \Mux62~16_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\Mux62~13_combout )) # (!\my_rf.rsel2[3]~input_o  & ((\Mux62~15_combout )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux62~13_combout ),
	.datad(\Mux62~15_combout ),
	.cin(gnd),
	.combout(\Mux62~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~16 .lut_mask = 16'hD9C8;
defparam \Mux62~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N29
dffeas \registerArray[22][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][2] .is_wysiwyg = "true";
defparam \registerArray[22][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N1
dffeas \registerArray[26][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][2] .is_wysiwyg = "true";
defparam \registerArray[26][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y38_N5
dffeas \registerArray[18][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][2] .is_wysiwyg = "true";
defparam \registerArray[18][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N0
cycloneive_lcell_comb \Mux61~2 (
// Equation(s):
// \Mux61~2_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & ((\registerArray[26][2]~q ))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[18][2]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[18][2]~q ),
	.datac(\registerArray[26][2]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux61~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~2 .lut_mask = 16'hFA44;
defparam \Mux61~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N3
dffeas \registerArray[30][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][2] .is_wysiwyg = "true";
defparam \registerArray[30][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N28
cycloneive_lcell_comb \Mux61~3 (
// Equation(s):
// \Mux61~3_combout  = (\Mux61~2_combout  & ((\registerArray[30][2]~q ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux61~2_combout  & (((\registerArray[22][2]~q  & \my_rf.rsel2[2]~input_o ))))

	.dataa(\registerArray[30][2]~q ),
	.datab(\Mux61~2_combout ),
	.datac(\registerArray[22][2]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux61~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~3 .lut_mask = 16'hB8CC;
defparam \Mux61~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N4
cycloneive_lcell_comb \Mux61~4 (
// Equation(s):
// \Mux61~4_combout  = (\my_rf.rsel2[3]~input_o  & (((\registerArray[24][2]~q ) # (\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[16][2]~q  & ((!\my_rf.rsel2[2]~input_o ))))

	.dataa(\registerArray[16][2]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][2]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux61~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~4 .lut_mask = 16'hCCE2;
defparam \Mux61~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N2
cycloneive_lcell_comb \Mux61~5 (
// Equation(s):
// \Mux61~5_combout  = (\Mux61~4_combout  & ((\registerArray[28][2]~q ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux61~4_combout  & (((\registerArray[20][2]~q  & \my_rf.rsel2[2]~input_o ))))

	.dataa(\Mux61~4_combout ),
	.datab(\registerArray[28][2]~q ),
	.datac(\registerArray[20][2]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux61~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~5 .lut_mask = 16'hD8AA;
defparam \Mux61~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N2
cycloneive_lcell_comb \Mux61~6 (
// Equation(s):
// \Mux61~6_combout  = (\my_rf.rsel2[0]~input_o  & (((\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\Mux61~3_combout )) # (!\my_rf.rsel2[1]~input_o  & ((\Mux61~5_combout )))))

	.dataa(\Mux61~3_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\my_rf.rsel2[1]~input_o ),
	.datad(\Mux61~5_combout ),
	.cin(gnd),
	.combout(\Mux61~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~6 .lut_mask = 16'hE3E0;
defparam \Mux61~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y31_N25
dffeas \registerArray[10][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][2] .is_wysiwyg = "true";
defparam \registerArray[10][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y31_N3
dffeas \registerArray[8][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][2] .is_wysiwyg = "true";
defparam \registerArray[8][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N24
cycloneive_lcell_comb \Mux61~10 (
// Equation(s):
// \Mux61~10_combout  = (\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o ) # ((\registerArray[10][2]~q )))) # (!\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & ((\registerArray[8][2]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[10][2]~q ),
	.datad(\registerArray[8][2]~q ),
	.cin(gnd),
	.combout(\Mux61~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~10 .lut_mask = 16'hB9A8;
defparam \Mux61~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N24
cycloneive_lcell_comb \Mux61~11 (
// Equation(s):
// \Mux61~11_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux61~10_combout  & (\registerArray[11][2]~q )) # (!\Mux61~10_combout  & ((\registerArray[9][2]~q ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux61~10_combout ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\registerArray[11][2]~q ),
	.datac(\registerArray[9][2]~q ),
	.datad(\Mux61~10_combout ),
	.cin(gnd),
	.combout(\Mux61~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~11 .lut_mask = 16'hDDA0;
defparam \Mux61~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y29_N19
dffeas \registerArray[4][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][2] .is_wysiwyg = "true";
defparam \registerArray[4][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y29_N27
dffeas \registerArray[7][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][2] .is_wysiwyg = "true";
defparam \registerArray[7][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N27
dffeas \registerArray[1][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][2] .is_wysiwyg = "true";
defparam \registerArray[1][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N17
dffeas \registerArray[13][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][2] .is_wysiwyg = "true";
defparam \registerArray[13][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N27
dffeas \registerArray[12][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][2] .is_wysiwyg = "true";
defparam \registerArray[12][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N16
cycloneive_lcell_comb \Mux61~17 (
// Equation(s):
// \Mux61~17_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & ((\registerArray[13][2]~q ))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[12][2]~q ))))

	.dataa(\registerArray[12][2]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[13][2]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux61~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~17 .lut_mask = 16'hFC22;
defparam \Mux61~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N7
dffeas \registerArray[17][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][3] .is_wysiwyg = "true";
defparam \registerArray[17][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y36_N13
dffeas \registerArray[22][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][3] .is_wysiwyg = "true";
defparam \registerArray[22][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y36_N15
dffeas \registerArray[18][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][3] .is_wysiwyg = "true";
defparam \registerArray[18][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N12
cycloneive_lcell_comb \Mux60~2 (
// Equation(s):
// \Mux60~2_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & ((\registerArray[22][3]~q ))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[18][3]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[18][3]~q ),
	.datac(\registerArray[22][3]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux60~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~2 .lut_mask = 16'hFA44;
defparam \Mux60~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N12
cycloneive_lcell_comb \Mux60~3 (
// Equation(s):
// \Mux60~3_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux60~2_combout  & (\registerArray[30][3]~q )) # (!\Mux60~2_combout  & ((\registerArray[26][3]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux60~2_combout ))))

	.dataa(\registerArray[30][3]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[26][3]~q ),
	.datad(\Mux60~2_combout ),
	.cin(gnd),
	.combout(\Mux60~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~3 .lut_mask = 16'hBBC0;
defparam \Mux60~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y36_N21
dffeas \registerArray[20][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][3] .is_wysiwyg = "true";
defparam \registerArray[20][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N31
dffeas \registerArray[16][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][3] .is_wysiwyg = "true";
defparam \registerArray[16][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N20
cycloneive_lcell_comb \Mux60~4 (
// Equation(s):
// \Mux60~4_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[20][3]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[16][3]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[16][3]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[20][3]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux60~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~4 .lut_mask = 16'hCCE2;
defparam \Mux60~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N30
cycloneive_lcell_comb \Mux60~5 (
// Equation(s):
// \Mux60~5_combout  = (\Mux60~4_combout  & ((\registerArray[28][3]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux60~4_combout  & (((\registerArray[24][3]~q  & \my_rf.rsel2[3]~input_o ))))

	.dataa(\Mux60~4_combout ),
	.datab(\registerArray[28][3]~q ),
	.datac(\registerArray[24][3]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux60~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~5 .lut_mask = 16'hD8AA;
defparam \Mux60~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N22
cycloneive_lcell_comb \Mux60~6 (
// Equation(s):
// \Mux60~6_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux60~3_combout ) # ((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux60~5_combout  & !\my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux60~3_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\Mux60~5_combout ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux60~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~6 .lut_mask = 16'hCCB8;
defparam \Mux60~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N12
cycloneive_lcell_comb \Mux60~10 (
// Equation(s):
// \Mux60~10_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[5][3]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][3]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[4][3]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][3]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux60~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~10 .lut_mask = 16'hCCE2;
defparam \Mux60~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y31_N31
dffeas \registerArray[8][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][3] .is_wysiwyg = "true";
defparam \registerArray[8][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y31_N23
dffeas \registerArray[11][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][3] .is_wysiwyg = "true";
defparam \registerArray[11][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N23
dffeas \registerArray[1][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][3] .is_wysiwyg = "true";
defparam \registerArray[1][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y36_N1
dffeas \registerArray[22][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][4] .is_wysiwyg = "true";
defparam \registerArray[22][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y32_N17
dffeas \registerArray[26][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][4] .is_wysiwyg = "true";
defparam \registerArray[26][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y36_N11
dffeas \registerArray[18][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][4] .is_wysiwyg = "true";
defparam \registerArray[18][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N16
cycloneive_lcell_comb \Mux59~2 (
// Equation(s):
// \Mux59~2_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[26][4]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[18][4]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[26][4]~q ),
	.datad(\registerArray[18][4]~q ),
	.cin(gnd),
	.combout(\Mux59~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~2 .lut_mask = 16'hD9C8;
defparam \Mux59~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y32_N11
dffeas \registerArray[30][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][4] .is_wysiwyg = "true";
defparam \registerArray[30][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N0
cycloneive_lcell_comb \Mux59~3 (
// Equation(s):
// \Mux59~3_combout  = (\Mux59~2_combout  & ((\registerArray[30][4]~q ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux59~2_combout  & (((\registerArray[22][4]~q  & \my_rf.rsel2[2]~input_o ))))

	.dataa(\registerArray[30][4]~q ),
	.datab(\Mux59~2_combout ),
	.datac(\registerArray[22][4]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux59~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~3 .lut_mask = 16'hB8CC;
defparam \Mux59~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N16
cycloneive_lcell_comb \Mux59~7 (
// Equation(s):
// \Mux59~7_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & ((\registerArray[23][4]~q ))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[19][4]~q ))))

	.dataa(\registerArray[19][4]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[23][4]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux59~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~7 .lut_mask = 16'hFC22;
defparam \Mux59~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y29_N17
dffeas \registerArray[6][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][4] .is_wysiwyg = "true";
defparam \registerArray[6][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y29_N17
dffeas \registerArray[5][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][4] .is_wysiwyg = "true";
defparam \registerArray[5][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y29_N27
dffeas \registerArray[4][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][4] .is_wysiwyg = "true";
defparam \registerArray[4][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N16
cycloneive_lcell_comb \Mux59~12 (
// Equation(s):
// \Mux59~12_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[5][4]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][4]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[4][4]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][4]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux59~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~12 .lut_mask = 16'hCCE2;
defparam \Mux59~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y29_N19
dffeas \registerArray[7][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][4] .is_wysiwyg = "true";
defparam \registerArray[7][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N16
cycloneive_lcell_comb \Mux59~13 (
// Equation(s):
// \Mux59~13_combout  = (\Mux59~12_combout  & (((\registerArray[7][4]~q )) # (!\my_rf.rsel2[1]~input_o ))) # (!\Mux59~12_combout  & (\my_rf.rsel2[1]~input_o  & (\registerArray[6][4]~q )))

	.dataa(\Mux59~12_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[6][4]~q ),
	.datad(\registerArray[7][4]~q ),
	.cin(gnd),
	.combout(\Mux59~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~13 .lut_mask = 16'hEA62;
defparam \Mux59~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N8
cycloneive_lcell_comb \Mux59~14 (
// Equation(s):
// \Mux59~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][4]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][4]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][4]~q ),
	.datad(\registerArray[1][4]~q ),
	.cin(gnd),
	.combout(\Mux59~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~14 .lut_mask = 16'hC480;
defparam \Mux59~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N22
cycloneive_lcell_comb \Mux59~15 (
// Equation(s):
// \Mux59~15_combout  = (\Mux59~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][4]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][4]~q ),
	.datad(\Mux59~14_combout ),
	.cin(gnd),
	.combout(\Mux59~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~15 .lut_mask = 16'hFF20;
defparam \Mux59~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N10
cycloneive_lcell_comb \Mux59~16 (
// Equation(s):
// \Mux59~16_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\Mux59~13_combout )) # (!\my_rf.rsel2[2]~input_o  & ((\Mux59~15_combout )))))

	.dataa(\Mux59~13_combout ),
	.datab(\Mux59~15_combout ),
	.datac(\my_rf.rsel2[3]~input_o ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux59~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~16 .lut_mask = 16'hFA0C;
defparam \Mux59~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y0_N3
dffeas \registerArray[21][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[5]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][5] .is_wysiwyg = "true";
defparam \registerArray[21][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y36_N23
dffeas \registerArray[18][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][5] .is_wysiwyg = "true";
defparam \registerArray[18][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y29_N5
dffeas \registerArray[5][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][5] .is_wysiwyg = "true";
defparam \registerArray[5][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y29_N7
dffeas \registerArray[4][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][5] .is_wysiwyg = "true";
defparam \registerArray[4][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N4
cycloneive_lcell_comb \Mux58~10 (
// Equation(s):
// \Mux58~10_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[5][5]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][5]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[4][5]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][5]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux58~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~10 .lut_mask = 16'hCCE2;
defparam \Mux58~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N4
cycloneive_lcell_comb \Mux58~11 (
// Equation(s):
// \Mux58~11_combout  = (\Mux58~10_combout  & ((\registerArray[7][5]~q ) # ((!\my_rf.rsel2[1]~input_o )))) # (!\Mux58~10_combout  & (((\registerArray[6][5]~q  & \my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[7][5]~q ),
	.datab(\Mux58~10_combout ),
	.datac(\registerArray[6][5]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux58~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~11 .lut_mask = 16'hB8CC;
defparam \Mux58~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y31_N13
dffeas \registerArray[9][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][5] .is_wysiwyg = "true";
defparam \registerArray[9][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N28
cycloneive_lcell_comb \Mux58~12 (
// Equation(s):
// \Mux58~12_combout  = (\my_rf.rsel2[0]~input_o  & (((\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[10][5]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[8][5]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\registerArray[8][5]~q ),
	.datac(\registerArray[10][5]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux58~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~12 .lut_mask = 16'hFA44;
defparam \Mux58~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N12
cycloneive_lcell_comb \Mux58~13 (
// Equation(s):
// \Mux58~13_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux58~12_combout  & (\registerArray[11][5]~q )) # (!\Mux58~12_combout  & ((\registerArray[9][5]~q ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux58~12_combout ))))

	.dataa(\registerArray[11][5]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[9][5]~q ),
	.datad(\Mux58~12_combout ),
	.cin(gnd),
	.combout(\Mux58~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~13 .lut_mask = 16'hBBC0;
defparam \Mux58~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N4
cycloneive_lcell_comb \Mux58~14 (
// Equation(s):
// \Mux58~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[3][5]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[1][5]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[1][5]~q ),
	.datac(\registerArray[3][5]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux58~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~14 .lut_mask = 16'hE400;
defparam \Mux58~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N28
cycloneive_lcell_comb \Mux57~0 (
// Equation(s):
// \Mux57~0_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[21][6]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[17][6]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[17][6]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[21][6]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux57~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~0 .lut_mask = 16'hCCE2;
defparam \Mux57~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N10
cycloneive_lcell_comb \Mux57~1 (
// Equation(s):
// \Mux57~1_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux57~0_combout  & (\registerArray[29][6]~q )) # (!\Mux57~0_combout  & ((\registerArray[25][6]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (\Mux57~0_combout ))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux57~0_combout ),
	.datac(\registerArray[29][6]~q ),
	.datad(\registerArray[25][6]~q ),
	.cin(gnd),
	.combout(\Mux57~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~1 .lut_mask = 16'hE6C4;
defparam \Mux57~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N8
cycloneive_lcell_comb \Mux57~2 (
// Equation(s):
// \Mux57~2_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[26][6]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[18][6]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[26][6]~q ),
	.datad(\registerArray[18][6]~q ),
	.cin(gnd),
	.combout(\Mux57~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~2 .lut_mask = 16'hD9C8;
defparam \Mux57~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N24
cycloneive_lcell_comb \Mux57~3 (
// Equation(s):
// \Mux57~3_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux57~2_combout  & (\registerArray[30][6]~q )) # (!\Mux57~2_combout  & ((\registerArray[22][6]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux57~2_combout ))))

	.dataa(\registerArray[30][6]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][6]~q ),
	.datad(\Mux57~2_combout ),
	.cin(gnd),
	.combout(\Mux57~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~3 .lut_mask = 16'hBBC0;
defparam \Mux57~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y32_N27
dffeas \registerArray[31][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][6] .is_wysiwyg = "true";
defparam \registerArray[31][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y29_N25
dffeas \registerArray[5][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][6] .is_wysiwyg = "true";
defparam \registerArray[5][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y29_N3
dffeas \registerArray[4][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][6] .is_wysiwyg = "true";
defparam \registerArray[4][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N24
cycloneive_lcell_comb \Mux57~12 (
// Equation(s):
// \Mux57~12_combout  = (\my_rf.rsel2[1]~input_o  & (\my_rf.rsel2[0]~input_o )) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & (\registerArray[5][6]~q )) # (!\my_rf.rsel2[0]~input_o  & ((\registerArray[4][6]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][6]~q ),
	.datad(\registerArray[4][6]~q ),
	.cin(gnd),
	.combout(\Mux57~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~12 .lut_mask = 16'hD9C8;
defparam \Mux57~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y31_N1
dffeas \registerArray[3][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][6] .is_wysiwyg = "true";
defparam \registerArray[3][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N19
dffeas \registerArray[1][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][6] .is_wysiwyg = "true";
defparam \registerArray[1][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N0
cycloneive_lcell_comb \Mux57~14 (
// Equation(s):
// \Mux57~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][6]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][6]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][6]~q ),
	.datad(\registerArray[1][6]~q ),
	.cin(gnd),
	.combout(\Mux57~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~14 .lut_mask = 16'hC480;
defparam \Mux57~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N19
dffeas \registerArray[2][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][6] .is_wysiwyg = "true";
defparam \registerArray[2][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N18
cycloneive_lcell_comb \Mux57~15 (
// Equation(s):
// \Mux57~15_combout  = (\Mux57~14_combout ) # ((!\my_rf.rsel2[0]~input_o  & (\registerArray[2][6]~q  & \my_rf.rsel2[1]~input_o )))

	.dataa(\Mux57~14_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][6]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux57~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~15 .lut_mask = 16'hBAAA;
defparam \Mux57~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N24
cycloneive_lcell_comb \Mux57~17 (
// Equation(s):
// \Mux57~17_combout  = (\my_rf.rsel2[1]~input_o  & (\my_rf.rsel2[0]~input_o )) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & (\registerArray[13][6]~q )) # (!\my_rf.rsel2[0]~input_o  & ((\registerArray[12][6]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[13][6]~q ),
	.datad(\registerArray[12][6]~q ),
	.cin(gnd),
	.combout(\Mux57~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~17 .lut_mask = 16'hD9C8;
defparam \Mux57~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N12
cycloneive_lcell_comb \Mux57~18 (
// Equation(s):
// \Mux57~18_combout  = (\Mux57~17_combout  & (((\registerArray[15][6]~q )) # (!\my_rf.rsel2[1]~input_o ))) # (!\Mux57~17_combout  & (\my_rf.rsel2[1]~input_o  & (\registerArray[14][6]~q )))

	.dataa(\Mux57~17_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][6]~q ),
	.datad(\registerArray[15][6]~q ),
	.cin(gnd),
	.combout(\Mux57~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~18 .lut_mask = 16'hEA62;
defparam \Mux57~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N31
dffeas \registerArray[25][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][7] .is_wysiwyg = "true";
defparam \registerArray[25][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N1
dffeas \registerArray[17][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][7] .is_wysiwyg = "true";
defparam \registerArray[17][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N30
cycloneive_lcell_comb \Mux56~0 (
// Equation(s):
// \Mux56~0_combout  = (\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o ) # ((\registerArray[25][7]~q )))) # (!\my_rf.rsel2[3]~input_o  & (!\my_rf.rsel2[2]~input_o  & ((\registerArray[17][7]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[25][7]~q ),
	.datad(\registerArray[17][7]~q ),
	.cin(gnd),
	.combout(\Mux56~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~0 .lut_mask = 16'hB9A8;
defparam \Mux56~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N12
cycloneive_lcell_comb \Mux56~1 (
// Equation(s):
// \Mux56~1_combout  = (\Mux56~0_combout  & ((\registerArray[29][7]~q ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux56~0_combout  & (((\my_rf.rsel2[2]~input_o  & \registerArray[21][7]~q ))))

	.dataa(\Mux56~0_combout ),
	.datab(\registerArray[29][7]~q ),
	.datac(\my_rf.rsel2[2]~input_o ),
	.datad(\registerArray[21][7]~q ),
	.cin(gnd),
	.combout(\Mux56~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~1 .lut_mask = 16'hDA8A;
defparam \Mux56~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N23
dffeas \registerArray[28][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][7] .is_wysiwyg = "true";
defparam \registerArray[28][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N8
cycloneive_lcell_comb \Mux56~7 (
// Equation(s):
// \Mux56~7_combout  = (\my_rf.rsel2[3]~input_o  & (((\registerArray[27][7]~q ) # (\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[19][7]~q  & ((!\my_rf.rsel2[2]~input_o ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[19][7]~q ),
	.datac(\registerArray[27][7]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux56~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~7 .lut_mask = 16'hAAE4;
defparam \Mux56~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N9
dffeas \registerArray[4][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][7] .is_wysiwyg = "true";
defparam \registerArray[4][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y33_N17
dffeas \registerArray[10][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][7] .is_wysiwyg = "true";
defparam \registerArray[10][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y33_N11
dffeas \registerArray[8][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][7] .is_wysiwyg = "true";
defparam \registerArray[8][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N16
cycloneive_lcell_comb \Mux56~12 (
// Equation(s):
// \Mux56~12_combout  = (\my_rf.rsel2[1]~input_o  & (((\registerArray[10][7]~q ) # (\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[8][7]~q  & ((!\my_rf.rsel2[0]~input_o ))))

	.dataa(\registerArray[8][7]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[10][7]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux56~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~12 .lut_mask = 16'hCCE2;
defparam \Mux56~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N28
cycloneive_lcell_comb \Mux56~13 (
// Equation(s):
// \Mux56~13_combout  = (\Mux56~12_combout  & ((\registerArray[11][7]~q ) # ((!\my_rf.rsel2[0]~input_o )))) # (!\Mux56~12_combout  & (((\registerArray[9][7]~q  & \my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux56~12_combout ),
	.datab(\registerArray[11][7]~q ),
	.datac(\registerArray[9][7]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux56~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~13 .lut_mask = 16'hD8AA;
defparam \Mux56~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N1
dffeas \registerArray[14][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][7] .is_wysiwyg = "true";
defparam \registerArray[14][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N27
dffeas \registerArray[13][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][7] .is_wysiwyg = "true";
defparam \registerArray[13][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N29
dffeas \registerArray[12][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][7] .is_wysiwyg = "true";
defparam \registerArray[12][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N26
cycloneive_lcell_comb \Mux56~17 (
// Equation(s):
// \Mux56~17_combout  = (\my_rf.rsel2[1]~input_o  & (\my_rf.rsel2[0]~input_o )) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & (\registerArray[13][7]~q )) # (!\my_rf.rsel2[0]~input_o  & ((\registerArray[12][7]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[13][7]~q ),
	.datad(\registerArray[12][7]~q ),
	.cin(gnd),
	.combout(\Mux56~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~17 .lut_mask = 16'hD9C8;
defparam \Mux56~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N11
dffeas \registerArray[15][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][7] .is_wysiwyg = "true";
defparam \registerArray[15][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N0
cycloneive_lcell_comb \Mux56~18 (
// Equation(s):
// \Mux56~18_combout  = (\Mux56~17_combout  & (((\registerArray[15][7]~q )) # (!\my_rf.rsel2[1]~input_o ))) # (!\Mux56~17_combout  & (\my_rf.rsel2[1]~input_o  & (\registerArray[14][7]~q )))

	.dataa(\Mux56~17_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][7]~q ),
	.datad(\registerArray[15][7]~q ),
	.cin(gnd),
	.combout(\Mux56~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~18 .lut_mask = 16'hEA62;
defparam \Mux56~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N16
cycloneive_lcell_comb \Mux55~2 (
// Equation(s):
// \Mux55~2_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & ((\registerArray[26][8]~q ))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[18][8]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[18][8]~q ),
	.datac(\registerArray[26][8]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux55~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~2 .lut_mask = 16'hFA44;
defparam \Mux55~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N0
cycloneive_lcell_comb \Mux55~4 (
// Equation(s):
// \Mux55~4_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[24][8]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][8]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][8]~q ),
	.datad(\registerArray[16][8]~q ),
	.cin(gnd),
	.combout(\Mux55~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~4 .lut_mask = 16'hD9C8;
defparam \Mux55~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y33_N11
dffeas \registerArray[27][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][8] .is_wysiwyg = "true";
defparam \registerArray[27][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N5
dffeas \registerArray[23][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][8] .is_wysiwyg = "true";
defparam \registerArray[23][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N4
cycloneive_lcell_comb \Mux55~7 (
// Equation(s):
// \Mux55~7_combout  = (\my_rf.rsel2[3]~input_o  & (\my_rf.rsel2[2]~input_o )) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\registerArray[23][8]~q )) # (!\my_rf.rsel2[2]~input_o  & ((\registerArray[19][8]~q )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[23][8]~q ),
	.datad(\registerArray[19][8]~q ),
	.cin(gnd),
	.combout(\Mux55~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~7 .lut_mask = 16'hD9C8;
defparam \Mux55~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N10
cycloneive_lcell_comb \Mux55~8 (
// Equation(s):
// \Mux55~8_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux55~7_combout  & ((\registerArray[31][8]~q ))) # (!\Mux55~7_combout  & (\registerArray[27][8]~q )))) # (!\my_rf.rsel2[3]~input_o  & (\Mux55~7_combout ))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux55~7_combout ),
	.datac(\registerArray[27][8]~q ),
	.datad(\registerArray[31][8]~q ),
	.cin(gnd),
	.combout(\Mux55~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~8 .lut_mask = 16'hEC64;
defparam \Mux55~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y37_N27
dffeas \registerArray[8][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][8] .is_wysiwyg = "true";
defparam \registerArray[8][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N17
dffeas \registerArray[4][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][8] .is_wysiwyg = "true";
defparam \registerArray[4][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N4
cycloneive_lcell_comb \Mux55~14 (
// Equation(s):
// \Mux55~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][8]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][8]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][8]~q ),
	.datad(\registerArray[1][8]~q ),
	.cin(gnd),
	.combout(\Mux55~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~14 .lut_mask = 16'hC480;
defparam \Mux55~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N12
cycloneive_lcell_comb \Mux54~0 (
// Equation(s):
// \Mux54~0_combout  = (\my_rf.rsel2[3]~input_o  & (((\registerArray[25][9]~q ) # (\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[17][9]~q  & ((!\my_rf.rsel2[2]~input_o ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[17][9]~q ),
	.datac(\registerArray[25][9]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux54~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~0 .lut_mask = 16'hAAE4;
defparam \Mux54~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N23
dffeas \registerArray[19][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][9] .is_wysiwyg = "true";
defparam \registerArray[19][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N29
dffeas \registerArray[5][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][9] .is_wysiwyg = "true";
defparam \registerArray[5][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N3
dffeas \registerArray[4][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][9] .is_wysiwyg = "true";
defparam \registerArray[4][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N28
cycloneive_lcell_comb \Mux54~10 (
// Equation(s):
// \Mux54~10_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[5][9]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][9]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[4][9]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][9]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux54~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~10 .lut_mask = 16'hCCE2;
defparam \Mux54~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y37_N29
dffeas \registerArray[9][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][9] .is_wysiwyg = "true";
defparam \registerArray[9][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y37_N29
dffeas \registerArray[10][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][9] .is_wysiwyg = "true";
defparam \registerArray[10][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y37_N7
dffeas \registerArray[8][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][9] .is_wysiwyg = "true";
defparam \registerArray[8][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y37_N28
cycloneive_lcell_comb \Mux54~12 (
// Equation(s):
// \Mux54~12_combout  = (\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o ) # ((\registerArray[10][9]~q )))) # (!\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & ((\registerArray[8][9]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[10][9]~q ),
	.datad(\registerArray[8][9]~q ),
	.cin(gnd),
	.combout(\Mux54~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~12 .lut_mask = 16'hB9A8;
defparam \Mux54~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y37_N31
dffeas \registerArray[11][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][9] .is_wysiwyg = "true";
defparam \registerArray[11][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y37_N28
cycloneive_lcell_comb \Mux54~13 (
// Equation(s):
// \Mux54~13_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux54~12_combout  & (\registerArray[11][9]~q )) # (!\Mux54~12_combout  & ((\registerArray[9][9]~q ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux54~12_combout ))))

	.dataa(\registerArray[11][9]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[9][9]~q ),
	.datad(\Mux54~12_combout ),
	.cin(gnd),
	.combout(\Mux54~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~13 .lut_mask = 16'hBBC0;
defparam \Mux54~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N8
cycloneive_lcell_comb \Mux54~14 (
// Equation(s):
// \Mux54~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][9]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][9]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][9]~q ),
	.datad(\registerArray[1][9]~q ),
	.cin(gnd),
	.combout(\Mux54~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~14 .lut_mask = 16'hC480;
defparam \Mux54~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N1
dffeas \registerArray[14][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][9] .is_wysiwyg = "true";
defparam \registerArray[14][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N11
dffeas \registerArray[13][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][9] .is_wysiwyg = "true";
defparam \registerArray[13][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N21
dffeas \registerArray[12][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][9] .is_wysiwyg = "true";
defparam \registerArray[12][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N10
cycloneive_lcell_comb \Mux54~17 (
// Equation(s):
// \Mux54~17_combout  = (\my_rf.rsel2[1]~input_o  & (\my_rf.rsel2[0]~input_o )) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & (\registerArray[13][9]~q )) # (!\my_rf.rsel2[0]~input_o  & ((\registerArray[12][9]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[13][9]~q ),
	.datad(\registerArray[12][9]~q ),
	.cin(gnd),
	.combout(\Mux54~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~17 .lut_mask = 16'hD9C8;
defparam \Mux54~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N19
dffeas \registerArray[15][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][9] .is_wysiwyg = "true";
defparam \registerArray[15][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N0
cycloneive_lcell_comb \Mux54~18 (
// Equation(s):
// \Mux54~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux54~17_combout  & ((\registerArray[15][9]~q ))) # (!\Mux54~17_combout  & (\registerArray[14][9]~q )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux54~17_combout ))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux54~17_combout ),
	.datac(\registerArray[14][9]~q ),
	.datad(\registerArray[15][9]~q ),
	.cin(gnd),
	.combout(\Mux54~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~18 .lut_mask = 16'hEC64;
defparam \Mux54~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y0_N3
dffeas \registerArray[25][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[10]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][10] .is_wysiwyg = "true";
defparam \registerArray[25][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N9
dffeas \registerArray[21][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][10] .is_wysiwyg = "true";
defparam \registerArray[21][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N27
dffeas \registerArray[17][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][10] .is_wysiwyg = "true";
defparam \registerArray[17][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N8
cycloneive_lcell_comb \Mux53~0 (
// Equation(s):
// \Mux53~0_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & ((\registerArray[21][10]~q ))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[17][10]~q ))))

	.dataa(\registerArray[17][10]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[21][10]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux53~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~0 .lut_mask = 16'hFC22;
defparam \Mux53~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y34_N1
dffeas \registerArray[29][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][10] .is_wysiwyg = "true";
defparam \registerArray[29][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N18
cycloneive_lcell_comb \Mux53~1 (
// Equation(s):
// \Mux53~1_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux53~0_combout  & (\registerArray[29][10]~q )) # (!\Mux53~0_combout  & ((\registerArray[25][10]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux53~0_combout ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[29][10]~q ),
	.datac(\registerArray[25][10]~q ),
	.datad(\Mux53~0_combout ),
	.cin(gnd),
	.combout(\Mux53~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~1 .lut_mask = 16'hDDA0;
defparam \Mux53~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y36_N21
dffeas \registerArray[22][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][10] .is_wysiwyg = "true";
defparam \registerArray[22][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y36_N25
dffeas \registerArray[26][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][10] .is_wysiwyg = "true";
defparam \registerArray[26][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y36_N23
dffeas \registerArray[18][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][10] .is_wysiwyg = "true";
defparam \registerArray[18][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N24
cycloneive_lcell_comb \Mux53~2 (
// Equation(s):
// \Mux53~2_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[26][10]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[18][10]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[26][10]~q ),
	.datad(\registerArray[18][10]~q ),
	.cin(gnd),
	.combout(\Mux53~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~2 .lut_mask = 16'hD9C8;
defparam \Mux53~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y36_N11
dffeas \registerArray[30][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][10] .is_wysiwyg = "true";
defparam \registerArray[30][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N20
cycloneive_lcell_comb \Mux53~3 (
// Equation(s):
// \Mux53~3_combout  = (\Mux53~2_combout  & (((\registerArray[30][10]~q )) # (!\my_rf.rsel2[2]~input_o ))) # (!\Mux53~2_combout  & (\my_rf.rsel2[2]~input_o  & (\registerArray[22][10]~q )))

	.dataa(\Mux53~2_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][10]~q ),
	.datad(\registerArray[30][10]~q ),
	.cin(gnd),
	.combout(\Mux53~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~3 .lut_mask = 16'hEA62;
defparam \Mux53~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y37_N9
dffeas \registerArray[10][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][10] .is_wysiwyg = "true";
defparam \registerArray[10][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y37_N11
dffeas \registerArray[8][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][10] .is_wysiwyg = "true";
defparam \registerArray[8][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y37_N8
cycloneive_lcell_comb \Mux53~10 (
// Equation(s):
// \Mux53~10_combout  = (\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o ) # ((\registerArray[10][10]~q )))) # (!\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & ((\registerArray[8][10]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[10][10]~q ),
	.datad(\registerArray[8][10]~q ),
	.cin(gnd),
	.combout(\Mux53~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~10 .lut_mask = 16'hB9A8;
defparam \Mux53~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y37_N8
cycloneive_lcell_comb \Mux53~11 (
// Equation(s):
// \Mux53~11_combout  = (\Mux53~10_combout  & (((\registerArray[11][10]~q )) # (!\my_rf.rsel2[0]~input_o ))) # (!\Mux53~10_combout  & (\my_rf.rsel2[0]~input_o  & (\registerArray[9][10]~q )))

	.dataa(\Mux53~10_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[9][10]~q ),
	.datad(\registerArray[11][10]~q ),
	.cin(gnd),
	.combout(\Mux53~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~11 .lut_mask = 16'hEA62;
defparam \Mux53~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X0_Y34_N10
dffeas \registerArray[21][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[11]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][11] .is_wysiwyg = "true";
defparam \registerArray[21][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N19
dffeas \registerArray[25][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][11] .is_wysiwyg = "true";
defparam \registerArray[25][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N18
cycloneive_lcell_comb \Mux52~0 (
// Equation(s):
// \Mux52~0_combout  = (\my_rf.rsel2[3]~input_o  & (((\registerArray[25][11]~q ) # (\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[17][11]~q  & ((!\my_rf.rsel2[2]~input_o ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[17][11]~q ),
	.datac(\registerArray[25][11]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux52~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~0 .lut_mask = 16'hAAE4;
defparam \Mux52~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N30
cycloneive_lcell_comb \Mux52~1 (
// Equation(s):
// \Mux52~1_combout  = (\Mux52~0_combout  & (((\registerArray[29][11]~q ) # (!\my_rf.rsel2[2]~input_o )))) # (!\Mux52~0_combout  & (\registerArray[21][11]~q  & ((\my_rf.rsel2[2]~input_o ))))

	.dataa(\registerArray[21][11]~q ),
	.datab(\Mux52~0_combout ),
	.datac(\registerArray[29][11]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux52~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~1 .lut_mask = 16'hE2CC;
defparam \Mux52~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N9
dffeas \registerArray[24][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][11] .is_wysiwyg = "true";
defparam \registerArray[24][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N0
cycloneive_lcell_comb \Mux52~4 (
// Equation(s):
// \Mux52~4_combout  = (\my_rf.rsel2[3]~input_o  & (\my_rf.rsel2[2]~input_o )) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\registerArray[20][11]~q )) # (!\my_rf.rsel2[2]~input_o  & ((\registerArray[16][11]~q )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[20][11]~q ),
	.datad(\registerArray[16][11]~q ),
	.cin(gnd),
	.combout(\Mux52~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~4 .lut_mask = 16'hD9C8;
defparam \Mux52~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N8
cycloneive_lcell_comb \Mux52~5 (
// Equation(s):
// \Mux52~5_combout  = (\Mux52~4_combout  & ((\registerArray[28][11]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux52~4_combout  & (((\registerArray[24][11]~q  & \my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[28][11]~q ),
	.datab(\Mux52~4_combout ),
	.datac(\registerArray[24][11]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux52~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~5 .lut_mask = 16'hB8CC;
defparam \Mux52~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y37_N5
dffeas \registerArray[10][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][11] .is_wysiwyg = "true";
defparam \registerArray[10][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y37_N31
dffeas \registerArray[8][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][11] .is_wysiwyg = "true";
defparam \registerArray[8][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y37_N4
cycloneive_lcell_comb \Mux52~12 (
// Equation(s):
// \Mux52~12_combout  = (\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o ) # ((\registerArray[10][11]~q )))) # (!\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & ((\registerArray[8][11]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[10][11]~q ),
	.datad(\registerArray[8][11]~q ),
	.cin(gnd),
	.combout(\Mux52~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~12 .lut_mask = 16'hB9A8;
defparam \Mux52~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y37_N29
dffeas \registerArray[13][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][11] .is_wysiwyg = "true";
defparam \registerArray[13][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N15
dffeas \registerArray[12][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][11] .is_wysiwyg = "true";
defparam \registerArray[12][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N28
cycloneive_lcell_comb \Mux52~17 (
// Equation(s):
// \Mux52~17_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & ((\registerArray[13][11]~q ))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[12][11]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[12][11]~q ),
	.datac(\registerArray[13][11]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux52~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~17 .lut_mask = 16'hFA44;
defparam \Mux52~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N16
cycloneive_lcell_comb \Mux52~18 (
// Equation(s):
// \Mux52~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux52~17_combout  & (\registerArray[15][11]~q )) # (!\Mux52~17_combout  & ((\registerArray[14][11]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux52~17_combout ))))

	.dataa(\registerArray[15][11]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][11]~q ),
	.datad(\Mux52~17_combout ),
	.cin(gnd),
	.combout(\Mux52~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~18 .lut_mask = 16'hBBC0;
defparam \Mux52~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y32_N31
dffeas \registerArray[21][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][12] .is_wysiwyg = "true";
defparam \registerArray[21][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N30
cycloneive_lcell_comb \Mux51~0 (
// Equation(s):
// \Mux51~0_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[21][12]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[17][12]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[21][12]~q ),
	.datad(\registerArray[17][12]~q ),
	.cin(gnd),
	.combout(\Mux51~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~0 .lut_mask = 16'hB9A8;
defparam \Mux51~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y36_N29
dffeas \registerArray[22][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][12] .is_wysiwyg = "true";
defparam \registerArray[22][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y37_N11
dffeas \registerArray[26][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][12] .is_wysiwyg = "true";
defparam \registerArray[26][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y36_N15
dffeas \registerArray[18][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][12] .is_wysiwyg = "true";
defparam \registerArray[18][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y37_N10
cycloneive_lcell_comb \Mux51~2 (
// Equation(s):
// \Mux51~2_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[26][12]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[18][12]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[26][12]~q ),
	.datad(\registerArray[18][12]~q ),
	.cin(gnd),
	.combout(\Mux51~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~2 .lut_mask = 16'hD9C8;
defparam \Mux51~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y35_N1
dffeas \registerArray[30][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][12] .is_wysiwyg = "true";
defparam \registerArray[30][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N28
cycloneive_lcell_comb \Mux51~3 (
// Equation(s):
// \Mux51~3_combout  = (\Mux51~2_combout  & (((\registerArray[30][12]~q )) # (!\my_rf.rsel2[2]~input_o ))) # (!\Mux51~2_combout  & (\my_rf.rsel2[2]~input_o  & (\registerArray[22][12]~q )))

	.dataa(\Mux51~2_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][12]~q ),
	.datad(\registerArray[30][12]~q ),
	.cin(gnd),
	.combout(\Mux51~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~3 .lut_mask = 16'hEA62;
defparam \Mux51~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y32_N1
dffeas \registerArray[23][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][12] .is_wysiwyg = "true";
defparam \registerArray[23][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N0
cycloneive_lcell_comb \Mux51~7 (
// Equation(s):
// \Mux51~7_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & ((\registerArray[23][12]~q ))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[19][12]~q ))))

	.dataa(\registerArray[19][12]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[23][12]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux51~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~7 .lut_mask = 16'hFC22;
defparam \Mux51~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N0
cycloneive_lcell_comb \Mux51~8 (
// Equation(s):
// \Mux51~8_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux51~7_combout  & ((\registerArray[31][12]~q ))) # (!\Mux51~7_combout  & (\registerArray[27][12]~q )))) # (!\my_rf.rsel2[3]~input_o  & (\Mux51~7_combout ))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux51~7_combout ),
	.datac(\registerArray[27][12]~q ),
	.datad(\registerArray[31][12]~q ),
	.cin(gnd),
	.combout(\Mux51~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~8 .lut_mask = 16'hEC64;
defparam \Mux51~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y37_N1
dffeas \registerArray[10][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][12] .is_wysiwyg = "true";
defparam \registerArray[10][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y37_N3
dffeas \registerArray[8][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][12] .is_wysiwyg = "true";
defparam \registerArray[8][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y37_N0
cycloneive_lcell_comb \Mux51~10 (
// Equation(s):
// \Mux51~10_combout  = (\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o ) # ((\registerArray[10][12]~q )))) # (!\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & ((\registerArray[8][12]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[10][12]~q ),
	.datad(\registerArray[8][12]~q ),
	.cin(gnd),
	.combout(\Mux51~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~10 .lut_mask = 16'hB9A8;
defparam \Mux51~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N27
dffeas \registerArray[7][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][12] .is_wysiwyg = "true";
defparam \registerArray[7][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N20
cycloneive_lcell_comb \Mux51~14 (
// Equation(s):
// \Mux51~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][12]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][12]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][12]~q ),
	.datad(\registerArray[1][12]~q ),
	.cin(gnd),
	.combout(\Mux51~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~14 .lut_mask = 16'hC480;
defparam \Mux51~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N12
cycloneive_lcell_comb \Mux51~15 (
// Equation(s):
// \Mux51~15_combout  = (\Mux51~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][12]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][12]~q ),
	.datad(\Mux51~14_combout ),
	.cin(gnd),
	.combout(\Mux51~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~15 .lut_mask = 16'hFF20;
defparam \Mux51~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N9
dffeas \registerArray[25][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][13] .is_wysiwyg = "true";
defparam \registerArray[25][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N11
dffeas \registerArray[17][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][13] .is_wysiwyg = "true";
defparam \registerArray[17][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N8
cycloneive_lcell_comb \Mux50~0 (
// Equation(s):
// \Mux50~0_combout  = (\my_rf.rsel2[3]~input_o  & (((\registerArray[25][13]~q ) # (\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[17][13]~q  & ((!\my_rf.rsel2[2]~input_o ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[17][13]~q ),
	.datac(\registerArray[25][13]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux50~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~0 .lut_mask = 16'hAAE4;
defparam \Mux50~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N4
cycloneive_lcell_comb \Mux50~1 (
// Equation(s):
// \Mux50~1_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux50~0_combout  & ((\registerArray[29][13]~q ))) # (!\Mux50~0_combout  & (\registerArray[21][13]~q )))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux50~0_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[21][13]~q ),
	.datac(\Mux50~0_combout ),
	.datad(\registerArray[29][13]~q ),
	.cin(gnd),
	.combout(\Mux50~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~1 .lut_mask = 16'hF858;
defparam \Mux50~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N24
cycloneive_lcell_comb \Mux50~2 (
// Equation(s):
// \Mux50~2_combout  = (\my_rf.rsel2[3]~input_o  & (\my_rf.rsel2[2]~input_o )) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\registerArray[22][13]~q )) # (!\my_rf.rsel2[2]~input_o  & ((\registerArray[18][13]~q )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][13]~q ),
	.datad(\registerArray[18][13]~q ),
	.cin(gnd),
	.combout(\Mux50~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~2 .lut_mask = 16'hD9C8;
defparam \Mux50~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N13
dffeas \registerArray[24][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][13] .is_wysiwyg = "true";
defparam \registerArray[24][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N8
cycloneive_lcell_comb \Mux50~4 (
// Equation(s):
// \Mux50~4_combout  = (\my_rf.rsel2[3]~input_o  & (\my_rf.rsel2[2]~input_o )) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\registerArray[20][13]~q )) # (!\my_rf.rsel2[2]~input_o  & ((\registerArray[16][13]~q )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[20][13]~q ),
	.datad(\registerArray[16][13]~q ),
	.cin(gnd),
	.combout(\Mux50~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~4 .lut_mask = 16'hD9C8;
defparam \Mux50~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N12
cycloneive_lcell_comb \Mux50~5 (
// Equation(s):
// \Mux50~5_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux50~4_combout  & (\registerArray[28][13]~q )) # (!\Mux50~4_combout  & ((\registerArray[24][13]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux50~4_combout ))))

	.dataa(\registerArray[28][13]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][13]~q ),
	.datad(\Mux50~4_combout ),
	.cin(gnd),
	.combout(\Mux50~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~5 .lut_mask = 16'hBBC0;
defparam \Mux50~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y37_N11
dffeas \registerArray[9][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][13] .is_wysiwyg = "true";
defparam \registerArray[9][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y37_N21
dffeas \registerArray[10][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][13] .is_wysiwyg = "true";
defparam \registerArray[10][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y37_N15
dffeas \registerArray[8][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][13] .is_wysiwyg = "true";
defparam \registerArray[8][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y37_N20
cycloneive_lcell_comb \Mux50~12 (
// Equation(s):
// \Mux50~12_combout  = (\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o ) # ((\registerArray[10][13]~q )))) # (!\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & ((\registerArray[8][13]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[10][13]~q ),
	.datad(\registerArray[8][13]~q ),
	.cin(gnd),
	.combout(\Mux50~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~12 .lut_mask = 16'hB9A8;
defparam \Mux50~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y37_N5
dffeas \registerArray[11][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][13] .is_wysiwyg = "true";
defparam \registerArray[11][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y37_N10
cycloneive_lcell_comb \Mux50~13 (
// Equation(s):
// \Mux50~13_combout  = (\Mux50~12_combout  & ((\registerArray[11][13]~q ) # ((!\my_rf.rsel2[0]~input_o )))) # (!\Mux50~12_combout  & (((\registerArray[9][13]~q  & \my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux50~12_combout ),
	.datab(\registerArray[11][13]~q ),
	.datac(\registerArray[9][13]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux50~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~13 .lut_mask = 16'hD8AA;
defparam \Mux50~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y36_N1
dffeas \registerArray[3][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][13] .is_wysiwyg = "true";
defparam \registerArray[3][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N27
dffeas \registerArray[1][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][13] .is_wysiwyg = "true";
defparam \registerArray[1][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N0
cycloneive_lcell_comb \Mux50~14 (
// Equation(s):
// \Mux50~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[3][13]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[1][13]~q ))))

	.dataa(\registerArray[1][13]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][13]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux50~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~14 .lut_mask = 16'hC088;
defparam \Mux50~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N17
dffeas \registerArray[2][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][13] .is_wysiwyg = "true";
defparam \registerArray[2][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N16
cycloneive_lcell_comb \Mux50~15 (
// Equation(s):
// \Mux50~15_combout  = (\Mux50~14_combout ) # ((!\my_rf.rsel2[0]~input_o  & (\registerArray[2][13]~q  & \my_rf.rsel2[1]~input_o )))

	.dataa(\Mux50~14_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][13]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux50~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~15 .lut_mask = 16'hBAAA;
defparam \Mux50~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y37_N6
cycloneive_lcell_comb \Mux50~16 (
// Equation(s):
// \Mux50~16_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o ) # (\Mux50~13_combout )))) # (!\my_rf.rsel2[3]~input_o  & (\Mux50~15_combout  & (!\my_rf.rsel2[2]~input_o )))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux50~15_combout ),
	.datac(\my_rf.rsel2[2]~input_o ),
	.datad(\Mux50~13_combout ),
	.cin(gnd),
	.combout(\Mux50~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~16 .lut_mask = 16'hAEA4;
defparam \Mux50~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y38_N21
dffeas \registerArray[30][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][14] .is_wysiwyg = "true";
defparam \registerArray[30][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y37_N23
dffeas \registerArray[28][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][14] .is_wysiwyg = "true";
defparam \registerArray[28][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y32_N19
dffeas \registerArray[23][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][14] .is_wysiwyg = "true";
defparam \registerArray[23][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N31
dffeas \registerArray[19][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][14] .is_wysiwyg = "true";
defparam \registerArray[19][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N18
cycloneive_lcell_comb \Mux49~7 (
// Equation(s):
// \Mux49~7_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & ((\registerArray[23][14]~q ))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[19][14]~q ))))

	.dataa(\registerArray[19][14]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[23][14]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux49~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~7 .lut_mask = 16'hFC22;
defparam \Mux49~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y37_N16
cycloneive_lcell_comb \Mux49~10 (
// Equation(s):
// \Mux49~10_combout  = (\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o ) # ((\registerArray[10][14]~q )))) # (!\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & ((\registerArray[8][14]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[10][14]~q ),
	.datad(\registerArray[8][14]~q ),
	.cin(gnd),
	.combout(\Mux49~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~10 .lut_mask = 16'hB9A8;
defparam \Mux49~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N9
dffeas \registerArray[5][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][14] .is_wysiwyg = "true";
defparam \registerArray[5][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N19
dffeas \registerArray[4][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][14] .is_wysiwyg = "true";
defparam \registerArray[4][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N8
cycloneive_lcell_comb \Mux49~12 (
// Equation(s):
// \Mux49~12_combout  = (\my_rf.rsel2[1]~input_o  & (\my_rf.rsel2[0]~input_o )) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & (\registerArray[5][14]~q )) # (!\my_rf.rsel2[0]~input_o  & ((\registerArray[4][14]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][14]~q ),
	.datad(\registerArray[4][14]~q ),
	.cin(gnd),
	.combout(\Mux49~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~12 .lut_mask = 16'hD9C8;
defparam \Mux49~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N0
cycloneive_lcell_comb \Mux49~13 (
// Equation(s):
// \Mux49~13_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux49~12_combout  & ((\registerArray[7][14]~q ))) # (!\Mux49~12_combout  & (\registerArray[6][14]~q )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux49~12_combout ))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux49~12_combout ),
	.datac(\registerArray[6][14]~q ),
	.datad(\registerArray[7][14]~q ),
	.cin(gnd),
	.combout(\Mux49~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~13 .lut_mask = 16'hEC64;
defparam \Mux49~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N4
cycloneive_lcell_comb \Mux49~14 (
// Equation(s):
// \Mux49~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[3][14]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[1][14]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\registerArray[1][14]~q ),
	.datac(\registerArray[3][14]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux49~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~14 .lut_mask = 16'hA088;
defparam \Mux49~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N22
cycloneive_lcell_comb \Mux49~15 (
// Equation(s):
// \Mux49~15_combout  = (\Mux49~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][14]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][14]~q ),
	.datad(\Mux49~14_combout ),
	.cin(gnd),
	.combout(\Mux49~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~15 .lut_mask = 16'hFF20;
defparam \Mux49~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y30_N0
cycloneive_lcell_comb \Mux49~16 (
// Equation(s):
// \Mux49~16_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\Mux49~13_combout )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\Mux49~15_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux49~13_combout ),
	.datad(\Mux49~15_combout ),
	.cin(gnd),
	.combout(\Mux49~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~16 .lut_mask = 16'hB9A8;
defparam \Mux49~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y36_N31
dffeas \registerArray[12][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][14] .is_wysiwyg = "true";
defparam \registerArray[12][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N0
cycloneive_lcell_comb \Mux48~2 (
// Equation(s):
// \Mux48~2_combout  = (\my_rf.rsel2[3]~input_o  & (\my_rf.rsel2[2]~input_o )) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\registerArray[22][15]~q )) # (!\my_rf.rsel2[2]~input_o  & ((\registerArray[18][15]~q )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][15]~q ),
	.datad(\registerArray[18][15]~q ),
	.cin(gnd),
	.combout(\Mux48~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~2 .lut_mask = 16'hD9C8;
defparam \Mux48~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y35_N1
dffeas \registerArray[28][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][15] .is_wysiwyg = "true";
defparam \registerArray[28][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y33_N27
dffeas \registerArray[31][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][15] .is_wysiwyg = "true";
defparam \registerArray[31][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y39_N1
dffeas \registerArray[9][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][15] .is_wysiwyg = "true";
defparam \registerArray[9][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y39_N9
dffeas \registerArray[10][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][15] .is_wysiwyg = "true";
defparam \registerArray[10][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y39_N19
dffeas \registerArray[8][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][15] .is_wysiwyg = "true";
defparam \registerArray[8][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N8
cycloneive_lcell_comb \Mux48~12 (
// Equation(s):
// \Mux48~12_combout  = (\my_rf.rsel2[0]~input_o  & (\my_rf.rsel2[1]~input_o )) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[10][15]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[8][15]~q )))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[10][15]~q ),
	.datad(\registerArray[8][15]~q ),
	.cin(gnd),
	.combout(\Mux48~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~12 .lut_mask = 16'hD9C8;
defparam \Mux48~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N19
dffeas \registerArray[11][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][15] .is_wysiwyg = "true";
defparam \registerArray[11][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N0
cycloneive_lcell_comb \Mux48~13 (
// Equation(s):
// \Mux48~13_combout  = (\Mux48~12_combout  & (((\registerArray[11][15]~q )) # (!\my_rf.rsel2[0]~input_o ))) # (!\Mux48~12_combout  & (\my_rf.rsel2[0]~input_o  & (\registerArray[9][15]~q )))

	.dataa(\Mux48~12_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[9][15]~q ),
	.datad(\registerArray[11][15]~q ),
	.cin(gnd),
	.combout(\Mux48~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~13 .lut_mask = 16'hEA62;
defparam \Mux48~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y36_N1
dffeas \registerArray[13][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][15] .is_wysiwyg = "true";
defparam \registerArray[13][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y36_N11
dffeas \registerArray[12][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][15] .is_wysiwyg = "true";
defparam \registerArray[12][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y36_N0
cycloneive_lcell_comb \Mux48~17 (
// Equation(s):
// \Mux48~17_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[13][15]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[12][15]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[13][15]~q ),
	.datad(\registerArray[12][15]~q ),
	.cin(gnd),
	.combout(\Mux48~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~17 .lut_mask = 16'hB9A8;
defparam \Mux48~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N4
cycloneive_lcell_comb \Mux48~18 (
// Equation(s):
// \Mux48~18_combout  = (\Mux48~17_combout  & ((\registerArray[15][15]~q ) # ((!\my_rf.rsel2[1]~input_o )))) # (!\Mux48~17_combout  & (((\registerArray[14][15]~q  & \my_rf.rsel2[1]~input_o ))))

	.dataa(\Mux48~17_combout ),
	.datab(\registerArray[15][15]~q ),
	.datac(\registerArray[14][15]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux48~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~18 .lut_mask = 16'hD8AA;
defparam \Mux48~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N14
cycloneive_lcell_comb \Mux47~2 (
// Equation(s):
// \Mux47~2_combout  = (\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o ) # ((\registerArray[26][16]~q )))) # (!\my_rf.rsel2[3]~input_o  & (!\my_rf.rsel2[2]~input_o  & ((\registerArray[18][16]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[26][16]~q ),
	.datad(\registerArray[18][16]~q ),
	.cin(gnd),
	.combout(\Mux47~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~2 .lut_mask = 16'hB9A8;
defparam \Mux47~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y35_N27
dffeas \registerArray[24][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][16] .is_wysiwyg = "true";
defparam \registerArray[24][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y35_N3
dffeas \registerArray[16][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][16] .is_wysiwyg = "true";
defparam \registerArray[16][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N26
cycloneive_lcell_comb \Mux47~4 (
// Equation(s):
// \Mux47~4_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & ((\registerArray[24][16]~q ))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[16][16]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[16][16]~q ),
	.datac(\registerArray[24][16]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux47~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~4 .lut_mask = 16'hFA44;
defparam \Mux47~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N8
cycloneive_lcell_comb \Mux47~5 (
// Equation(s):
// \Mux47~5_combout  = (\Mux47~4_combout  & ((\registerArray[28][16]~q ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux47~4_combout  & (((\registerArray[20][16]~q  & \my_rf.rsel2[2]~input_o ))))

	.dataa(\registerArray[28][16]~q ),
	.datab(\Mux47~4_combout ),
	.datac(\registerArray[20][16]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux47~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~5 .lut_mask = 16'hB8CC;
defparam \Mux47~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y33_N31
dffeas \registerArray[27][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][16] .is_wysiwyg = "true";
defparam \registerArray[27][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y33_N29
dffeas \registerArray[23][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][16] .is_wysiwyg = "true";
defparam \registerArray[23][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y33_N25
dffeas \registerArray[19][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][16] .is_wysiwyg = "true";
defparam \registerArray[19][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N28
cycloneive_lcell_comb \Mux47~7 (
// Equation(s):
// \Mux47~7_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[23][16]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[19][16]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[23][16]~q ),
	.datad(\registerArray[19][16]~q ),
	.cin(gnd),
	.combout(\Mux47~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~7 .lut_mask = 16'hB9A8;
defparam \Mux47~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y33_N15
dffeas \registerArray[31][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][16] .is_wysiwyg = "true";
defparam \registerArray[31][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N30
cycloneive_lcell_comb \Mux47~8 (
// Equation(s):
// \Mux47~8_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux47~7_combout  & (\registerArray[31][16]~q )) # (!\Mux47~7_combout  & ((\registerArray[27][16]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux47~7_combout ))))

	.dataa(\registerArray[31][16]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][16]~q ),
	.datad(\Mux47~7_combout ),
	.cin(gnd),
	.combout(\Mux47~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~8 .lut_mask = 16'hBBC0;
defparam \Mux47~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N28
cycloneive_lcell_comb \Mux47~10 (
// Equation(s):
// \Mux47~10_combout  = (\my_rf.rsel2[0]~input_o  & (\my_rf.rsel2[1]~input_o )) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[10][16]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[8][16]~q )))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[10][16]~q ),
	.datad(\registerArray[8][16]~q ),
	.cin(gnd),
	.combout(\Mux47~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~10 .lut_mask = 16'hD9C8;
defparam \Mux47~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y37_N13
dffeas \registerArray[6][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][16] .is_wysiwyg = "true";
defparam \registerArray[6][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N25
dffeas \registerArray[5][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][16] .is_wysiwyg = "true";
defparam \registerArray[5][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N19
dffeas \registerArray[4][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][16] .is_wysiwyg = "true";
defparam \registerArray[4][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N24
cycloneive_lcell_comb \Mux47~12 (
// Equation(s):
// \Mux47~12_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[5][16]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[4][16]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[5][16]~q ),
	.datad(\registerArray[4][16]~q ),
	.cin(gnd),
	.combout(\Mux47~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~12 .lut_mask = 16'hB9A8;
defparam \Mux47~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y37_N15
dffeas \registerArray[7][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][16] .is_wysiwyg = "true";
defparam \registerArray[7][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N12
cycloneive_lcell_comb \Mux47~13 (
// Equation(s):
// \Mux47~13_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux47~12_combout  & (\registerArray[7][16]~q )) # (!\Mux47~12_combout  & ((\registerArray[6][16]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux47~12_combout ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[7][16]~q ),
	.datac(\registerArray[6][16]~q ),
	.datad(\Mux47~12_combout ),
	.cin(gnd),
	.combout(\Mux47~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~13 .lut_mask = 16'hDDA0;
defparam \Mux47~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N8
cycloneive_lcell_comb \Mux47~14 (
// Equation(s):
// \Mux47~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][16]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][16]~q )))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[3][16]~q ),
	.datad(\registerArray[1][16]~q ),
	.cin(gnd),
	.combout(\Mux47~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~14 .lut_mask = 16'hA280;
defparam \Mux47~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N0
cycloneive_lcell_comb \Mux47~15 (
// Equation(s):
// \Mux47~15_combout  = (\Mux47~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][16]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][16]~q ),
	.datad(\Mux47~14_combout ),
	.cin(gnd),
	.combout(\Mux47~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~15 .lut_mask = 16'hFF20;
defparam \Mux47~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N22
cycloneive_lcell_comb \Mux47~16 (
// Equation(s):
// \Mux47~16_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux47~13_combout ) # ((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux47~15_combout  & !\my_rf.rsel2[3]~input_o ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux47~13_combout ),
	.datac(\Mux47~15_combout ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux47~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~16 .lut_mask = 16'hAAD8;
defparam \Mux47~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y36_N13
dffeas \registerArray[13][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][16] .is_wysiwyg = "true";
defparam \registerArray[13][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y36_N7
dffeas \registerArray[12][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][16] .is_wysiwyg = "true";
defparam \registerArray[12][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y36_N12
cycloneive_lcell_comb \Mux47~17 (
// Equation(s):
// \Mux47~17_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[13][16]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[12][16]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[13][16]~q ),
	.datad(\registerArray[12][16]~q ),
	.cin(gnd),
	.combout(\Mux47~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~17 .lut_mask = 16'hB9A8;
defparam \Mux47~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N31
dffeas \registerArray[25][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][17] .is_wysiwyg = "true";
defparam \registerArray[25][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N23
dffeas \registerArray[17][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][17] .is_wysiwyg = "true";
defparam \registerArray[17][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N30
cycloneive_lcell_comb \Mux46~0 (
// Equation(s):
// \Mux46~0_combout  = (\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o ) # ((\registerArray[25][17]~q )))) # (!\my_rf.rsel2[3]~input_o  & (!\my_rf.rsel2[2]~input_o  & ((\registerArray[17][17]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[25][17]~q ),
	.datad(\registerArray[17][17]~q ),
	.cin(gnd),
	.combout(\Mux46~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~0 .lut_mask = 16'hB9A8;
defparam \Mux46~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N4
cycloneive_lcell_comb \Mux46~4 (
// Equation(s):
// \Mux46~4_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[20][17]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][17]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[20][17]~q ),
	.datad(\registerArray[16][17]~q ),
	.cin(gnd),
	.combout(\Mux46~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~4 .lut_mask = 16'hB9A8;
defparam \Mux46~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N18
cycloneive_lcell_comb \Mux46~5 (
// Equation(s):
// \Mux46~5_combout  = (\Mux46~4_combout  & (((\registerArray[28][17]~q )) # (!\my_rf.rsel2[3]~input_o ))) # (!\Mux46~4_combout  & (\my_rf.rsel2[3]~input_o  & (\registerArray[24][17]~q )))

	.dataa(\Mux46~4_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][17]~q ),
	.datad(\registerArray[28][17]~q ),
	.cin(gnd),
	.combout(\Mux46~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~5 .lut_mask = 16'hEA62;
defparam \Mux46~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N5
dffeas \registerArray[27][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][17] .is_wysiwyg = "true";
defparam \registerArray[27][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N15
dffeas \registerArray[19][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][17] .is_wysiwyg = "true";
defparam \registerArray[19][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N4
cycloneive_lcell_comb \Mux46~7 (
// Equation(s):
// \Mux46~7_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & ((\registerArray[27][17]~q ))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[19][17]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[19][17]~q ),
	.datac(\registerArray[27][17]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux46~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~7 .lut_mask = 16'hFA44;
defparam \Mux46~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N24
cycloneive_lcell_comb \Mux46~8 (
// Equation(s):
// \Mux46~8_combout  = (\Mux46~7_combout  & ((\registerArray[31][17]~q ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux46~7_combout  & (((\registerArray[23][17]~q  & \my_rf.rsel2[2]~input_o ))))

	.dataa(\registerArray[31][17]~q ),
	.datab(\Mux46~7_combout ),
	.datac(\registerArray[23][17]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux46~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~8 .lut_mask = 16'hB8CC;
defparam \Mux46~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N21
dffeas \registerArray[5][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][17] .is_wysiwyg = "true";
defparam \registerArray[5][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N23
dffeas \registerArray[4][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][17] .is_wysiwyg = "true";
defparam \registerArray[4][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N20
cycloneive_lcell_comb \Mux46~10 (
// Equation(s):
// \Mux46~10_combout  = (\my_rf.rsel2[1]~input_o  & (\my_rf.rsel2[0]~input_o )) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & (\registerArray[5][17]~q )) # (!\my_rf.rsel2[0]~input_o  & ((\registerArray[4][17]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][17]~q ),
	.datad(\registerArray[4][17]~q ),
	.cin(gnd),
	.combout(\Mux46~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~10 .lut_mask = 16'hD9C8;
defparam \Mux46~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N9
dffeas \registerArray[9][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][17] .is_wysiwyg = "true";
defparam \registerArray[9][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y39_N17
dffeas \registerArray[10][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][17] .is_wysiwyg = "true";
defparam \registerArray[10][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y39_N3
dffeas \registerArray[8][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][17] .is_wysiwyg = "true";
defparam \registerArray[8][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N16
cycloneive_lcell_comb \Mux46~12 (
// Equation(s):
// \Mux46~12_combout  = (\my_rf.rsel2[0]~input_o  & (\my_rf.rsel2[1]~input_o )) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[10][17]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[8][17]~q )))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[10][17]~q ),
	.datad(\registerArray[8][17]~q ),
	.cin(gnd),
	.combout(\Mux46~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~12 .lut_mask = 16'hD9C8;
defparam \Mux46~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N3
dffeas \registerArray[11][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][17] .is_wysiwyg = "true";
defparam \registerArray[11][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N8
cycloneive_lcell_comb \Mux46~13 (
// Equation(s):
// \Mux46~13_combout  = (\Mux46~12_combout  & (((\registerArray[11][17]~q )) # (!\my_rf.rsel2[0]~input_o ))) # (!\Mux46~12_combout  & (\my_rf.rsel2[0]~input_o  & (\registerArray[9][17]~q )))

	.dataa(\Mux46~12_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[9][17]~q ),
	.datad(\registerArray[11][17]~q ),
	.cin(gnd),
	.combout(\Mux46~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~13 .lut_mask = 16'hEA62;
defparam \Mux46~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y32_N13
dffeas \registerArray[3][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][17] .is_wysiwyg = "true";
defparam \registerArray[3][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N12
cycloneive_lcell_comb \Mux46~14 (
// Equation(s):
// \Mux46~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][17]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][17]~q )))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[3][17]~q ),
	.datad(\registerArray[1][17]~q ),
	.cin(gnd),
	.combout(\Mux46~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~14 .lut_mask = 16'hA280;
defparam \Mux46~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N2
cycloneive_lcell_comb \Mux46~15 (
// Equation(s):
// \Mux46~15_combout  = (\Mux46~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][17]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][17]~q ),
	.datad(\Mux46~14_combout ),
	.cin(gnd),
	.combout(\Mux46~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~15 .lut_mask = 16'hFF20;
defparam \Mux46~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N16
cycloneive_lcell_comb \Mux46~16 (
// Equation(s):
// \Mux46~16_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & ((\Mux46~13_combout ))) # (!\my_rf.rsel2[3]~input_o  & (\Mux46~15_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux46~15_combout ),
	.datad(\Mux46~13_combout ),
	.cin(gnd),
	.combout(\Mux46~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~16 .lut_mask = 16'hDC98;
defparam \Mux46~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y35_N25
dffeas \registerArray[13][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][17] .is_wysiwyg = "true";
defparam \registerArray[13][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y35_N3
dffeas \registerArray[12][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][17] .is_wysiwyg = "true";
defparam \registerArray[12][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N24
cycloneive_lcell_comb \Mux46~17 (
// Equation(s):
// \Mux46~17_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[13][17]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[12][17]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[13][17]~q ),
	.datad(\registerArray[12][17]~q ),
	.cin(gnd),
	.combout(\Mux46~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~17 .lut_mask = 16'hB9A8;
defparam \Mux46~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N17
dffeas \registerArray[24][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][18] .is_wysiwyg = "true";
defparam \registerArray[24][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y35_N1
dffeas \registerArray[16][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][18] .is_wysiwyg = "true";
defparam \registerArray[16][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N16
cycloneive_lcell_comb \Mux45~4 (
// Equation(s):
// \Mux45~4_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[24][18]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][18]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][18]~q ),
	.datad(\registerArray[16][18]~q ),
	.cin(gnd),
	.combout(\Mux45~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~4 .lut_mask = 16'hD9C8;
defparam \Mux45~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N5
dffeas \registerArray[10][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][18] .is_wysiwyg = "true";
defparam \registerArray[10][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y33_N31
dffeas \registerArray[8][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][18] .is_wysiwyg = "true";
defparam \registerArray[8][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N4
cycloneive_lcell_comb \Mux45~10 (
// Equation(s):
// \Mux45~10_combout  = (\my_rf.rsel2[1]~input_o  & (((\registerArray[10][18]~q ) # (\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[8][18]~q  & ((!\my_rf.rsel2[0]~input_o ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[8][18]~q ),
	.datac(\registerArray[10][18]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux45~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~10 .lut_mask = 16'hAAE4;
defparam \Mux45~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y29_N15
dffeas \registerArray[4][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][18] .is_wysiwyg = "true";
defparam \registerArray[4][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y29_N31
dffeas \registerArray[7][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][18] .is_wysiwyg = "true";
defparam \registerArray[7][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y38_N31
dffeas \registerArray[26][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][19] .is_wysiwyg = "true";
defparam \registerArray[26][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y36_N29
dffeas \registerArray[22][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][19] .is_wysiwyg = "true";
defparam \registerArray[22][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y36_N31
dffeas \registerArray[18][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][19] .is_wysiwyg = "true";
defparam \registerArray[18][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N28
cycloneive_lcell_comb \Mux44~2 (
// Equation(s):
// \Mux44~2_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[22][19]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[18][19]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[18][19]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][19]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux44~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~2 .lut_mask = 16'hCCE2;
defparam \Mux44~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y38_N9
dffeas \registerArray[30][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][19] .is_wysiwyg = "true";
defparam \registerArray[30][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y38_N30
cycloneive_lcell_comb \Mux44~3 (
// Equation(s):
// \Mux44~3_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux44~2_combout  & (\registerArray[30][19]~q )) # (!\Mux44~2_combout  & ((\registerArray[26][19]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux44~2_combout ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[30][19]~q ),
	.datac(\registerArray[26][19]~q ),
	.datad(\Mux44~2_combout ),
	.cin(gnd),
	.combout(\Mux44~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~3 .lut_mask = 16'hDDA0;
defparam \Mux44~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y35_N31
dffeas \registerArray[24][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][19] .is_wysiwyg = "true";
defparam \registerArray[24][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N4
cycloneive_lcell_comb \Mux44~4 (
// Equation(s):
// \Mux44~4_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[20][19]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[16][19]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[16][19]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[20][19]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux44~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~4 .lut_mask = 16'hCCE2;
defparam \Mux44~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N30
cycloneive_lcell_comb \Mux44~5 (
// Equation(s):
// \Mux44~5_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux44~4_combout  & (\registerArray[28][19]~q )) # (!\Mux44~4_combout  & ((\registerArray[24][19]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux44~4_combout ))))

	.dataa(\registerArray[28][19]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][19]~q ),
	.datad(\Mux44~4_combout ),
	.cin(gnd),
	.combout(\Mux44~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~5 .lut_mask = 16'hBBC0;
defparam \Mux44~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N0
cycloneive_lcell_comb \Mux44~6 (
// Equation(s):
// \Mux44~6_combout  = (\my_rf.rsel2[1]~input_o  & (((\Mux44~3_combout ) # (\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux44~5_combout  & ((!\my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux44~5_combout ),
	.datab(\Mux44~3_combout ),
	.datac(\my_rf.rsel2[1]~input_o ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux44~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~6 .lut_mask = 16'hF0CA;
defparam \Mux44~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N25
dffeas \registerArray[27][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][19] .is_wysiwyg = "true";
defparam \registerArray[27][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N11
dffeas \registerArray[19][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][19] .is_wysiwyg = "true";
defparam \registerArray[19][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N24
cycloneive_lcell_comb \Mux44~7 (
// Equation(s):
// \Mux44~7_combout  = (\my_rf.rsel2[3]~input_o  & (((\registerArray[27][19]~q ) # (\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[19][19]~q  & ((!\my_rf.rsel2[2]~input_o ))))

	.dataa(\registerArray[19][19]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][19]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux44~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~7 .lut_mask = 16'hCCE2;
defparam \Mux44~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y31_N23
dffeas \registerArray[8][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][19] .is_wysiwyg = "true";
defparam \registerArray[8][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N15
dffeas \registerArray[11][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][19] .is_wysiwyg = "true";
defparam \registerArray[11][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N31
dffeas \registerArray[1][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][19] .is_wysiwyg = "true";
defparam \registerArray[1][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N27
dffeas \registerArray[17][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][20] .is_wysiwyg = "true";
defparam \registerArray[17][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y38_N23
dffeas \registerArray[26][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][20] .is_wysiwyg = "true";
defparam \registerArray[26][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y38_N9
dffeas \registerArray[18][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][20] .is_wysiwyg = "true";
defparam \registerArray[18][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N22
cycloneive_lcell_comb \Mux43~2 (
// Equation(s):
// \Mux43~2_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & ((\registerArray[26][20]~q ))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[18][20]~q ))))

	.dataa(\registerArray[18][20]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[26][20]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux43~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~2 .lut_mask = 16'hFC22;
defparam \Mux43~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N20
cycloneive_lcell_comb \Mux43~3 (
// Equation(s):
// \Mux43~3_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux43~2_combout  & (\registerArray[30][20]~q )) # (!\Mux43~2_combout  & ((\registerArray[22][20]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux43~2_combout ))))

	.dataa(\registerArray[30][20]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][20]~q ),
	.datad(\Mux43~2_combout ),
	.cin(gnd),
	.combout(\Mux43~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~3 .lut_mask = 16'hBBC0;
defparam \Mux43~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y35_N11
dffeas \registerArray[20][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][20] .is_wysiwyg = "true";
defparam \registerArray[20][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N8
cycloneive_lcell_comb \Mux43~4 (
// Equation(s):
// \Mux43~4_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[24][20]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][20]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][20]~q ),
	.datad(\registerArray[16][20]~q ),
	.cin(gnd),
	.combout(\Mux43~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~4 .lut_mask = 16'hD9C8;
defparam \Mux43~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N10
cycloneive_lcell_comb \Mux43~5 (
// Equation(s):
// \Mux43~5_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux43~4_combout  & (\registerArray[28][20]~q )) # (!\Mux43~4_combout  & ((\registerArray[20][20]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux43~4_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[28][20]~q ),
	.datac(\registerArray[20][20]~q ),
	.datad(\Mux43~4_combout ),
	.cin(gnd),
	.combout(\Mux43~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~5 .lut_mask = 16'hDDA0;
defparam \Mux43~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N22
cycloneive_lcell_comb \Mux43~6 (
// Equation(s):
// \Mux43~6_combout  = (\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o ) # ((\Mux43~3_combout )))) # (!\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & ((\Mux43~5_combout ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux43~3_combout ),
	.datad(\Mux43~5_combout ),
	.cin(gnd),
	.combout(\Mux43~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~6 .lut_mask = 16'hB9A8;
defparam \Mux43~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y32_N25
dffeas \registerArray[3][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][20] .is_wysiwyg = "true";
defparam \registerArray[3][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y32_N27
dffeas \registerArray[1][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][20] .is_wysiwyg = "true";
defparam \registerArray[1][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N24
cycloneive_lcell_comb \Mux43~14 (
// Equation(s):
// \Mux43~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][20]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][20]~q )))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[3][20]~q ),
	.datad(\registerArray[1][20]~q ),
	.cin(gnd),
	.combout(\Mux43~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~14 .lut_mask = 16'hA280;
defparam \Mux43~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N30
cycloneive_lcell_comb \Mux43~15 (
// Equation(s):
// \Mux43~15_combout  = (\Mux43~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][20]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][20]~q ),
	.datad(\Mux43~14_combout ),
	.cin(gnd),
	.combout(\Mux43~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~15 .lut_mask = 16'hFF20;
defparam \Mux43~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y35_N21
dffeas \registerArray[13][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][20] .is_wysiwyg = "true";
defparam \registerArray[13][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y35_N23
dffeas \registerArray[12][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][20] .is_wysiwyg = "true";
defparam \registerArray[12][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N20
cycloneive_lcell_comb \Mux43~17 (
// Equation(s):
// \Mux43~17_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[13][20]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[12][20]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[12][20]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[13][20]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux43~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~17 .lut_mask = 16'hCCE2;
defparam \Mux43~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N0
cycloneive_lcell_comb \Mux43~18 (
// Equation(s):
// \Mux43~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux43~17_combout  & (\registerArray[15][20]~q )) # (!\Mux43~17_combout  & ((\registerArray[14][20]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux43~17_combout ))))

	.dataa(\registerArray[15][20]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][20]~q ),
	.datad(\Mux43~17_combout ),
	.cin(gnd),
	.combout(\Mux43~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~18 .lut_mask = 16'hBBC0;
defparam \Mux43~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X0_Y32_N24
dffeas \registerArray[21][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[21]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][21] .is_wysiwyg = "true";
defparam \registerArray[21][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N14
cycloneive_lcell_comb \Mux42~0 (
// Equation(s):
// \Mux42~0_combout  = (\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o ) # ((\registerArray[25][21]~q )))) # (!\my_rf.rsel2[3]~input_o  & (!\my_rf.rsel2[2]~input_o  & ((\registerArray[17][21]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[25][21]~q ),
	.datad(\registerArray[17][21]~q ),
	.cin(gnd),
	.combout(\Mux42~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~0 .lut_mask = 16'hB9A8;
defparam \Mux42~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N2
cycloneive_lcell_comb \Mux42~1 (
// Equation(s):
// \Mux42~1_combout  = (\Mux42~0_combout  & (((\registerArray[29][21]~q ) # (!\my_rf.rsel2[2]~input_o )))) # (!\Mux42~0_combout  & (\registerArray[21][21]~q  & (\my_rf.rsel2[2]~input_o )))

	.dataa(\registerArray[21][21]~q ),
	.datab(\Mux42~0_combout ),
	.datac(\my_rf.rsel2[2]~input_o ),
	.datad(\registerArray[29][21]~q ),
	.cin(gnd),
	.combout(\Mux42~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~1 .lut_mask = 16'hEC2C;
defparam \Mux42~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y35_N23
dffeas \registerArray[24][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][21] .is_wysiwyg = "true";
defparam \registerArray[24][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N20
cycloneive_lcell_comb \Mux42~4 (
// Equation(s):
// \Mux42~4_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[20][21]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[16][21]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[16][21]~q ),
	.datac(\registerArray[20][21]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux42~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~4 .lut_mask = 16'hAAE4;
defparam \Mux42~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N22
cycloneive_lcell_comb \Mux42~5 (
// Equation(s):
// \Mux42~5_combout  = (\Mux42~4_combout  & ((\registerArray[28][21]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux42~4_combout  & (((\registerArray[24][21]~q  & \my_rf.rsel2[3]~input_o ))))

	.dataa(\Mux42~4_combout ),
	.datab(\registerArray[28][21]~q ),
	.datac(\registerArray[24][21]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux42~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~5 .lut_mask = 16'hD8AA;
defparam \Mux42~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y39_N25
dffeas \registerArray[10][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][21] .is_wysiwyg = "true";
defparam \registerArray[10][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y39_N27
dffeas \registerArray[8][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][21] .is_wysiwyg = "true";
defparam \registerArray[8][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N24
cycloneive_lcell_comb \Mux42~12 (
// Equation(s):
// \Mux42~12_combout  = (\my_rf.rsel2[0]~input_o  & (\my_rf.rsel2[1]~input_o )) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[10][21]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[8][21]~q )))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[10][21]~q ),
	.datad(\registerArray[8][21]~q ),
	.cin(gnd),
	.combout(\Mux42~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~12 .lut_mask = 16'hD9C8;
defparam \Mux42~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N28
cycloneive_lcell_comb \Mux42~14 (
// Equation(s):
// \Mux42~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][21]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][21]~q )))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[3][21]~q ),
	.datad(\registerArray[1][21]~q ),
	.cin(gnd),
	.combout(\Mux42~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~14 .lut_mask = 16'hA280;
defparam \Mux42~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y34_N25
dffeas \registerArray[13][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][21] .is_wysiwyg = "true";
defparam \registerArray[13][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y34_N3
dffeas \registerArray[12][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][21] .is_wysiwyg = "true";
defparam \registerArray[12][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N24
cycloneive_lcell_comb \Mux42~17 (
// Equation(s):
// \Mux42~17_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[13][21]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[12][21]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[13][21]~q ),
	.datad(\registerArray[12][21]~q ),
	.cin(gnd),
	.combout(\Mux42~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~17 .lut_mask = 16'hB9A8;
defparam \Mux42~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N23
dffeas \registerArray[22][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][22] .is_wysiwyg = "true";
defparam \registerArray[22][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y38_N31
dffeas \registerArray[26][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][22] .is_wysiwyg = "true";
defparam \registerArray[26][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y38_N25
dffeas \registerArray[18][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][22] .is_wysiwyg = "true";
defparam \registerArray[18][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N30
cycloneive_lcell_comb \Mux41~2 (
// Equation(s):
// \Mux41~2_combout  = (\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o ) # ((\registerArray[26][22]~q )))) # (!\my_rf.rsel2[3]~input_o  & (!\my_rf.rsel2[2]~input_o  & ((\registerArray[18][22]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[26][22]~q ),
	.datad(\registerArray[18][22]~q ),
	.cin(gnd),
	.combout(\Mux41~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~2 .lut_mask = 16'hB9A8;
defparam \Mux41~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N21
dffeas \registerArray[30][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][22] .is_wysiwyg = "true";
defparam \registerArray[30][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N22
cycloneive_lcell_comb \Mux41~3 (
// Equation(s):
// \Mux41~3_combout  = (\Mux41~2_combout  & ((\registerArray[30][22]~q ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux41~2_combout  & (((\registerArray[22][22]~q  & \my_rf.rsel2[2]~input_o ))))

	.dataa(\Mux41~2_combout ),
	.datab(\registerArray[30][22]~q ),
	.datac(\registerArray[22][22]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux41~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~3 .lut_mask = 16'hD8AA;
defparam \Mux41~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y35_N25
dffeas \registerArray[20][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][22] .is_wysiwyg = "true";
defparam \registerArray[20][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N13
dffeas \registerArray[24][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][22] .is_wysiwyg = "true";
defparam \registerArray[24][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N23
dffeas \registerArray[16][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][22] .is_wysiwyg = "true";
defparam \registerArray[16][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N12
cycloneive_lcell_comb \Mux41~4 (
// Equation(s):
// \Mux41~4_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[24][22]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][22]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][22]~q ),
	.datad(\registerArray[16][22]~q ),
	.cin(gnd),
	.combout(\Mux41~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~4 .lut_mask = 16'hD9C8;
defparam \Mux41~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y35_N27
dffeas \registerArray[28][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][22] .is_wysiwyg = "true";
defparam \registerArray[28][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N24
cycloneive_lcell_comb \Mux41~5 (
// Equation(s):
// \Mux41~5_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux41~4_combout  & (\registerArray[28][22]~q )) # (!\Mux41~4_combout  & ((\registerArray[20][22]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux41~4_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[28][22]~q ),
	.datac(\registerArray[20][22]~q ),
	.datad(\Mux41~4_combout ),
	.cin(gnd),
	.combout(\Mux41~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~5 .lut_mask = 16'hDDA0;
defparam \Mux41~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y31_N22
cycloneive_lcell_comb \Mux41~6 (
// Equation(s):
// \Mux41~6_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o ) # (\Mux41~3_combout )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux41~5_combout  & (!\my_rf.rsel2[0]~input_o )))

	.dataa(\Mux41~5_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux41~3_combout ),
	.cin(gnd),
	.combout(\Mux41~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~6 .lut_mask = 16'hCEC2;
defparam \Mux41~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y31_N27
dffeas \registerArray[19][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][22] .is_wysiwyg = "true";
defparam \registerArray[19][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y32_N17
dffeas \registerArray[3][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][22] .is_wysiwyg = "true";
defparam \registerArray[3][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y32_N11
dffeas \registerArray[1][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][22] .is_wysiwyg = "true";
defparam \registerArray[1][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N16
cycloneive_lcell_comb \Mux41~14 (
// Equation(s):
// \Mux41~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][22]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][22]~q )))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[3][22]~q ),
	.datad(\registerArray[1][22]~q ),
	.cin(gnd),
	.combout(\Mux41~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~14 .lut_mask = 16'hA280;
defparam \Mux41~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y35_N9
dffeas \registerArray[13][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][22] .is_wysiwyg = "true";
defparam \registerArray[13][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y35_N19
dffeas \registerArray[12][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][22] .is_wysiwyg = "true";
defparam \registerArray[12][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N8
cycloneive_lcell_comb \Mux41~17 (
// Equation(s):
// \Mux41~17_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[13][22]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[12][22]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[13][22]~q ),
	.datad(\registerArray[12][22]~q ),
	.cin(gnd),
	.combout(\Mux41~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~17 .lut_mask = 16'hB9A8;
defparam \Mux41~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N27
dffeas \registerArray[25][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][23] .is_wysiwyg = "true";
defparam \registerArray[25][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N15
dffeas \registerArray[17][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][23] .is_wysiwyg = "true";
defparam \registerArray[17][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N26
cycloneive_lcell_comb \Mux40~0 (
// Equation(s):
// \Mux40~0_combout  = (\my_rf.rsel2[3]~input_o  & (((\registerArray[25][23]~q ) # (\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[17][23]~q  & ((!\my_rf.rsel2[2]~input_o ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[17][23]~q ),
	.datac(\registerArray[25][23]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux40~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~0 .lut_mask = 16'hAAE4;
defparam \Mux40~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y37_N25
dffeas \registerArray[22][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][23] .is_wysiwyg = "true";
defparam \registerArray[22][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y37_N11
dffeas \registerArray[18][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][23] .is_wysiwyg = "true";
defparam \registerArray[18][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N24
cycloneive_lcell_comb \Mux40~2 (
// Equation(s):
// \Mux40~2_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[22][23]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[18][23]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[22][23]~q ),
	.datad(\registerArray[18][23]~q ),
	.cin(gnd),
	.combout(\Mux40~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~2 .lut_mask = 16'hB9A8;
defparam \Mux40~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y37_N20
cycloneive_lcell_comb \Mux40~3 (
// Equation(s):
// \Mux40~3_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux40~2_combout  & (\registerArray[30][23]~q )) # (!\Mux40~2_combout  & ((\registerArray[26][23]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux40~2_combout ))))

	.dataa(\registerArray[30][23]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[26][23]~q ),
	.datad(\Mux40~2_combout ),
	.cin(gnd),
	.combout(\Mux40~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~3 .lut_mask = 16'hBBC0;
defparam \Mux40~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y35_N13
dffeas \registerArray[24][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][23] .is_wysiwyg = "true";
defparam \registerArray[24][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N27
dffeas \registerArray[20][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][23] .is_wysiwyg = "true";
defparam \registerArray[20][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N17
dffeas \registerArray[16][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][23] .is_wysiwyg = "true";
defparam \registerArray[16][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N26
cycloneive_lcell_comb \Mux40~4 (
// Equation(s):
// \Mux40~4_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[20][23]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][23]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[20][23]~q ),
	.datad(\registerArray[16][23]~q ),
	.cin(gnd),
	.combout(\Mux40~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~4 .lut_mask = 16'hB9A8;
defparam \Mux40~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y35_N7
dffeas \registerArray[28][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][23] .is_wysiwyg = "true";
defparam \registerArray[28][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N12
cycloneive_lcell_comb \Mux40~5 (
// Equation(s):
// \Mux40~5_combout  = (\Mux40~4_combout  & (((\registerArray[28][23]~q )) # (!\my_rf.rsel2[3]~input_o ))) # (!\Mux40~4_combout  & (\my_rf.rsel2[3]~input_o  & (\registerArray[24][23]~q )))

	.dataa(\Mux40~4_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][23]~q ),
	.datad(\registerArray[28][23]~q ),
	.cin(gnd),
	.combout(\Mux40~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~5 .lut_mask = 16'hEA62;
defparam \Mux40~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N12
cycloneive_lcell_comb \Mux40~6 (
// Equation(s):
// \Mux40~6_combout  = (\my_rf.rsel2[1]~input_o  & (((\Mux40~3_combout ) # (\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux40~5_combout  & ((!\my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux40~5_combout ),
	.datab(\Mux40~3_combout ),
	.datac(\my_rf.rsel2[1]~input_o ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux40~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~6 .lut_mask = 16'hF0CA;
defparam \Mux40~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N0
cycloneive_lcell_comb \Mux40~12 (
// Equation(s):
// \Mux40~12_combout  = (\my_rf.rsel2[0]~input_o  & (\my_rf.rsel2[1]~input_o )) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[10][23]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[8][23]~q )))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[10][23]~q ),
	.datad(\registerArray[8][23]~q ),
	.cin(gnd),
	.combout(\Mux40~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~12 .lut_mask = 16'hD9C8;
defparam \Mux40~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N24
cycloneive_lcell_comb \Mux40~13 (
// Equation(s):
// \Mux40~13_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux40~12_combout  & (\registerArray[11][23]~q )) # (!\Mux40~12_combout  & ((\registerArray[9][23]~q ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux40~12_combout ))))

	.dataa(\registerArray[11][23]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[9][23]~q ),
	.datad(\Mux40~12_combout ),
	.cin(gnd),
	.combout(\Mux40~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~13 .lut_mask = 16'hBBC0;
defparam \Mux40~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y32_N21
dffeas \registerArray[3][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][23] .is_wysiwyg = "true";
defparam \registerArray[3][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y32_N31
dffeas \registerArray[1][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][23] .is_wysiwyg = "true";
defparam \registerArray[1][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N20
cycloneive_lcell_comb \Mux40~14 (
// Equation(s):
// \Mux40~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[3][23]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[1][23]~q ))))

	.dataa(\registerArray[1][23]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[3][23]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux40~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~14 .lut_mask = 16'hE200;
defparam \Mux40~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N27
dffeas \registerArray[2][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][23] .is_wysiwyg = "true";
defparam \registerArray[2][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N26
cycloneive_lcell_comb \Mux40~15 (
// Equation(s):
// \Mux40~15_combout  = (\Mux40~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][23]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][23]~q ),
	.datad(\Mux40~14_combout ),
	.cin(gnd),
	.combout(\Mux40~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~15 .lut_mask = 16'hFF20;
defparam \Mux40~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y31_N24
cycloneive_lcell_comb \Mux40~16 (
// Equation(s):
// \Mux40~16_combout  = (\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o ) # ((\Mux40~13_combout )))) # (!\my_rf.rsel2[3]~input_o  & (!\my_rf.rsel2[2]~input_o  & ((\Mux40~15_combout ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\Mux40~13_combout ),
	.datad(\Mux40~15_combout ),
	.cin(gnd),
	.combout(\Mux40~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~16 .lut_mask = 16'hB9A8;
defparam \Mux40~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N8
cycloneive_lcell_comb \Mux39~0 (
// Equation(s):
// \Mux39~0_combout  = (\my_rf.rsel2[3]~input_o  & (\my_rf.rsel2[2]~input_o )) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\registerArray[21][24]~q )) # (!\my_rf.rsel2[2]~input_o  & ((\registerArray[17][24]~q )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[21][24]~q ),
	.datad(\registerArray[17][24]~q ),
	.cin(gnd),
	.combout(\Mux39~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~0 .lut_mask = 16'hD9C8;
defparam \Mux39~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y37_N29
dffeas \registerArray[22][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][24] .is_wysiwyg = "true";
defparam \registerArray[22][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y37_N17
dffeas \registerArray[26][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][24] .is_wysiwyg = "true";
defparam \registerArray[26][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y37_N15
dffeas \registerArray[18][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][24] .is_wysiwyg = "true";
defparam \registerArray[18][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y37_N16
cycloneive_lcell_comb \Mux39~2 (
// Equation(s):
// \Mux39~2_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[26][24]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[18][24]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[26][24]~q ),
	.datad(\registerArray[18][24]~q ),
	.cin(gnd),
	.combout(\Mux39~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~2 .lut_mask = 16'hD9C8;
defparam \Mux39~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y37_N27
dffeas \registerArray[30][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][24] .is_wysiwyg = "true";
defparam \registerArray[30][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N28
cycloneive_lcell_comb \Mux39~3 (
// Equation(s):
// \Mux39~3_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux39~2_combout  & ((\registerArray[30][24]~q ))) # (!\Mux39~2_combout  & (\registerArray[22][24]~q )))) # (!\my_rf.rsel2[2]~input_o  & (\Mux39~2_combout ))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux39~2_combout ),
	.datac(\registerArray[22][24]~q ),
	.datad(\registerArray[30][24]~q ),
	.cin(gnd),
	.combout(\Mux39~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~3 .lut_mask = 16'hEC64;
defparam \Mux39~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y35_N17
dffeas \registerArray[28][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][24] .is_wysiwyg = "true";
defparam \registerArray[28][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y31_N29
dffeas \registerArray[23][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][24] .is_wysiwyg = "true";
defparam \registerArray[23][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y31_N15
dffeas \registerArray[19][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][24] .is_wysiwyg = "true";
defparam \registerArray[19][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N28
cycloneive_lcell_comb \Mux39~7 (
// Equation(s):
// \Mux39~7_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[23][24]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[19][24]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[19][24]~q ),
	.datac(\registerArray[23][24]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux39~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~7 .lut_mask = 16'hAAE4;
defparam \Mux39~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N12
cycloneive_lcell_comb \Mux39~8 (
// Equation(s):
// \Mux39~8_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux39~7_combout  & (\registerArray[31][24]~q )) # (!\Mux39~7_combout  & ((\registerArray[27][24]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux39~7_combout ))))

	.dataa(\registerArray[31][24]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][24]~q ),
	.datad(\Mux39~7_combout ),
	.cin(gnd),
	.combout(\Mux39~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~8 .lut_mask = 16'hBBC0;
defparam \Mux39~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N27
dffeas \registerArray[8][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][24] .is_wysiwyg = "true";
defparam \registerArray[8][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N0
cycloneive_lcell_comb \Mux39~14 (
// Equation(s):
// \Mux39~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][24]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][24]~q )))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[3][24]~q ),
	.datad(\registerArray[1][24]~q ),
	.cin(gnd),
	.combout(\Mux39~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~14 .lut_mask = 16'hA280;
defparam \Mux39~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N20
cycloneive_lcell_comb \Mux39~15 (
// Equation(s):
// \Mux39~15_combout  = (\Mux39~14_combout ) # ((!\my_rf.rsel2[0]~input_o  & (\my_rf.rsel2[1]~input_o  & \registerArray[2][24]~q )))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[2][24]~q ),
	.datad(\Mux39~14_combout ),
	.cin(gnd),
	.combout(\Mux39~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~15 .lut_mask = 16'hFF40;
defparam \Mux39~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y34_N9
dffeas \registerArray[13][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][24] .is_wysiwyg = "true";
defparam \registerArray[13][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y34_N19
dffeas \registerArray[12][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][24] .is_wysiwyg = "true";
defparam \registerArray[12][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N8
cycloneive_lcell_comb \Mux39~17 (
// Equation(s):
// \Mux39~17_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[13][24]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[12][24]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[13][24]~q ),
	.datad(\registerArray[12][24]~q ),
	.cin(gnd),
	.combout(\Mux39~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~17 .lut_mask = 16'hB9A8;
defparam \Mux39~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N28
cycloneive_lcell_comb \Mux39~18 (
// Equation(s):
// \Mux39~18_combout  = (\Mux39~17_combout  & ((\registerArray[15][24]~q ) # ((!\my_rf.rsel2[1]~input_o )))) # (!\Mux39~17_combout  & (((\registerArray[14][24]~q  & \my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[15][24]~q ),
	.datab(\Mux39~17_combout ),
	.datac(\registerArray[14][24]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux39~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~18 .lut_mask = 16'hB8CC;
defparam \Mux39~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y35_N21
dffeas \registerArray[20][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][25] .is_wysiwyg = "true";
defparam \registerArray[20][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N29
dffeas \registerArray[16][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][25] .is_wysiwyg = "true";
defparam \registerArray[16][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N20
cycloneive_lcell_comb \Mux38~4 (
// Equation(s):
// \Mux38~4_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[20][25]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][25]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[20][25]~q ),
	.datad(\registerArray[16][25]~q ),
	.cin(gnd),
	.combout(\Mux38~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~4 .lut_mask = 16'hB9A8;
defparam \Mux38~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N2
cycloneive_lcell_comb \Mux38~5 (
// Equation(s):
// \Mux38~5_combout  = (\Mux38~4_combout  & (((\registerArray[28][25]~q )) # (!\my_rf.rsel2[3]~input_o ))) # (!\Mux38~4_combout  & (\my_rf.rsel2[3]~input_o  & (\registerArray[24][25]~q )))

	.dataa(\Mux38~4_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][25]~q ),
	.datad(\registerArray[28][25]~q ),
	.cin(gnd),
	.combout(\Mux38~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~5 .lut_mask = 16'hEA62;
defparam \Mux38~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N14
cycloneive_lcell_comb \Mux38~7 (
// Equation(s):
// \Mux38~7_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[27][25]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[19][25]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][25]~q ),
	.datad(\registerArray[19][25]~q ),
	.cin(gnd),
	.combout(\Mux38~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~7 .lut_mask = 16'hD9C8;
defparam \Mux38~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N30
cycloneive_lcell_comb \Mux38~8 (
// Equation(s):
// \Mux38~8_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux38~7_combout  & ((\registerArray[31][25]~q ))) # (!\Mux38~7_combout  & (\registerArray[23][25]~q )))) # (!\my_rf.rsel2[2]~input_o  & (\Mux38~7_combout ))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux38~7_combout ),
	.datac(\registerArray[23][25]~q ),
	.datad(\registerArray[31][25]~q ),
	.cin(gnd),
	.combout(\Mux38~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~8 .lut_mask = 16'hEC64;
defparam \Mux38~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N15
dffeas \registerArray[4][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][25] .is_wysiwyg = "true";
defparam \registerArray[4][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y33_N23
dffeas \registerArray[11][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][25] .is_wysiwyg = "true";
defparam \registerArray[11][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X0_Y34_N24
dffeas \registerArray[25][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[26]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][26] .is_wysiwyg = "true";
defparam \registerArray[25][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y37_N5
dffeas \registerArray[22][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][26] .is_wysiwyg = "true";
defparam \registerArray[22][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y37_N29
dffeas \registerArray[26][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][26] .is_wysiwyg = "true";
defparam \registerArray[26][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y37_N31
dffeas \registerArray[18][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][26] .is_wysiwyg = "true";
defparam \registerArray[18][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y37_N28
cycloneive_lcell_comb \Mux37~2 (
// Equation(s):
// \Mux37~2_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[26][26]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[18][26]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[26][26]~q ),
	.datad(\registerArray[18][26]~q ),
	.cin(gnd),
	.combout(\Mux37~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~2 .lut_mask = 16'hD9C8;
defparam \Mux37~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y35_N3
dffeas \registerArray[30][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][26] .is_wysiwyg = "true";
defparam \registerArray[30][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N4
cycloneive_lcell_comb \Mux37~3 (
// Equation(s):
// \Mux37~3_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux37~2_combout  & ((\registerArray[30][26]~q ))) # (!\Mux37~2_combout  & (\registerArray[22][26]~q )))) # (!\my_rf.rsel2[2]~input_o  & (\Mux37~2_combout ))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux37~2_combout ),
	.datac(\registerArray[22][26]~q ),
	.datad(\registerArray[30][26]~q ),
	.cin(gnd),
	.combout(\Mux37~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~3 .lut_mask = 16'hEC64;
defparam \Mux37~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y35_N7
dffeas \registerArray[24][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][26] .is_wysiwyg = "true";
defparam \registerArray[24][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N25
dffeas \registerArray[16][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][26] .is_wysiwyg = "true";
defparam \registerArray[16][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N6
cycloneive_lcell_comb \Mux37~4 (
// Equation(s):
// \Mux37~4_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[24][26]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][26]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][26]~q ),
	.datad(\registerArray[16][26]~q ),
	.cin(gnd),
	.combout(\Mux37~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~4 .lut_mask = 16'hD9C8;
defparam \Mux37~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N26
cycloneive_lcell_comb \Mux37~5 (
// Equation(s):
// \Mux37~5_combout  = (\Mux37~4_combout  & ((\registerArray[28][26]~q ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux37~4_combout  & (((\registerArray[20][26]~q  & \my_rf.rsel2[2]~input_o ))))

	.dataa(\Mux37~4_combout ),
	.datab(\registerArray[28][26]~q ),
	.datac(\registerArray[20][26]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux37~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~5 .lut_mask = 16'hD8AA;
defparam \Mux37~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N26
cycloneive_lcell_comb \Mux37~6 (
// Equation(s):
// \Mux37~6_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o ) # (\Mux37~3_combout )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux37~5_combout  & (!\my_rf.rsel2[0]~input_o )))

	.dataa(\Mux37~5_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux37~3_combout ),
	.cin(gnd),
	.combout(\Mux37~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~6 .lut_mask = 16'hCEC2;
defparam \Mux37~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y32_N17
dffeas \registerArray[23][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][26] .is_wysiwyg = "true";
defparam \registerArray[23][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N5
dffeas \registerArray[19][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][26] .is_wysiwyg = "true";
defparam \registerArray[19][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N16
cycloneive_lcell_comb \Mux37~7 (
// Equation(s):
// \Mux37~7_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[23][26]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[19][26]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[23][26]~q ),
	.datad(\registerArray[19][26]~q ),
	.cin(gnd),
	.combout(\Mux37~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~7 .lut_mask = 16'hB9A8;
defparam \Mux37~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y33_N9
dffeas \registerArray[9][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][26] .is_wysiwyg = "true";
defparam \registerArray[9][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y33_N9
dffeas \registerArray[10][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][26] .is_wysiwyg = "true";
defparam \registerArray[10][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y33_N19
dffeas \registerArray[8][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][26] .is_wysiwyg = "true";
defparam \registerArray[8][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N8
cycloneive_lcell_comb \Mux37~10 (
// Equation(s):
// \Mux37~10_combout  = (\my_rf.rsel2[1]~input_o  & (((\registerArray[10][26]~q ) # (\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[8][26]~q  & ((!\my_rf.rsel2[0]~input_o ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[8][26]~q ),
	.datac(\registerArray[10][26]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux37~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~10 .lut_mask = 16'hAAE4;
defparam \Mux37~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y33_N11
dffeas \registerArray[11][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][26] .is_wysiwyg = "true";
defparam \registerArray[11][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N8
cycloneive_lcell_comb \Mux37~11 (
// Equation(s):
// \Mux37~11_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux37~10_combout  & (\registerArray[11][26]~q )) # (!\Mux37~10_combout  & ((\registerArray[9][26]~q ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux37~10_combout ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\registerArray[11][26]~q ),
	.datac(\registerArray[9][26]~q ),
	.datad(\Mux37~10_combout ),
	.cin(gnd),
	.combout(\Mux37~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~11 .lut_mask = 16'hDDA0;
defparam \Mux37~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N27
dffeas \registerArray[4][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][26] .is_wysiwyg = "true";
defparam \registerArray[4][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y34_N27
dffeas \registerArray[12][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][26] .is_wysiwyg = "true";
defparam \registerArray[12][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X38_Y0_N10
dffeas \registerArray[21][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[27]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][27] .is_wysiwyg = "true";
defparam \registerArray[21][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y34_N7
dffeas \registerArray[26][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][27] .is_wysiwyg = "true";
defparam \registerArray[26][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y38_N11
dffeas \registerArray[22][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][27] .is_wysiwyg = "true";
defparam \registerArray[22][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y38_N11
dffeas \registerArray[18][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][27] .is_wysiwyg = "true";
defparam \registerArray[18][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N10
cycloneive_lcell_comb \Mux36~2 (
// Equation(s):
// \Mux36~2_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & ((\registerArray[22][27]~q ))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[18][27]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[18][27]~q ),
	.datac(\registerArray[22][27]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux36~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~2 .lut_mask = 16'hFA44;
defparam \Mux36~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y38_N29
dffeas \registerArray[30][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][27] .is_wysiwyg = "true";
defparam \registerArray[30][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N6
cycloneive_lcell_comb \Mux36~3 (
// Equation(s):
// \Mux36~3_combout  = (\Mux36~2_combout  & (((\registerArray[30][27]~q )) # (!\my_rf.rsel2[3]~input_o ))) # (!\Mux36~2_combout  & (\my_rf.rsel2[3]~input_o  & (\registerArray[26][27]~q )))

	.dataa(\Mux36~2_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[26][27]~q ),
	.datad(\registerArray[30][27]~q ),
	.cin(gnd),
	.combout(\Mux36~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~3 .lut_mask = 16'hEA62;
defparam \Mux36~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y35_N21
dffeas \registerArray[28][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][27] .is_wysiwyg = "true";
defparam \registerArray[28][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N30
cycloneive_lcell_comb \Mux36~7 (
// Equation(s):
// \Mux36~7_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[27][27]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[19][27]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][27]~q ),
	.datad(\registerArray[19][27]~q ),
	.cin(gnd),
	.combout(\Mux36~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~7 .lut_mask = 16'hD9C8;
defparam \Mux36~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N26
cycloneive_lcell_comb \Mux36~8 (
// Equation(s):
// \Mux36~8_combout  = (\Mux36~7_combout  & ((\registerArray[31][27]~q ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux36~7_combout  & (((\registerArray[23][27]~q  & \my_rf.rsel2[2]~input_o ))))

	.dataa(\Mux36~7_combout ),
	.datab(\registerArray[31][27]~q ),
	.datac(\registerArray[23][27]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux36~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~8 .lut_mask = 16'hD8AA;
defparam \Mux36~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N23
dffeas \registerArray[8][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][27] .is_wysiwyg = "true";
defparam \registerArray[8][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y33_N27
dffeas \registerArray[11][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][27] .is_wysiwyg = "true";
defparam \registerArray[11][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N4
cycloneive_lcell_comb \Mux36~17 (
// Equation(s):
// \Mux36~17_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[13][27]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[12][27]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[12][27]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[13][27]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux36~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~17 .lut_mask = 16'hCCE2;
defparam \Mux36~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N12
cycloneive_lcell_comb \Mux35~0 (
// Equation(s):
// \Mux35~0_combout  = (\my_rf.rsel2[3]~input_o  & (\my_rf.rsel2[2]~input_o )) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\registerArray[21][28]~q )) # (!\my_rf.rsel2[2]~input_o  & ((\registerArray[17][28]~q )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[21][28]~q ),
	.datad(\registerArray[17][28]~q ),
	.cin(gnd),
	.combout(\Mux35~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~0 .lut_mask = 16'hD9C8;
defparam \Mux35~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N0
cycloneive_lcell_comb \Mux35~2 (
// Equation(s):
// \Mux35~2_combout  = (\my_rf.rsel2[3]~input_o  & (((\registerArray[26][28]~q ) # (\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[18][28]~q  & ((!\my_rf.rsel2[2]~input_o ))))

	.dataa(\registerArray[18][28]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[26][28]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux35~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~2 .lut_mask = 16'hCCE2;
defparam \Mux35~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N8
cycloneive_lcell_comb \Mux35~3 (
// Equation(s):
// \Mux35~3_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux35~2_combout  & ((\registerArray[30][28]~q ))) # (!\Mux35~2_combout  & (\registerArray[22][28]~q )))) # (!\my_rf.rsel2[2]~input_o  & (\Mux35~2_combout ))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux35~2_combout ),
	.datac(\registerArray[22][28]~q ),
	.datad(\registerArray[30][28]~q ),
	.cin(gnd),
	.combout(\Mux35~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~3 .lut_mask = 16'hEC64;
defparam \Mux35~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y33_N25
dffeas \registerArray[27][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][28] .is_wysiwyg = "true";
defparam \registerArray[27][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y32_N29
dffeas \registerArray[23][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][28] .is_wysiwyg = "true";
defparam \registerArray[23][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N27
dffeas \registerArray[19][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][28] .is_wysiwyg = "true";
defparam \registerArray[19][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N28
cycloneive_lcell_comb \Mux35~7 (
// Equation(s):
// \Mux35~7_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & ((\registerArray[23][28]~q ))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[19][28]~q ))))

	.dataa(\registerArray[19][28]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[23][28]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux35~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~7 .lut_mask = 16'hFC22;
defparam \Mux35~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N15
dffeas \registerArray[31][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][28] .is_wysiwyg = "true";
defparam \registerArray[31][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N24
cycloneive_lcell_comb \Mux35~8 (
// Equation(s):
// \Mux35~8_combout  = (\Mux35~7_combout  & (((\registerArray[31][28]~q )) # (!\my_rf.rsel2[3]~input_o ))) # (!\Mux35~7_combout  & (\my_rf.rsel2[3]~input_o  & (\registerArray[27][28]~q )))

	.dataa(\Mux35~7_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][28]~q ),
	.datad(\registerArray[31][28]~q ),
	.cin(gnd),
	.combout(\Mux35~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~8 .lut_mask = 16'hEA62;
defparam \Mux35~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y34_N1
dffeas \registerArray[13][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][28] .is_wysiwyg = "true";
defparam \registerArray[13][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y34_N11
dffeas \registerArray[12][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][28] .is_wysiwyg = "true";
defparam \registerArray[12][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N0
cycloneive_lcell_comb \Mux35~17 (
// Equation(s):
// \Mux35~17_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[13][28]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[12][28]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[13][28]~q ),
	.datad(\registerArray[12][28]~q ),
	.cin(gnd),
	.combout(\Mux35~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~17 .lut_mask = 16'hB9A8;
defparam \Mux35~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N8
cycloneive_lcell_comb \Mux34~0 (
// Equation(s):
// \Mux34~0_combout  = (\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o ) # ((\registerArray[25][29]~q )))) # (!\my_rf.rsel2[3]~input_o  & (!\my_rf.rsel2[2]~input_o  & ((\registerArray[17][29]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[25][29]~q ),
	.datad(\registerArray[17][29]~q ),
	.cin(gnd),
	.combout(\Mux34~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~0 .lut_mask = 16'hB9A8;
defparam \Mux34~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N20
cycloneive_lcell_comb \Mux34~1 (
// Equation(s):
// \Mux34~1_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux34~0_combout  & ((\registerArray[29][29]~q ))) # (!\Mux34~0_combout  & (\registerArray[21][29]~q )))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux34~0_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[21][29]~q ),
	.datac(\Mux34~0_combout ),
	.datad(\registerArray[29][29]~q ),
	.cin(gnd),
	.combout(\Mux34~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~1 .lut_mask = 16'hF858;
defparam \Mux34~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y37_N13
dffeas \registerArray[22][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][29] .is_wysiwyg = "true";
defparam \registerArray[22][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y37_N7
dffeas \registerArray[18][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][29] .is_wysiwyg = "true";
defparam \registerArray[18][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N12
cycloneive_lcell_comb \Mux34~2 (
// Equation(s):
// \Mux34~2_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[22][29]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[18][29]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[22][29]~q ),
	.datad(\registerArray[18][29]~q ),
	.cin(gnd),
	.combout(\Mux34~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~2 .lut_mask = 16'hB9A8;
defparam \Mux34~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y35_N31
dffeas \registerArray[20][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][29] .is_wysiwyg = "true";
defparam \registerArray[20][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N30
cycloneive_lcell_comb \Mux34~4 (
// Equation(s):
// \Mux34~4_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[20][29]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][29]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[20][29]~q ),
	.datad(\registerArray[16][29]~q ),
	.cin(gnd),
	.combout(\Mux34~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~4 .lut_mask = 16'hB9A8;
defparam \Mux34~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N10
cycloneive_lcell_comb \Mux34~5 (
// Equation(s):
// \Mux34~5_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux34~4_combout  & (\registerArray[28][29]~q )) # (!\Mux34~4_combout  & ((\registerArray[24][29]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux34~4_combout ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[28][29]~q ),
	.datac(\registerArray[24][29]~q ),
	.datad(\Mux34~4_combout ),
	.cin(gnd),
	.combout(\Mux34~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~5 .lut_mask = 16'hDDA0;
defparam \Mux34~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N11
dffeas \registerArray[4][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][29] .is_wysiwyg = "true";
defparam \registerArray[4][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y34_N31
dffeas \registerArray[12][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][29] .is_wysiwyg = "true";
defparam \registerArray[12][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N31
dffeas \registerArray[15][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][29] .is_wysiwyg = "true";
defparam \registerArray[15][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N21
dffeas \registerArray[21][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][30] .is_wysiwyg = "true";
defparam \registerArray[21][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N15
dffeas \registerArray[17][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][30] .is_wysiwyg = "true";
defparam \registerArray[17][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N20
cycloneive_lcell_comb \Mux33~0 (
// Equation(s):
// \Mux33~0_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[21][30]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[17][30]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[17][30]~q ),
	.datac(\registerArray[21][30]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux33~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~0 .lut_mask = 16'hAAE4;
defparam \Mux33~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N18
cycloneive_lcell_comb \Mux33~1 (
// Equation(s):
// \Mux33~1_combout  = (\Mux33~0_combout  & ((\registerArray[29][30]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux33~0_combout  & (((\registerArray[25][30]~q  & \my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[29][30]~q ),
	.datab(\registerArray[25][30]~q ),
	.datac(\Mux33~0_combout ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux33~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~1 .lut_mask = 16'hACF0;
defparam \Mux33~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y38_N7
dffeas \registerArray[18][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][30] .is_wysiwyg = "true";
defparam \registerArray[18][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N27
dffeas \registerArray[24][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][30] .is_wysiwyg = "true";
defparam \registerArray[24][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N21
dffeas \registerArray[16][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][30] .is_wysiwyg = "true";
defparam \registerArray[16][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N26
cycloneive_lcell_comb \Mux33~4 (
// Equation(s):
// \Mux33~4_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[24][30]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][30]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][30]~q ),
	.datad(\registerArray[16][30]~q ),
	.cin(gnd),
	.combout(\Mux33~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~4 .lut_mask = 16'hD9C8;
defparam \Mux33~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N31
dffeas \registerArray[11][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][30] .is_wysiwyg = "true";
defparam \registerArray[11][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N27
dffeas \registerArray[5][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][30] .is_wysiwyg = "true";
defparam \registerArray[5][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N13
dffeas \registerArray[4][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][30] .is_wysiwyg = "true";
defparam \registerArray[4][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N26
cycloneive_lcell_comb \Mux33~12 (
// Equation(s):
// \Mux33~12_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[5][30]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[4][30]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[5][30]~q ),
	.datad(\registerArray[4][30]~q ),
	.cin(gnd),
	.combout(\Mux33~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~12 .lut_mask = 16'hB9A8;
defparam \Mux33~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y31_N2
cycloneive_lcell_comb \Mux33~13 (
// Equation(s):
// \Mux33~13_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux33~12_combout  & (\registerArray[7][30]~q )) # (!\Mux33~12_combout  & ((\registerArray[6][30]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux33~12_combout ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[7][30]~q ),
	.datac(\registerArray[6][30]~q ),
	.datad(\Mux33~12_combout ),
	.cin(gnd),
	.combout(\Mux33~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~13 .lut_mask = 16'hDDA0;
defparam \Mux33~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y32_N1
dffeas \registerArray[3][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][30] .is_wysiwyg = "true";
defparam \registerArray[3][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y32_N3
dffeas \registerArray[1][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][30] .is_wysiwyg = "true";
defparam \registerArray[1][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N0
cycloneive_lcell_comb \Mux33~14 (
// Equation(s):
// \Mux33~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][30]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][30]~q )))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[3][30]~q ),
	.datad(\registerArray[1][30]~q ),
	.cin(gnd),
	.combout(\Mux33~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~14 .lut_mask = 16'hA280;
defparam \Mux33~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y32_N21
dffeas \registerArray[2][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][30] .is_wysiwyg = "true";
defparam \registerArray[2][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y32_N20
cycloneive_lcell_comb \Mux33~15 (
// Equation(s):
// \Mux33~15_combout  = (\Mux33~14_combout ) # ((!\my_rf.rsel2[0]~input_o  & (\registerArray[2][30]~q  & \my_rf.rsel2[1]~input_o )))

	.dataa(\Mux33~14_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][30]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux33~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~15 .lut_mask = 16'hBAAA;
defparam \Mux33~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y32_N14
cycloneive_lcell_comb \Mux33~16 (
// Equation(s):
// \Mux33~16_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o ) # (\Mux33~13_combout )))) # (!\my_rf.rsel2[2]~input_o  & (\Mux33~15_combout  & (!\my_rf.rsel2[3]~input_o )))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux33~15_combout ),
	.datac(\my_rf.rsel2[3]~input_o ),
	.datad(\Mux33~13_combout ),
	.cin(gnd),
	.combout(\Mux33~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~16 .lut_mask = 16'hAEA4;
defparam \Mux33~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y0_N10
dffeas \registerArray[21][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[31]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][31] .is_wysiwyg = "true";
defparam \registerArray[21][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y38_N15
dffeas \registerArray[26][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][31] .is_wysiwyg = "true";
defparam \registerArray[26][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y36_N13
dffeas \registerArray[22][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][31] .is_wysiwyg = "true";
defparam \registerArray[22][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y36_N7
dffeas \registerArray[18][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][31] .is_wysiwyg = "true";
defparam \registerArray[18][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N12
cycloneive_lcell_comb \Mux32~2 (
// Equation(s):
// \Mux32~2_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[22][31]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[18][31]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[18][31]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][31]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux32~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~2 .lut_mask = 16'hCCE2;
defparam \Mux32~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y38_N9
dffeas \registerArray[30][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][31] .is_wysiwyg = "true";
defparam \registerArray[30][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N14
cycloneive_lcell_comb \Mux32~3 (
// Equation(s):
// \Mux32~3_combout  = (\Mux32~2_combout  & ((\registerArray[30][31]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux32~2_combout  & (((\registerArray[26][31]~q  & \my_rf.rsel2[3]~input_o ))))

	.dataa(\Mux32~2_combout ),
	.datab(\registerArray[30][31]~q ),
	.datac(\registerArray[26][31]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux32~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~3 .lut_mask = 16'hD8AA;
defparam \Mux32~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N16
cycloneive_lcell_comb \Mux32~4 (
// Equation(s):
// \Mux32~4_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[20][31]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][31]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[20][31]~q ),
	.datad(\registerArray[16][31]~q ),
	.cin(gnd),
	.combout(\Mux32~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~4 .lut_mask = 16'hB9A8;
defparam \Mux32~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N24
cycloneive_lcell_comb \Mux32~5 (
// Equation(s):
// \Mux32~5_combout  = (\Mux32~4_combout  & (((\registerArray[28][31]~q )) # (!\my_rf.rsel2[3]~input_o ))) # (!\Mux32~4_combout  & (\my_rf.rsel2[3]~input_o  & (\registerArray[24][31]~q )))

	.dataa(\Mux32~4_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][31]~q ),
	.datad(\registerArray[28][31]~q ),
	.cin(gnd),
	.combout(\Mux32~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~5 .lut_mask = 16'hEA62;
defparam \Mux32~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N6
cycloneive_lcell_comb \Mux32~6 (
// Equation(s):
// \Mux32~6_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux32~3_combout ) # ((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (((!\my_rf.rsel2[0]~input_o  & \Mux32~5_combout ))))

	.dataa(\Mux32~3_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux32~5_combout ),
	.cin(gnd),
	.combout(\Mux32~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~6 .lut_mask = 16'hCBC8;
defparam \Mux32~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N29
dffeas \registerArray[27][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][31] .is_wysiwyg = "true";
defparam \registerArray[27][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N7
dffeas \registerArray[19][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][31] .is_wysiwyg = "true";
defparam \registerArray[19][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N28
cycloneive_lcell_comb \Mux32~7 (
// Equation(s):
// \Mux32~7_combout  = (\my_rf.rsel2[3]~input_o  & (((\registerArray[27][31]~q ) # (\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[19][31]~q  & ((!\my_rf.rsel2[2]~input_o ))))

	.dataa(\registerArray[19][31]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][31]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux32~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~7 .lut_mask = 16'hCCE2;
defparam \Mux32~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N12
cycloneive_lcell_comb \Mux32~10 (
// Equation(s):
// \Mux32~10_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & ((\registerArray[5][31]~q ))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][31]~q ))))

	.dataa(\registerArray[4][31]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[5][31]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux32~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~10 .lut_mask = 16'hFC22;
defparam \Mux32~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N10
cycloneive_lcell_comb \Mux32~11 (
// Equation(s):
// \Mux32~11_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux32~10_combout  & ((\registerArray[7][31]~q ))) # (!\Mux32~10_combout  & (\registerArray[6][31]~q )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux32~10_combout ))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux32~10_combout ),
	.datac(\registerArray[6][31]~q ),
	.datad(\registerArray[7][31]~q ),
	.cin(gnd),
	.combout(\Mux32~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~11 .lut_mask = 16'hEC64;
defparam \Mux32~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y37_N13
dffeas \registerArray[9][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][31] .is_wysiwyg = "true";
defparam \registerArray[9][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y37_N13
dffeas \registerArray[10][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][31] .is_wysiwyg = "true";
defparam \registerArray[10][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y37_N23
dffeas \registerArray[8][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][31] .is_wysiwyg = "true";
defparam \registerArray[8][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y37_N12
cycloneive_lcell_comb \Mux32~12 (
// Equation(s):
// \Mux32~12_combout  = (\my_rf.rsel2[0]~input_o  & (((\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[10][31]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[8][31]~q ))))

	.dataa(\registerArray[8][31]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[10][31]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux32~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~12 .lut_mask = 16'hFC22;
defparam \Mux32~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y37_N23
dffeas \registerArray[11][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][31] .is_wysiwyg = "true";
defparam \registerArray[11][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y37_N12
cycloneive_lcell_comb \Mux32~13 (
// Equation(s):
// \Mux32~13_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux32~12_combout  & (\registerArray[11][31]~q )) # (!\Mux32~12_combout  & ((\registerArray[9][31]~q ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux32~12_combout ))))

	.dataa(\registerArray[11][31]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[9][31]~q ),
	.datad(\Mux32~12_combout ),
	.cin(gnd),
	.combout(\Mux32~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~13 .lut_mask = 16'hBBC0;
defparam \Mux32~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y36_N31
dffeas \registerArray[1][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][31] .is_wysiwyg = "true";
defparam \registerArray[1][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y36_N13
dffeas \registerArray[15][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][31] .is_wysiwyg = "true";
defparam \registerArray[15][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N2
cycloneive_lcell_comb \Mux31~0 (
// Equation(s):
// \Mux31~0_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[21][0]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[17][0]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[17][0]~q ),
	.datad(\registerArray[21][0]~q ),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~0 .lut_mask = 16'hDC98;
defparam \Mux31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N24
cycloneive_lcell_comb \Mux31~1 (
// Equation(s):
// \Mux31~1_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux31~0_combout  & ((\registerArray[29][0]~q ))) # (!\Mux31~0_combout  & (\registerArray[25][0]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux31~0_combout ))))

	.dataa(\registerArray[25][0]~q ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[29][0]~q ),
	.datad(\Mux31~0_combout ),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~1 .lut_mask = 16'hF388;
defparam \Mux31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N18
cycloneive_lcell_comb \Mux31~2 (
// Equation(s):
// \Mux31~2_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[26][0]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[18][0]~q )))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[26][0]~q ),
	.datac(\registerArray[18][0]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux31~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~2 .lut_mask = 16'hEE50;
defparam \Mux31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y38_N16
cycloneive_lcell_comb \Mux31~3 (
// Equation(s):
// \Mux31~3_combout  = (\Mux31~2_combout  & (((\registerArray[30][0]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux31~2_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[22][0]~q ))))

	.dataa(\Mux31~2_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[30][0]~q ),
	.datad(\registerArray[22][0]~q ),
	.cin(gnd),
	.combout(\Mux31~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~3 .lut_mask = 16'hE6A2;
defparam \Mux31~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N26
cycloneive_lcell_comb \Mux31~4 (
// Equation(s):
// \Mux31~4_combout  = (\my_rf.rsel1[2]~input_o  & (\my_rf.rsel1[3]~input_o )) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & ((\registerArray[24][0]~q ))) # (!\my_rf.rsel1[3]~input_o  & (\registerArray[16][0]~q ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[16][0]~q ),
	.datad(\registerArray[24][0]~q ),
	.cin(gnd),
	.combout(\Mux31~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~4 .lut_mask = 16'hDC98;
defparam \Mux31~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N2
cycloneive_lcell_comb \Mux31~7 (
// Equation(s):
// \Mux31~7_combout  = (\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o ) # ((\registerArray[23][0]~q )))) # (!\my_rf.rsel1[2]~input_o  & (!\my_rf.rsel1[3]~input_o  & (\registerArray[19][0]~q )))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[19][0]~q ),
	.datad(\registerArray[23][0]~q ),
	.cin(gnd),
	.combout(\Mux31~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~7 .lut_mask = 16'hBA98;
defparam \Mux31~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N10
cycloneive_lcell_comb \Mux31~10 (
// Equation(s):
// \Mux31~10_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\registerArray[10][0]~q )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & (\registerArray[8][0]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[8][0]~q ),
	.datad(\registerArray[10][0]~q ),
	.cin(gnd),
	.combout(\Mux31~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~10 .lut_mask = 16'hBA98;
defparam \Mux31~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N10
cycloneive_lcell_comb \Mux31~12 (
// Equation(s):
// \Mux31~12_combout  = (\my_rf.rsel1[0]~input_o  & ((\registerArray[5][0]~q ) # ((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & (((\registerArray[4][0]~q  & !\my_rf.rsel1[1]~input_o ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\registerArray[5][0]~q ),
	.datac(\registerArray[4][0]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux31~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~12 .lut_mask = 16'hAAD8;
defparam \Mux31~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N2
cycloneive_lcell_comb \Mux31~13 (
// Equation(s):
// \Mux31~13_combout  = (\Mux31~12_combout  & (((\registerArray[7][0]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux31~12_combout  & (\registerArray[6][0]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux31~12_combout ),
	.datab(\registerArray[6][0]~q ),
	.datac(\registerArray[7][0]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux31~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~13 .lut_mask = 16'hE4AA;
defparam \Mux31~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N2
cycloneive_lcell_comb \Mux31~14 (
// Equation(s):
// \Mux31~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][0]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][0]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[1][0]~q ),
	.datad(\registerArray[3][0]~q ),
	.cin(gnd),
	.combout(\Mux31~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~14 .lut_mask = 16'hA820;
defparam \Mux31~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N20
cycloneive_lcell_comb \Mux31~15 (
// Equation(s):
// \Mux31~15_combout  = (\Mux31~14_combout ) # ((!\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o  & \registerArray[2][0]~q )))

	.dataa(\Mux31~14_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\registerArray[2][0]~q ),
	.cin(gnd),
	.combout(\Mux31~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~15 .lut_mask = 16'hBAAA;
defparam \Mux31~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N22
cycloneive_lcell_comb \Mux31~16 (
// Equation(s):
// \Mux31~16_combout  = (\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o ) # ((\Mux31~13_combout )))) # (!\my_rf.rsel1[2]~input_o  & (!\my_rf.rsel1[3]~input_o  & ((\Mux31~15_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\Mux31~13_combout ),
	.datad(\Mux31~15_combout ),
	.cin(gnd),
	.combout(\Mux31~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~16 .lut_mask = 16'hB9A8;
defparam \Mux31~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N2
cycloneive_lcell_comb \Mux31~17 (
// Equation(s):
// \Mux31~17_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[13][0]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[12][0]~q )))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[13][0]~q ),
	.datac(\registerArray[12][0]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux31~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~17 .lut_mask = 16'hEE50;
defparam \Mux31~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N2
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// \Mux30~0_combout  = (\my_rf.rsel1[2]~input_o  & (\my_rf.rsel1[3]~input_o )) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & ((\registerArray[25][1]~q ))) # (!\my_rf.rsel1[3]~input_o  & (\registerArray[17][1]~q ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[17][1]~q ),
	.datad(\registerArray[25][1]~q ),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'hDC98;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N24
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// \Mux30~1_combout  = (\Mux30~0_combout  & (((\registerArray[29][1]~q ) # (!\my_rf.rsel1[2]~input_o )))) # (!\Mux30~0_combout  & (\registerArray[21][1]~q  & ((\my_rf.rsel1[2]~input_o ))))

	.dataa(\Mux30~0_combout ),
	.datab(\registerArray[21][1]~q ),
	.datac(\registerArray[29][1]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'hE4AA;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N26
cycloneive_lcell_comb \Mux30~2 (
// Equation(s):
// \Mux30~2_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[22][1]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][1]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][1]~q ),
	.datad(\registerArray[22][1]~q ),
	.cin(gnd),
	.combout(\Mux30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~2 .lut_mask = 16'hDC98;
defparam \Mux30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N2
cycloneive_lcell_comb \Mux30~4 (
// Equation(s):
// \Mux30~4_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[20][1]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[16][1]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[16][1]~q ),
	.datad(\registerArray[20][1]~q ),
	.cin(gnd),
	.combout(\Mux30~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~4 .lut_mask = 16'hDC98;
defparam \Mux30~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N18
cycloneive_lcell_comb \Mux30~5 (
// Equation(s):
// \Mux30~5_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux30~4_combout  & ((\registerArray[28][1]~q ))) # (!\Mux30~4_combout  & (\registerArray[24][1]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux30~4_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[24][1]~q ),
	.datac(\registerArray[28][1]~q ),
	.datad(\Mux30~4_combout ),
	.cin(gnd),
	.combout(\Mux30~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~5 .lut_mask = 16'hF588;
defparam \Mux30~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N6
cycloneive_lcell_comb \Mux30~7 (
// Equation(s):
// \Mux30~7_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[27][1]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[19][1]~q )))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[27][1]~q ),
	.datac(\registerArray[19][1]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux30~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~7 .lut_mask = 16'hEE50;
defparam \Mux30~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N6
cycloneive_lcell_comb \Mux30~12 (
// Equation(s):
// \Mux30~12_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\registerArray[10][1]~q )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & (\registerArray[8][1]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[8][1]~q ),
	.datad(\registerArray[10][1]~q ),
	.cin(gnd),
	.combout(\Mux30~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~12 .lut_mask = 16'hBA98;
defparam \Mux30~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N30
cycloneive_lcell_comb \Mux30~13 (
// Equation(s):
// \Mux30~13_combout  = (\Mux30~12_combout  & (((\registerArray[11][1]~q )) # (!\my_rf.rsel1[0]~input_o ))) # (!\Mux30~12_combout  & (\my_rf.rsel1[0]~input_o  & ((\registerArray[9][1]~q ))))

	.dataa(\Mux30~12_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[11][1]~q ),
	.datad(\registerArray[9][1]~q ),
	.cin(gnd),
	.combout(\Mux30~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~13 .lut_mask = 16'hE6A2;
defparam \Mux30~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N6
cycloneive_lcell_comb \Mux30~14 (
// Equation(s):
// \Mux30~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][1]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][1]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[1][1]~q ),
	.datad(\registerArray[3][1]~q ),
	.cin(gnd),
	.combout(\Mux30~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~14 .lut_mask = 16'hA820;
defparam \Mux30~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N24
cycloneive_lcell_comb \Mux30~15 (
// Equation(s):
// \Mux30~15_combout  = (\Mux30~14_combout ) # ((\registerArray[2][1]~q  & (!\my_rf.rsel1[0]~input_o  & \my_rf.rsel1[1]~input_o )))

	.dataa(\registerArray[2][1]~q ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\Mux30~14_combout ),
	.cin(gnd),
	.combout(\Mux30~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~15 .lut_mask = 16'hFF20;
defparam \Mux30~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N26
cycloneive_lcell_comb \Mux30~16 (
// Equation(s):
// \Mux30~16_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux30~13_combout ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((!\my_rf.rsel1[2]~input_o  & \Mux30~15_combout ))))

	.dataa(\Mux30~13_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux30~15_combout ),
	.cin(gnd),
	.combout(\Mux30~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~16 .lut_mask = 16'hCBC8;
defparam \Mux30~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N28
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[21][2]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[17][2]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[17][2]~q ),
	.datad(\registerArray[21][2]~q ),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'hDC98;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N4
cycloneive_lcell_comb \Mux29~2 (
// Equation(s):
// \Mux29~2_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[26][2]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[18][2]~q )))))

	.dataa(\registerArray[26][2]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][2]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux29~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~2 .lut_mask = 16'hEE30;
defparam \Mux29~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N2
cycloneive_lcell_comb \Mux29~3 (
// Equation(s):
// \Mux29~3_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux29~2_combout  & (\registerArray[30][2]~q )) # (!\Mux29~2_combout  & ((\registerArray[22][2]~q ))))) # (!\my_rf.rsel1[2]~input_o  & (\Mux29~2_combout ))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux29~2_combout ),
	.datac(\registerArray[30][2]~q ),
	.datad(\registerArray[22][2]~q ),
	.cin(gnd),
	.combout(\Mux29~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~3 .lut_mask = 16'hE6C4;
defparam \Mux29~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N18
cycloneive_lcell_comb \Mux29~7 (
// Equation(s):
// \Mux29~7_combout  = (\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o ) # ((\registerArray[23][2]~q )))) # (!\my_rf.rsel1[2]~input_o  & (!\my_rf.rsel1[3]~input_o  & (\registerArray[19][2]~q )))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[19][2]~q ),
	.datad(\registerArray[23][2]~q ),
	.cin(gnd),
	.combout(\Mux29~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~7 .lut_mask = 16'hBA98;
defparam \Mux29~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N18
cycloneive_lcell_comb \Mux29~8 (
// Equation(s):
// \Mux29~8_combout  = (\Mux29~7_combout  & (((\registerArray[31][2]~q ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux29~7_combout  & (\registerArray[27][2]~q  & ((\my_rf.rsel1[3]~input_o ))))

	.dataa(\Mux29~7_combout ),
	.datab(\registerArray[27][2]~q ),
	.datac(\registerArray[31][2]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux29~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~8 .lut_mask = 16'hE4AA;
defparam \Mux29~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N2
cycloneive_lcell_comb \Mux29~10 (
// Equation(s):
// \Mux29~10_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\registerArray[10][2]~q )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & (\registerArray[8][2]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[8][2]~q ),
	.datad(\registerArray[10][2]~q ),
	.cin(gnd),
	.combout(\Mux29~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~10 .lut_mask = 16'hBA98;
defparam \Mux29~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N18
cycloneive_lcell_comb \Mux29~12 (
// Equation(s):
// \Mux29~12_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o ) # ((\registerArray[5][2]~q )))) # (!\my_rf.rsel1[0]~input_o  & (!\my_rf.rsel1[1]~input_o  & (\registerArray[4][2]~q )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[4][2]~q ),
	.datad(\registerArray[5][2]~q ),
	.cin(gnd),
	.combout(\Mux29~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~12 .lut_mask = 16'hBA98;
defparam \Mux29~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N26
cycloneive_lcell_comb \Mux29~13 (
// Equation(s):
// \Mux29~13_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux29~12_combout  & ((\registerArray[7][2]~q ))) # (!\Mux29~12_combout  & (\registerArray[6][2]~q )))) # (!\my_rf.rsel1[1]~input_o  & (((\Mux29~12_combout ))))

	.dataa(\registerArray[6][2]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[7][2]~q ),
	.datad(\Mux29~12_combout ),
	.cin(gnd),
	.combout(\Mux29~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~13 .lut_mask = 16'hF388;
defparam \Mux29~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N26
cycloneive_lcell_comb \Mux29~14 (
// Equation(s):
// \Mux29~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][2]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][2]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[1][2]~q ),
	.datad(\registerArray[3][2]~q ),
	.cin(gnd),
	.combout(\Mux29~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~14 .lut_mask = 16'hA820;
defparam \Mux29~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N4
cycloneive_lcell_comb \Mux29~15 (
// Equation(s):
// \Mux29~15_combout  = (\Mux29~14_combout ) # ((!\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o  & \registerArray[2][2]~q )))

	.dataa(\Mux29~14_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\registerArray[2][2]~q ),
	.cin(gnd),
	.combout(\Mux29~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~15 .lut_mask = 16'hBAAA;
defparam \Mux29~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N22
cycloneive_lcell_comb \Mux29~16 (
// Equation(s):
// \Mux29~16_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & (\Mux29~13_combout )) # (!\my_rf.rsel1[2]~input_o  & ((\Mux29~15_combout )))))

	.dataa(\Mux29~13_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\Mux29~15_combout ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux29~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~16 .lut_mask = 16'hEE30;
defparam \Mux29~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N26
cycloneive_lcell_comb \Mux29~17 (
// Equation(s):
// \Mux29~17_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[13][2]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[12][2]~q )))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[13][2]~q ),
	.datac(\registerArray[12][2]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux29~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~17 .lut_mask = 16'hEE50;
defparam \Mux29~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N6
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[25][3]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[17][3]~q )))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[25][3]~q ),
	.datac(\registerArray[17][3]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'hEE50;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N8
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// \Mux28~1_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux28~0_combout  & ((\registerArray[29][3]~q ))) # (!\Mux28~0_combout  & (\registerArray[21][3]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux28~0_combout ))))

	.dataa(\registerArray[21][3]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[29][3]~q ),
	.datad(\Mux28~0_combout ),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hF388;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N14
cycloneive_lcell_comb \Mux28~2 (
// Equation(s):
// \Mux28~2_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[22][3]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][3]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][3]~q ),
	.datad(\registerArray[22][3]~q ),
	.cin(gnd),
	.combout(\Mux28~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~2 .lut_mask = 16'hDC98;
defparam \Mux28~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N30
cycloneive_lcell_comb \Mux28~4 (
// Equation(s):
// \Mux28~4_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[20][3]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[16][3]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[16][3]~q ),
	.datad(\registerArray[20][3]~q ),
	.cin(gnd),
	.combout(\Mux28~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~4 .lut_mask = 16'hDC98;
defparam \Mux28~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N30
cycloneive_lcell_comb \Mux28~7 (
// Equation(s):
// \Mux28~7_combout  = (\my_rf.rsel1[2]~input_o  & (\my_rf.rsel1[3]~input_o )) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & ((\registerArray[27][3]~q ))) # (!\my_rf.rsel1[3]~input_o  & (\registerArray[19][3]~q ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[19][3]~q ),
	.datad(\registerArray[27][3]~q ),
	.cin(gnd),
	.combout(\Mux28~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~7 .lut_mask = 16'hDC98;
defparam \Mux28~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N30
cycloneive_lcell_comb \Mux28~12 (
// Equation(s):
// \Mux28~12_combout  = (\my_rf.rsel1[1]~input_o  & ((\registerArray[10][3]~q ) # ((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & (((\registerArray[8][3]~q  & !\my_rf.rsel1[0]~input_o ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[10][3]~q ),
	.datac(\registerArray[8][3]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux28~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~12 .lut_mask = 16'hAAD8;
defparam \Mux28~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N22
cycloneive_lcell_comb \Mux28~13 (
// Equation(s):
// \Mux28~13_combout  = (\Mux28~12_combout  & (((\registerArray[11][3]~q ) # (!\my_rf.rsel1[0]~input_o )))) # (!\Mux28~12_combout  & (\registerArray[9][3]~q  & ((\my_rf.rsel1[0]~input_o ))))

	.dataa(\Mux28~12_combout ),
	.datab(\registerArray[9][3]~q ),
	.datac(\registerArray[11][3]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux28~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~13 .lut_mask = 16'hE4AA;
defparam \Mux28~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N22
cycloneive_lcell_comb \Mux28~14 (
// Equation(s):
// \Mux28~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][3]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][3]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[1][3]~q ),
	.datad(\registerArray[3][3]~q ),
	.cin(gnd),
	.combout(\Mux28~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~14 .lut_mask = 16'hA820;
defparam \Mux28~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N14
cycloneive_lcell_comb \Mux28~17 (
// Equation(s):
// \Mux28~17_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[13][3]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[12][3]~q )))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[13][3]~q ),
	.datac(\registerArray[12][3]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux28~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~17 .lut_mask = 16'hEE50;
defparam \Mux28~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N10
cycloneive_lcell_comb \Mux27~2 (
// Equation(s):
// \Mux27~2_combout  = (\my_rf.rsel1[3]~input_o  & ((\registerArray[26][4]~q ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((\registerArray[18][4]~q  & !\my_rf.rsel1[2]~input_o ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[26][4]~q ),
	.datac(\registerArray[18][4]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux27~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~2 .lut_mask = 16'hAAD8;
defparam \Mux27~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N10
cycloneive_lcell_comb \Mux27~3 (
// Equation(s):
// \Mux27~3_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux27~2_combout  & ((\registerArray[30][4]~q ))) # (!\Mux27~2_combout  & (\registerArray[22][4]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux27~2_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[22][4]~q ),
	.datac(\registerArray[30][4]~q ),
	.datad(\Mux27~2_combout ),
	.cin(gnd),
	.combout(\Mux27~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~3 .lut_mask = 16'hF588;
defparam \Mux27~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N26
cycloneive_lcell_comb \Mux27~12 (
// Equation(s):
// \Mux27~12_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o ) # ((\registerArray[5][4]~q )))) # (!\my_rf.rsel1[0]~input_o  & (!\my_rf.rsel1[1]~input_o  & (\registerArray[4][4]~q )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[4][4]~q ),
	.datad(\registerArray[5][4]~q ),
	.cin(gnd),
	.combout(\Mux27~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~12 .lut_mask = 16'hBA98;
defparam \Mux27~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N18
cycloneive_lcell_comb \Mux27~13 (
// Equation(s):
// \Mux27~13_combout  = (\Mux27~12_combout  & (((\registerArray[7][4]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux27~12_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[6][4]~q ))))

	.dataa(\Mux27~12_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[7][4]~q ),
	.datad(\registerArray[6][4]~q ),
	.cin(gnd),
	.combout(\Mux27~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~13 .lut_mask = 16'hE6A2;
defparam \Mux27~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N18
cycloneive_lcell_comb \Mux27~17 (
// Equation(s):
// \Mux27~17_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[13][4]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[12][4]~q )))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[13][4]~q ),
	.datac(\registerArray[12][4]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux27~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~17 .lut_mask = 16'hEE50;
defparam \Mux27~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N2
cycloneive_lcell_comb \Mux27~18 (
// Equation(s):
// \Mux27~18_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux27~17_combout  & ((\registerArray[15][4]~q ))) # (!\Mux27~17_combout  & (\registerArray[14][4]~q )))) # (!\my_rf.rsel1[1]~input_o  & (((\Mux27~17_combout ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[14][4]~q ),
	.datac(\registerArray[15][4]~q ),
	.datad(\Mux27~17_combout ),
	.cin(gnd),
	.combout(\Mux27~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~18 .lut_mask = 16'hF588;
defparam \Mux27~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N22
cycloneive_lcell_comb \Mux26~2 (
// Equation(s):
// \Mux26~2_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[22][5]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][5]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][5]~q ),
	.datad(\registerArray[22][5]~q ),
	.cin(gnd),
	.combout(\Mux26~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~2 .lut_mask = 16'hDC98;
defparam \Mux26~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N6
cycloneive_lcell_comb \Mux26~10 (
// Equation(s):
// \Mux26~10_combout  = (\my_rf.rsel1[0]~input_o  & ((\registerArray[5][5]~q ) # ((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & (((\registerArray[4][5]~q  & !\my_rf.rsel1[1]~input_o ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\registerArray[5][5]~q ),
	.datac(\registerArray[4][5]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux26~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~10 .lut_mask = 16'hAAD8;
defparam \Mux26~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N8
cycloneive_lcell_comb \Mux25~7 (
// Equation(s):
// \Mux25~7_combout  = (\my_rf.rsel1[2]~input_o  & ((\registerArray[23][6]~q ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\registerArray[19][6]~q  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\registerArray[23][6]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[19][6]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux25~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~7 .lut_mask = 16'hCCB8;
defparam \Mux25~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N26
cycloneive_lcell_comb \Mux25~8 (
// Equation(s):
// \Mux25~8_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux25~7_combout  & (\registerArray[31][6]~q )) # (!\Mux25~7_combout  & ((\registerArray[27][6]~q ))))) # (!\my_rf.rsel1[3]~input_o  & (\Mux25~7_combout ))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux25~7_combout ),
	.datac(\registerArray[31][6]~q ),
	.datad(\registerArray[27][6]~q ),
	.cin(gnd),
	.combout(\Mux25~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~8 .lut_mask = 16'hE6C4;
defparam \Mux25~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N2
cycloneive_lcell_comb \Mux25~12 (
// Equation(s):
// \Mux25~12_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o ) # ((\registerArray[5][6]~q )))) # (!\my_rf.rsel1[0]~input_o  & (!\my_rf.rsel1[1]~input_o  & (\registerArray[4][6]~q )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[4][6]~q ),
	.datad(\registerArray[5][6]~q ),
	.cin(gnd),
	.combout(\Mux25~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~12 .lut_mask = 16'hBA98;
defparam \Mux25~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N24
cycloneive_lcell_comb \Mux25~13 (
// Equation(s):
// \Mux25~13_combout  = (\Mux25~12_combout  & (((\registerArray[7][6]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux25~12_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[6][6]~q ))))

	.dataa(\Mux25~12_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[7][6]~q ),
	.datad(\registerArray[6][6]~q ),
	.cin(gnd),
	.combout(\Mux25~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~13 .lut_mask = 16'hE6A2;
defparam \Mux25~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N18
cycloneive_lcell_comb \Mux25~14 (
// Equation(s):
// \Mux25~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][6]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][6]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[1][6]~q ),
	.datad(\registerArray[3][6]~q ),
	.cin(gnd),
	.combout(\Mux25~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~14 .lut_mask = 16'hA820;
defparam \Mux25~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N4
cycloneive_lcell_comb \Mux25~15 (
// Equation(s):
// \Mux25~15_combout  = (\Mux25~14_combout ) # ((\my_rf.rsel1[1]~input_o  & (\registerArray[2][6]~q  & !\my_rf.rsel1[0]~input_o )))

	.dataa(\Mux25~14_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[2][6]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux25~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~15 .lut_mask = 16'hAAEA;
defparam \Mux25~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N30
cycloneive_lcell_comb \Mux25~16 (
// Equation(s):
// \Mux25~16_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\Mux25~13_combout ))) # (!\my_rf.rsel1[2]~input_o  & (\Mux25~15_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux25~15_combout ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux25~13_combout ),
	.cin(gnd),
	.combout(\Mux25~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~16 .lut_mask = 16'hF4A4;
defparam \Mux25~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N0
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[25][7]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[17][7]~q )))))

	.dataa(\registerArray[25][7]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[17][7]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'hEE30;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N6
cycloneive_lcell_comb \Mux24~2 (
// Equation(s):
// \Mux24~2_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & (\registerArray[22][7]~q )) # (!\my_rf.rsel1[2]~input_o  & ((\registerArray[18][7]~q )))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[22][7]~q ),
	.datac(\registerArray[18][7]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux24~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~2 .lut_mask = 16'hEE50;
defparam \Mux24~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N14
cycloneive_lcell_comb \Mux24~3 (
// Equation(s):
// \Mux24~3_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux24~2_combout  & ((\registerArray[30][7]~q ))) # (!\Mux24~2_combout  & (\registerArray[26][7]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux24~2_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[26][7]~q ),
	.datac(\registerArray[30][7]~q ),
	.datad(\Mux24~2_combout ),
	.cin(gnd),
	.combout(\Mux24~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~3 .lut_mask = 16'hF588;
defparam \Mux24~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N10
cycloneive_lcell_comb \Mux24~4 (
// Equation(s):
// \Mux24~4_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & (\registerArray[20][7]~q )) # (!\my_rf.rsel1[2]~input_o  & ((\registerArray[16][7]~q )))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[20][7]~q ),
	.datac(\registerArray[16][7]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux24~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~4 .lut_mask = 16'hEE50;
defparam \Mux24~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N22
cycloneive_lcell_comb \Mux24~5 (
// Equation(s):
// \Mux24~5_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux24~4_combout  & ((\registerArray[28][7]~q ))) # (!\Mux24~4_combout  & (\registerArray[24][7]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux24~4_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[24][7]~q ),
	.datac(\registerArray[28][7]~q ),
	.datad(\Mux24~4_combout ),
	.cin(gnd),
	.combout(\Mux24~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~5 .lut_mask = 16'hF588;
defparam \Mux24~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N20
cycloneive_lcell_comb \Mux24~6 (
// Equation(s):
// \Mux24~6_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\Mux24~3_combout )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & ((\Mux24~5_combout ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux24~3_combout ),
	.datad(\Mux24~5_combout ),
	.cin(gnd),
	.combout(\Mux24~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~6 .lut_mask = 16'hB9A8;
defparam \Mux24~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N8
cycloneive_lcell_comb \Mux24~10 (
// Equation(s):
// \Mux24~10_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[5][7]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[4][7]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[4][7]~q ),
	.datad(\registerArray[5][7]~q ),
	.cin(gnd),
	.combout(\Mux24~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~10 .lut_mask = 16'hDC98;
defparam \Mux24~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N10
cycloneive_lcell_comb \Mux24~12 (
// Equation(s):
// \Mux24~12_combout  = (\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o )) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[10][7]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[8][7]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[8][7]~q ),
	.datad(\registerArray[10][7]~q ),
	.cin(gnd),
	.combout(\Mux24~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~12 .lut_mask = 16'hDC98;
defparam \Mux24~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N28
cycloneive_lcell_comb \Mux24~17 (
// Equation(s):
// \Mux24~17_combout  = (\my_rf.rsel1[0]~input_o  & ((\registerArray[13][7]~q ) # ((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & (((\registerArray[12][7]~q  & !\my_rf.rsel1[1]~input_o ))))

	.dataa(\registerArray[13][7]~q ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][7]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux24~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~17 .lut_mask = 16'hCCB8;
defparam \Mux24~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N10
cycloneive_lcell_comb \Mux24~18 (
// Equation(s):
// \Mux24~18_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux24~17_combout  & (\registerArray[15][7]~q )) # (!\Mux24~17_combout  & ((\registerArray[14][7]~q ))))) # (!\my_rf.rsel1[1]~input_o  & (\Mux24~17_combout ))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\Mux24~17_combout ),
	.datac(\registerArray[15][7]~q ),
	.datad(\registerArray[14][7]~q ),
	.cin(gnd),
	.combout(\Mux24~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~18 .lut_mask = 16'hE6C4;
defparam \Mux24~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y37_N26
cycloneive_lcell_comb \Mux23~10 (
// Equation(s):
// \Mux23~10_combout  = (\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o )) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[10][8]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[8][8]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[8][8]~q ),
	.datad(\registerArray[10][8]~q ),
	.cin(gnd),
	.combout(\Mux23~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~10 .lut_mask = 16'hDC98;
defparam \Mux23~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N16
cycloneive_lcell_comb \Mux23~12 (
// Equation(s):
// \Mux23~12_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[5][8]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[4][8]~q )))))

	.dataa(\registerArray[5][8]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[4][8]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux23~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~12 .lut_mask = 16'hEE30;
defparam \Mux23~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N10
cycloneive_lcell_comb \Mux23~17 (
// Equation(s):
// \Mux23~17_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o ) # ((\registerArray[13][8]~q )))) # (!\my_rf.rsel1[0]~input_o  & (!\my_rf.rsel1[1]~input_o  & (\registerArray[12][8]~q )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[12][8]~q ),
	.datad(\registerArray[13][8]~q ),
	.cin(gnd),
	.combout(\Mux23~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~17 .lut_mask = 16'hBA98;
defparam \Mux23~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N20
cycloneive_lcell_comb \Mux23~18 (
// Equation(s):
// \Mux23~18_combout  = (\Mux23~17_combout  & (((\registerArray[15][8]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux23~17_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[14][8]~q ))))

	.dataa(\Mux23~17_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][8]~q ),
	.datad(\registerArray[14][8]~q ),
	.cin(gnd),
	.combout(\Mux23~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~18 .lut_mask = 16'hE6A2;
defparam \Mux23~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N22
cycloneive_lcell_comb \Mux22~7 (
// Equation(s):
// \Mux22~7_combout  = (\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o ) # ((\registerArray[27][9]~q )))) # (!\my_rf.rsel1[3]~input_o  & (!\my_rf.rsel1[2]~input_o  & (\registerArray[19][9]~q )))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[19][9]~q ),
	.datad(\registerArray[27][9]~q ),
	.cin(gnd),
	.combout(\Mux22~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~7 .lut_mask = 16'hBA98;
defparam \Mux22~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N2
cycloneive_lcell_comb \Mux22~10 (
// Equation(s):
// \Mux22~10_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[5][9]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[4][9]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[4][9]~q ),
	.datad(\registerArray[5][9]~q ),
	.cin(gnd),
	.combout(\Mux22~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~10 .lut_mask = 16'hDC98;
defparam \Mux22~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y37_N6
cycloneive_lcell_comb \Mux22~12 (
// Equation(s):
// \Mux22~12_combout  = (\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o )) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[10][9]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[8][9]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[8][9]~q ),
	.datad(\registerArray[10][9]~q ),
	.cin(gnd),
	.combout(\Mux22~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~12 .lut_mask = 16'hDC98;
defparam \Mux22~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y37_N30
cycloneive_lcell_comb \Mux22~13 (
// Equation(s):
// \Mux22~13_combout  = (\Mux22~12_combout  & (((\registerArray[11][9]~q )) # (!\my_rf.rsel1[0]~input_o ))) # (!\Mux22~12_combout  & (\my_rf.rsel1[0]~input_o  & ((\registerArray[9][9]~q ))))

	.dataa(\Mux22~12_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[11][9]~q ),
	.datad(\registerArray[9][9]~q ),
	.cin(gnd),
	.combout(\Mux22~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~13 .lut_mask = 16'hE6A2;
defparam \Mux22~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N20
cycloneive_lcell_comb \Mux22~17 (
// Equation(s):
// \Mux22~17_combout  = (\my_rf.rsel1[0]~input_o  & ((\registerArray[13][9]~q ) # ((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & (((\registerArray[12][9]~q  & !\my_rf.rsel1[1]~input_o ))))

	.dataa(\registerArray[13][9]~q ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][9]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux22~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~17 .lut_mask = 16'hCCB8;
defparam \Mux22~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N18
cycloneive_lcell_comb \Mux22~18 (
// Equation(s):
// \Mux22~18_combout  = (\Mux22~17_combout  & (((\registerArray[15][9]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux22~17_combout  & (\registerArray[14][9]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux22~17_combout ),
	.datab(\registerArray[14][9]~q ),
	.datac(\registerArray[15][9]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux22~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~18 .lut_mask = 16'hE4AA;
defparam \Mux22~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N26
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// \Mux21~0_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & (\registerArray[21][10]~q )) # (!\my_rf.rsel1[2]~input_o  & ((\registerArray[17][10]~q )))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[21][10]~q ),
	.datac(\registerArray[17][10]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hEE50;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N0
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// \Mux21~1_combout  = (\Mux21~0_combout  & (((\registerArray[29][10]~q ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux21~0_combout  & (\registerArray[25][10]~q  & ((\my_rf.rsel1[3]~input_o ))))

	.dataa(\Mux21~0_combout ),
	.datab(\registerArray[25][10]~q ),
	.datac(\registerArray[29][10]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'hE4AA;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N22
cycloneive_lcell_comb \Mux21~2 (
// Equation(s):
// \Mux21~2_combout  = (\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o ) # ((\registerArray[26][10]~q )))) # (!\my_rf.rsel1[3]~input_o  & (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][10]~q )))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][10]~q ),
	.datad(\registerArray[26][10]~q ),
	.cin(gnd),
	.combout(\Mux21~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~2 .lut_mask = 16'hBA98;
defparam \Mux21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N10
cycloneive_lcell_comb \Mux21~3 (
// Equation(s):
// \Mux21~3_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux21~2_combout  & (\registerArray[30][10]~q )) # (!\Mux21~2_combout  & ((\registerArray[22][10]~q ))))) # (!\my_rf.rsel1[2]~input_o  & (\Mux21~2_combout ))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux21~2_combout ),
	.datac(\registerArray[30][10]~q ),
	.datad(\registerArray[22][10]~q ),
	.cin(gnd),
	.combout(\Mux21~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~3 .lut_mask = 16'hE6C4;
defparam \Mux21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y37_N10
cycloneive_lcell_comb \Mux21~10 (
// Equation(s):
// \Mux21~10_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\registerArray[10][10]~q )) # (!\my_rf.rsel1[1]~input_o  & ((\registerArray[8][10]~q )))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\registerArray[10][10]~q ),
	.datac(\registerArray[8][10]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux21~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~10 .lut_mask = 16'hEE50;
defparam \Mux21~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N2
cycloneive_lcell_comb \Mux21~12 (
// Equation(s):
// \Mux21~12_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[5][10]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[4][10]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[4][10]~q ),
	.datad(\registerArray[5][10]~q ),
	.cin(gnd),
	.combout(\Mux21~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~12 .lut_mask = 16'hDC98;
defparam \Mux21~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N26
cycloneive_lcell_comb \Mux20~7 (
// Equation(s):
// \Mux20~7_combout  = (\my_rf.rsel1[3]~input_o  & ((\registerArray[27][11]~q ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((\registerArray[19][11]~q  & !\my_rf.rsel1[2]~input_o ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[27][11]~q ),
	.datac(\registerArray[19][11]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux20~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~7 .lut_mask = 16'hAAD8;
defparam \Mux20~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N30
cycloneive_lcell_comb \Mux20~10 (
// Equation(s):
// \Mux20~10_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[5][11]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[4][11]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[4][11]~q ),
	.datad(\registerArray[5][11]~q ),
	.cin(gnd),
	.combout(\Mux20~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~10 .lut_mask = 16'hDC98;
defparam \Mux20~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y37_N30
cycloneive_lcell_comb \Mux20~12 (
// Equation(s):
// \Mux20~12_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\registerArray[10][11]~q )) # (!\my_rf.rsel1[1]~input_o  & ((\registerArray[8][11]~q )))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\registerArray[10][11]~q ),
	.datac(\registerArray[8][11]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux20~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~12 .lut_mask = 16'hEE50;
defparam \Mux20~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y37_N14
cycloneive_lcell_comb \Mux20~13 (
// Equation(s):
// \Mux20~13_combout  = (\Mux20~12_combout  & (((\registerArray[11][11]~q ) # (!\my_rf.rsel1[0]~input_o )))) # (!\Mux20~12_combout  & (\registerArray[9][11]~q  & ((\my_rf.rsel1[0]~input_o ))))

	.dataa(\registerArray[9][11]~q ),
	.datab(\Mux20~12_combout ),
	.datac(\registerArray[11][11]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux20~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~13 .lut_mask = 16'hE2CC;
defparam \Mux20~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N18
cycloneive_lcell_comb \Mux20~14 (
// Equation(s):
// \Mux20~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][11]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][11]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[1][11]~q ),
	.datad(\registerArray[3][11]~q ),
	.cin(gnd),
	.combout(\Mux20~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~14 .lut_mask = 16'hC840;
defparam \Mux20~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N10
cycloneive_lcell_comb \Mux20~15 (
// Equation(s):
// \Mux20~15_combout  = (\Mux20~14_combout ) # ((\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & \registerArray[2][11]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux20~14_combout ),
	.datad(\registerArray[2][11]~q ),
	.cin(gnd),
	.combout(\Mux20~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~15 .lut_mask = 16'hF2F0;
defparam \Mux20~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N12
cycloneive_lcell_comb \Mux20~16 (
// Equation(s):
// \Mux20~16_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\Mux20~13_combout )) # (!\my_rf.rsel1[3]~input_o  & ((\Mux20~15_combout )))))

	.dataa(\Mux20~13_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\my_rf.rsel1[3]~input_o ),
	.datad(\Mux20~15_combout ),
	.cin(gnd),
	.combout(\Mux20~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~16 .lut_mask = 16'hE3E0;
defparam \Mux20~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N14
cycloneive_lcell_comb \Mux20~17 (
// Equation(s):
// \Mux20~17_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[13][11]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[12][11]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][11]~q ),
	.datad(\registerArray[13][11]~q ),
	.cin(gnd),
	.combout(\Mux20~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~17 .lut_mask = 16'hDC98;
defparam \Mux20~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N14
cycloneive_lcell_comb \Mux19~2 (
// Equation(s):
// \Mux19~2_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[26][12]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[18][12]~q )))))

	.dataa(\registerArray[26][12]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][12]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~2 .lut_mask = 16'hEE30;
defparam \Mux19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N0
cycloneive_lcell_comb \Mux19~3 (
// Equation(s):
// \Mux19~3_combout  = (\Mux19~2_combout  & (((\registerArray[30][12]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux19~2_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[22][12]~q ))))

	.dataa(\Mux19~2_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[30][12]~q ),
	.datad(\registerArray[22][12]~q ),
	.cin(gnd),
	.combout(\Mux19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~3 .lut_mask = 16'hE6A2;
defparam \Mux19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N6
cycloneive_lcell_comb \Mux19~4 (
// Equation(s):
// \Mux19~4_combout  = (\my_rf.rsel1[2]~input_o  & (\my_rf.rsel1[3]~input_o )) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & ((\registerArray[24][12]~q ))) # (!\my_rf.rsel1[3]~input_o  & (\registerArray[16][12]~q ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[16][12]~q ),
	.datad(\registerArray[24][12]~q ),
	.cin(gnd),
	.combout(\Mux19~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~4 .lut_mask = 16'hDC98;
defparam \Mux19~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N14
cycloneive_lcell_comb \Mux19~5 (
// Equation(s):
// \Mux19~5_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux19~4_combout  & (\registerArray[28][12]~q )) # (!\Mux19~4_combout  & ((\registerArray[20][12]~q ))))) # (!\my_rf.rsel1[2]~input_o  & (\Mux19~4_combout ))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux19~4_combout ),
	.datac(\registerArray[28][12]~q ),
	.datad(\registerArray[20][12]~q ),
	.cin(gnd),
	.combout(\Mux19~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~5 .lut_mask = 16'hE6C4;
defparam \Mux19~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N22
cycloneive_lcell_comb \Mux19~6 (
// Equation(s):
// \Mux19~6_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux19~3_combout ) # ((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & (((\Mux19~5_combout  & !\my_rf.rsel1[0]~input_o ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\Mux19~3_combout ),
	.datac(\Mux19~5_combout ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux19~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~6 .lut_mask = 16'hAAD8;
defparam \Mux19~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y37_N2
cycloneive_lcell_comb \Mux19~10 (
// Equation(s):
// \Mux19~10_combout  = (\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o )) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[10][12]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[8][12]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[8][12]~q ),
	.datad(\registerArray[10][12]~q ),
	.cin(gnd),
	.combout(\Mux19~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~10 .lut_mask = 16'hDC98;
defparam \Mux19~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N16
cycloneive_lcell_comb \Mux19~11 (
// Equation(s):
// \Mux19~11_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux19~10_combout  & ((\registerArray[11][12]~q ))) # (!\Mux19~10_combout  & (\registerArray[9][12]~q )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux19~10_combout ))))

	.dataa(\registerArray[9][12]~q ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[11][12]~q ),
	.datad(\Mux19~10_combout ),
	.cin(gnd),
	.combout(\Mux19~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~11 .lut_mask = 16'hF388;
defparam \Mux19~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N10
cycloneive_lcell_comb \Mux19~12 (
// Equation(s):
// \Mux19~12_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[5][12]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[4][12]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[4][12]~q ),
	.datad(\registerArray[5][12]~q ),
	.cin(gnd),
	.combout(\Mux19~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~12 .lut_mask = 16'hDC98;
defparam \Mux19~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N26
cycloneive_lcell_comb \Mux19~13 (
// Equation(s):
// \Mux19~13_combout  = (\Mux19~12_combout  & (((\registerArray[7][12]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux19~12_combout  & (\registerArray[6][12]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux19~12_combout ),
	.datab(\registerArray[6][12]~q ),
	.datac(\registerArray[7][12]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux19~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~13 .lut_mask = 16'hE4AA;
defparam \Mux19~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N10
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// \Mux18~0_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[25][13]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[17][13]~q )))))

	.dataa(\registerArray[25][13]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[17][13]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'hEE30;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N14
cycloneive_lcell_comb \Mux18~10 (
// Equation(s):
// \Mux18~10_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[5][13]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[4][13]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[4][13]~q ),
	.datad(\registerArray[5][13]~q ),
	.cin(gnd),
	.combout(\Mux18~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~10 .lut_mask = 16'hDC98;
defparam \Mux18~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y37_N14
cycloneive_lcell_comb \Mux18~12 (
// Equation(s):
// \Mux18~12_combout  = (\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o )) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[10][13]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[8][13]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[8][13]~q ),
	.datad(\registerArray[10][13]~q ),
	.cin(gnd),
	.combout(\Mux18~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~12 .lut_mask = 16'hDC98;
defparam \Mux18~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y37_N4
cycloneive_lcell_comb \Mux18~13 (
// Equation(s):
// \Mux18~13_combout  = (\Mux18~12_combout  & (((\registerArray[11][13]~q )) # (!\my_rf.rsel1[0]~input_o ))) # (!\Mux18~12_combout  & (\my_rf.rsel1[0]~input_o  & ((\registerArray[9][13]~q ))))

	.dataa(\Mux18~12_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[11][13]~q ),
	.datad(\registerArray[9][13]~q ),
	.cin(gnd),
	.combout(\Mux18~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~13 .lut_mask = 16'hE6A2;
defparam \Mux18~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N26
cycloneive_lcell_comb \Mux18~14 (
// Equation(s):
// \Mux18~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][13]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][13]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[1][13]~q ),
	.datad(\registerArray[3][13]~q ),
	.cin(gnd),
	.combout(\Mux18~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~14 .lut_mask = 16'hC840;
defparam \Mux18~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y36_N20
cycloneive_lcell_comb \Mux18~15 (
// Equation(s):
// \Mux18~15_combout  = (\Mux18~14_combout ) # ((\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & \registerArray[2][13]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[2][13]~q ),
	.datad(\Mux18~14_combout ),
	.cin(gnd),
	.combout(\Mux18~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~15 .lut_mask = 16'hFF20;
defparam \Mux18~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N18
cycloneive_lcell_comb \Mux18~16 (
// Equation(s):
// \Mux18~16_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\Mux18~13_combout )) # (!\my_rf.rsel1[3]~input_o  & ((\Mux18~15_combout )))))

	.dataa(\Mux18~13_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\my_rf.rsel1[3]~input_o ),
	.datad(\Mux18~15_combout ),
	.cin(gnd),
	.combout(\Mux18~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~16 .lut_mask = 16'hE3E0;
defparam \Mux18~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N30
cycloneive_lcell_comb \Mux17~2 (
// Equation(s):
// \Mux17~2_combout  = (\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o ) # ((\registerArray[26][14]~q )))) # (!\my_rf.rsel1[3]~input_o  & (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][14]~q )))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][14]~q ),
	.datad(\registerArray[26][14]~q ),
	.cin(gnd),
	.combout(\Mux17~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~2 .lut_mask = 16'hBA98;
defparam \Mux17~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y38_N20
cycloneive_lcell_comb \Mux17~3 (
// Equation(s):
// \Mux17~3_combout  = (\Mux17~2_combout  & (((\registerArray[30][14]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux17~2_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[22][14]~q ))))

	.dataa(\Mux17~2_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[30][14]~q ),
	.datad(\registerArray[22][14]~q ),
	.cin(gnd),
	.combout(\Mux17~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~3 .lut_mask = 16'hE6A2;
defparam \Mux17~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N18
cycloneive_lcell_comb \Mux17~4 (
// Equation(s):
// \Mux17~4_combout  = (\my_rf.rsel1[2]~input_o  & (\my_rf.rsel1[3]~input_o )) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & ((\registerArray[24][14]~q ))) # (!\my_rf.rsel1[3]~input_o  & (\registerArray[16][14]~q ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[16][14]~q ),
	.datad(\registerArray[24][14]~q ),
	.cin(gnd),
	.combout(\Mux17~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~4 .lut_mask = 16'hDC98;
defparam \Mux17~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N22
cycloneive_lcell_comb \Mux17~5 (
// Equation(s):
// \Mux17~5_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux17~4_combout  & (\registerArray[28][14]~q )) # (!\Mux17~4_combout  & ((\registerArray[20][14]~q ))))) # (!\my_rf.rsel1[2]~input_o  & (\Mux17~4_combout ))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux17~4_combout ),
	.datac(\registerArray[28][14]~q ),
	.datad(\registerArray[20][14]~q ),
	.cin(gnd),
	.combout(\Mux17~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~5 .lut_mask = 16'hE6C4;
defparam \Mux17~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y38_N26
cycloneive_lcell_comb \Mux17~6 (
// Equation(s):
// \Mux17~6_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\Mux17~3_combout )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & (\Mux17~5_combout )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux17~5_combout ),
	.datad(\Mux17~3_combout ),
	.cin(gnd),
	.combout(\Mux17~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~6 .lut_mask = 16'hBA98;
defparam \Mux17~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N30
cycloneive_lcell_comb \Mux17~7 (
// Equation(s):
// \Mux17~7_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[23][14]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[19][14]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[19][14]~q ),
	.datad(\registerArray[23][14]~q ),
	.cin(gnd),
	.combout(\Mux17~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~7 .lut_mask = 16'hDC98;
defparam \Mux17~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N18
cycloneive_lcell_comb \Mux17~12 (
// Equation(s):
// \Mux17~12_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[5][14]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[4][14]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[4][14]~q ),
	.datad(\registerArray[5][14]~q ),
	.cin(gnd),
	.combout(\Mux17~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~12 .lut_mask = 16'hDC98;
defparam \Mux17~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y36_N30
cycloneive_lcell_comb \Mux17~17 (
// Equation(s):
// \Mux17~17_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[13][14]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[12][14]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][14]~q ),
	.datad(\registerArray[13][14]~q ),
	.cin(gnd),
	.combout(\Mux17~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~17 .lut_mask = 16'hDC98;
defparam \Mux17~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N22
cycloneive_lcell_comb \Mux16~4 (
// Equation(s):
// \Mux16~4_combout  = (\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o ) # ((\registerArray[20][15]~q )))) # (!\my_rf.rsel1[2]~input_o  & (!\my_rf.rsel1[3]~input_o  & (\registerArray[16][15]~q )))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[16][15]~q ),
	.datad(\registerArray[20][15]~q ),
	.cin(gnd),
	.combout(\Mux16~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~4 .lut_mask = 16'hBA98;
defparam \Mux16~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N0
cycloneive_lcell_comb \Mux16~5 (
// Equation(s):
// \Mux16~5_combout  = (\Mux16~4_combout  & (((\registerArray[28][15]~q ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux16~4_combout  & (\registerArray[24][15]~q  & ((\my_rf.rsel1[3]~input_o ))))

	.dataa(\Mux16~4_combout ),
	.datab(\registerArray[24][15]~q ),
	.datac(\registerArray[28][15]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux16~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~5 .lut_mask = 16'hE4AA;
defparam \Mux16~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N18
cycloneive_lcell_comb \Mux16~7 (
// Equation(s):
// \Mux16~7_combout  = (\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o ) # ((\registerArray[27][15]~q )))) # (!\my_rf.rsel1[3]~input_o  & (!\my_rf.rsel1[2]~input_o  & (\registerArray[19][15]~q )))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[19][15]~q ),
	.datad(\registerArray[27][15]~q ),
	.cin(gnd),
	.combout(\Mux16~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~7 .lut_mask = 16'hBA98;
defparam \Mux16~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N26
cycloneive_lcell_comb \Mux16~8 (
// Equation(s):
// \Mux16~8_combout  = (\Mux16~7_combout  & (((\registerArray[31][15]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux16~7_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[23][15]~q ))))

	.dataa(\Mux16~7_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[31][15]~q ),
	.datad(\registerArray[23][15]~q ),
	.cin(gnd),
	.combout(\Mux16~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~8 .lut_mask = 16'hE6A2;
defparam \Mux16~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N18
cycloneive_lcell_comb \Mux16~12 (
// Equation(s):
// \Mux16~12_combout  = (\my_rf.rsel1[1]~input_o  & ((\registerArray[10][15]~q ) # ((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & (((\registerArray[8][15]~q  & !\my_rf.rsel1[0]~input_o ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[10][15]~q ),
	.datac(\registerArray[8][15]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux16~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~12 .lut_mask = 16'hAAD8;
defparam \Mux16~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N18
cycloneive_lcell_comb \Mux16~13 (
// Equation(s):
// \Mux16~13_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux16~12_combout  & (\registerArray[11][15]~q )) # (!\Mux16~12_combout  & ((\registerArray[9][15]~q ))))) # (!\my_rf.rsel1[0]~input_o  & (\Mux16~12_combout ))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux16~12_combout ),
	.datac(\registerArray[11][15]~q ),
	.datad(\registerArray[9][15]~q ),
	.cin(gnd),
	.combout(\Mux16~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~13 .lut_mask = 16'hE6C4;
defparam \Mux16~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N2
cycloneive_lcell_comb \Mux16~14 (
// Equation(s):
// \Mux16~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][15]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][15]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[1][15]~q ),
	.datad(\registerArray[3][15]~q ),
	.cin(gnd),
	.combout(\Mux16~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~14 .lut_mask = 16'hC840;
defparam \Mux16~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y36_N18
cycloneive_lcell_comb \Mux16~15 (
// Equation(s):
// \Mux16~15_combout  = (\Mux16~14_combout ) # ((\registerArray[2][15]~q  & (!\my_rf.rsel1[0]~input_o  & \my_rf.rsel1[1]~input_o )))

	.dataa(\registerArray[2][15]~q ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\Mux16~14_combout ),
	.cin(gnd),
	.combout(\Mux16~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~15 .lut_mask = 16'hFF20;
defparam \Mux16~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y38_N22
cycloneive_lcell_comb \Mux16~16 (
// Equation(s):
// \Mux16~16_combout  = (\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o ) # ((\Mux16~13_combout )))) # (!\my_rf.rsel1[3]~input_o  & (!\my_rf.rsel1[2]~input_o  & ((\Mux16~15_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux16~13_combout ),
	.datad(\Mux16~15_combout ),
	.cin(gnd),
	.combout(\Mux16~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~16 .lut_mask = 16'hB9A8;
defparam \Mux16~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y36_N10
cycloneive_lcell_comb \Mux16~17 (
// Equation(s):
// \Mux16~17_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[13][15]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[12][15]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][15]~q ),
	.datad(\registerArray[13][15]~q ),
	.cin(gnd),
	.combout(\Mux16~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~17 .lut_mask = 16'hDC98;
defparam \Mux16~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N2
cycloneive_lcell_comb \Mux15~4 (
// Equation(s):
// \Mux15~4_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[24][16]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[16][16]~q )))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[24][16]~q ),
	.datac(\registerArray[16][16]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux15~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~4 .lut_mask = 16'hEE50;
defparam \Mux15~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N24
cycloneive_lcell_comb \Mux15~7 (
// Equation(s):
// \Mux15~7_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & (\registerArray[23][16]~q )) # (!\my_rf.rsel1[2]~input_o  & ((\registerArray[19][16]~q )))))

	.dataa(\registerArray[23][16]~q ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[19][16]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux15~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~7 .lut_mask = 16'hEE30;
defparam \Mux15~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N14
cycloneive_lcell_comb \Mux15~8 (
// Equation(s):
// \Mux15~8_combout  = (\Mux15~7_combout  & (((\registerArray[31][16]~q ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux15~7_combout  & (\registerArray[27][16]~q  & ((\my_rf.rsel1[3]~input_o ))))

	.dataa(\registerArray[27][16]~q ),
	.datab(\Mux15~7_combout ),
	.datac(\registerArray[31][16]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux15~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~8 .lut_mask = 16'hE2CC;
defparam \Mux15~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N18
cycloneive_lcell_comb \Mux15~12 (
// Equation(s):
// \Mux15~12_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[5][16]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[4][16]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[4][16]~q ),
	.datad(\registerArray[5][16]~q ),
	.cin(gnd),
	.combout(\Mux15~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~12 .lut_mask = 16'hDC98;
defparam \Mux15~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N14
cycloneive_lcell_comb \Mux15~13 (
// Equation(s):
// \Mux15~13_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux15~12_combout  & (\registerArray[7][16]~q )) # (!\Mux15~12_combout  & ((\registerArray[6][16]~q ))))) # (!\my_rf.rsel1[1]~input_o  & (\Mux15~12_combout ))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\Mux15~12_combout ),
	.datac(\registerArray[7][16]~q ),
	.datad(\registerArray[6][16]~q ),
	.cin(gnd),
	.combout(\Mux15~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~13 .lut_mask = 16'hE6C4;
defparam \Mux15~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y36_N6
cycloneive_lcell_comb \Mux15~17 (
// Equation(s):
// \Mux15~17_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[13][16]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[12][16]~q )))))

	.dataa(\registerArray[13][16]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[12][16]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux15~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~17 .lut_mask = 16'hEE30;
defparam \Mux15~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N2
cycloneive_lcell_comb \Mux15~18 (
// Equation(s):
// \Mux15~18_combout  = (\Mux15~17_combout  & (((\registerArray[15][16]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux15~17_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[14][16]~q ))))

	.dataa(\Mux15~17_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][16]~q ),
	.datad(\registerArray[14][16]~q ),
	.cin(gnd),
	.combout(\Mux15~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~18 .lut_mask = 16'hE6A2;
defparam \Mux15~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N22
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// \Mux14~0_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[25][17]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[17][17]~q )))))

	.dataa(\registerArray[25][17]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[17][17]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hEE30;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N24
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// \Mux14~1_combout  = (\Mux14~0_combout  & (((\registerArray[29][17]~q ) # (!\my_rf.rsel1[2]~input_o )))) # (!\Mux14~0_combout  & (\registerArray[21][17]~q  & ((\my_rf.rsel1[2]~input_o ))))

	.dataa(\Mux14~0_combout ),
	.datab(\registerArray[21][17]~q ),
	.datac(\registerArray[29][17]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hE4AA;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N14
cycloneive_lcell_comb \Mux14~7 (
// Equation(s):
// \Mux14~7_combout  = (\my_rf.rsel1[3]~input_o  & ((\registerArray[27][17]~q ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((\registerArray[19][17]~q  & !\my_rf.rsel1[2]~input_o ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[27][17]~q ),
	.datac(\registerArray[19][17]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux14~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~7 .lut_mask = 16'hAAD8;
defparam \Mux14~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N22
cycloneive_lcell_comb \Mux14~10 (
// Equation(s):
// \Mux14~10_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[5][17]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[4][17]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[4][17]~q ),
	.datad(\registerArray[5][17]~q ),
	.cin(gnd),
	.combout(\Mux14~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~10 .lut_mask = 16'hDC98;
defparam \Mux14~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N18
cycloneive_lcell_comb \Mux14~11 (
// Equation(s):
// \Mux14~11_combout  = (\Mux14~10_combout  & (((\registerArray[7][17]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux14~10_combout  & (\registerArray[6][17]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux14~10_combout ),
	.datab(\registerArray[6][17]~q ),
	.datac(\registerArray[7][17]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux14~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~11 .lut_mask = 16'hE4AA;
defparam \Mux14~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N2
cycloneive_lcell_comb \Mux14~12 (
// Equation(s):
// \Mux14~12_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\registerArray[10][17]~q )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & (\registerArray[8][17]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[8][17]~q ),
	.datad(\registerArray[10][17]~q ),
	.cin(gnd),
	.combout(\Mux14~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~12 .lut_mask = 16'hBA98;
defparam \Mux14~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N2
cycloneive_lcell_comb \Mux14~13 (
// Equation(s):
// \Mux14~13_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux14~12_combout  & ((\registerArray[11][17]~q ))) # (!\Mux14~12_combout  & (\registerArray[9][17]~q )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux14~12_combout ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\registerArray[9][17]~q ),
	.datac(\registerArray[11][17]~q ),
	.datad(\Mux14~12_combout ),
	.cin(gnd),
	.combout(\Mux14~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~13 .lut_mask = 16'hF588;
defparam \Mux14~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N2
cycloneive_lcell_comb \Mux14~17 (
// Equation(s):
// \Mux14~17_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[13][17]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[12][17]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][17]~q ),
	.datad(\registerArray[13][17]~q ),
	.cin(gnd),
	.combout(\Mux14~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~17 .lut_mask = 16'hDC98;
defparam \Mux14~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N24
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// \Mux13~0_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[21][18]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[17][18]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[17][18]~q ),
	.datad(\registerArray[21][18]~q ),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hDC98;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N28
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// \Mux13~1_combout  = (\Mux13~0_combout  & (((\registerArray[29][18]~q ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux13~0_combout  & (\registerArray[25][18]~q  & ((\my_rf.rsel1[3]~input_o ))))

	.dataa(\registerArray[25][18]~q ),
	.datab(\Mux13~0_combout ),
	.datac(\registerArray[29][18]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'hE2CC;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N0
cycloneive_lcell_comb \Mux13~4 (
// Equation(s):
// \Mux13~4_combout  = (\my_rf.rsel1[3]~input_o  & ((\registerArray[24][18]~q ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((\registerArray[16][18]~q  & !\my_rf.rsel1[2]~input_o ))))

	.dataa(\registerArray[24][18]~q ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[16][18]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux13~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~4 .lut_mask = 16'hCCB8;
defparam \Mux13~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N30
cycloneive_lcell_comb \Mux13~10 (
// Equation(s):
// \Mux13~10_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\registerArray[10][18]~q )) # (!\my_rf.rsel1[1]~input_o  & ((\registerArray[8][18]~q )))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\registerArray[10][18]~q ),
	.datac(\registerArray[8][18]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux13~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~10 .lut_mask = 16'hEE50;
defparam \Mux13~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N14
cycloneive_lcell_comb \Mux13~12 (
// Equation(s):
// \Mux13~12_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o ) # ((\registerArray[5][18]~q )))) # (!\my_rf.rsel1[0]~input_o  & (!\my_rf.rsel1[1]~input_o  & (\registerArray[4][18]~q )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[4][18]~q ),
	.datad(\registerArray[5][18]~q ),
	.cin(gnd),
	.combout(\Mux13~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~12 .lut_mask = 16'hBA98;
defparam \Mux13~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N30
cycloneive_lcell_comb \Mux13~13 (
// Equation(s):
// \Mux13~13_combout  = (\Mux13~12_combout  & (((\registerArray[7][18]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux13~12_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[6][18]~q ))))

	.dataa(\Mux13~12_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[7][18]~q ),
	.datad(\registerArray[6][18]~q ),
	.cin(gnd),
	.combout(\Mux13~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~13 .lut_mask = 16'hE6A2;
defparam \Mux13~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N18
cycloneive_lcell_comb \Mux13~14 (
// Equation(s):
// \Mux13~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][18]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][18]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[1][18]~q ),
	.datad(\registerArray[3][18]~q ),
	.cin(gnd),
	.combout(\Mux13~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~14 .lut_mask = 16'hC840;
defparam \Mux13~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N8
cycloneive_lcell_comb \Mux13~15 (
// Equation(s):
// \Mux13~15_combout  = (\Mux13~14_combout ) # ((!\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o  & \registerArray[2][18]~q )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux13~14_combout ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\registerArray[2][18]~q ),
	.cin(gnd),
	.combout(\Mux13~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~15 .lut_mask = 16'hDCCC;
defparam \Mux13~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N10
cycloneive_lcell_comb \Mux13~16 (
// Equation(s):
// \Mux13~16_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux13~13_combout ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux13~15_combout  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux13~13_combout ),
	.datac(\Mux13~15_combout ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux13~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~16 .lut_mask = 16'hAAD8;
defparam \Mux13~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N18
cycloneive_lcell_comb \Mux13~17 (
// Equation(s):
// \Mux13~17_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o ) # ((\registerArray[13][18]~q )))) # (!\my_rf.rsel1[0]~input_o  & (!\my_rf.rsel1[1]~input_o  & (\registerArray[12][18]~q )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[12][18]~q ),
	.datad(\registerArray[13][18]~q ),
	.cin(gnd),
	.combout(\Mux13~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~17 .lut_mask = 16'hBA98;
defparam \Mux13~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N18
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (\my_rf.rsel1[2]~input_o  & (\my_rf.rsel1[3]~input_o )) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & ((\registerArray[25][19]~q ))) # (!\my_rf.rsel1[3]~input_o  & (\registerArray[17][19]~q ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[17][19]~q ),
	.datad(\registerArray[25][19]~q ),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hDC98;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N30
cycloneive_lcell_comb \Mux12~2 (
// Equation(s):
// \Mux12~2_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[22][19]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][19]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][19]~q ),
	.datad(\registerArray[22][19]~q ),
	.cin(gnd),
	.combout(\Mux12~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~2 .lut_mask = 16'hDC98;
defparam \Mux12~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y38_N8
cycloneive_lcell_comb \Mux12~3 (
// Equation(s):
// \Mux12~3_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux12~2_combout  & (\registerArray[30][19]~q )) # (!\Mux12~2_combout  & ((\registerArray[26][19]~q ))))) # (!\my_rf.rsel1[3]~input_o  & (\Mux12~2_combout ))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux12~2_combout ),
	.datac(\registerArray[30][19]~q ),
	.datad(\registerArray[26][19]~q ),
	.cin(gnd),
	.combout(\Mux12~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~3 .lut_mask = 16'hE6C4;
defparam \Mux12~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N10
cycloneive_lcell_comb \Mux12~7 (
// Equation(s):
// \Mux12~7_combout  = (\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o ) # ((\registerArray[27][19]~q )))) # (!\my_rf.rsel1[3]~input_o  & (!\my_rf.rsel1[2]~input_o  & (\registerArray[19][19]~q )))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[19][19]~q ),
	.datad(\registerArray[27][19]~q ),
	.cin(gnd),
	.combout(\Mux12~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~7 .lut_mask = 16'hBA98;
defparam \Mux12~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N16
cycloneive_lcell_comb \Mux12~8 (
// Equation(s):
// \Mux12~8_combout  = (\Mux12~7_combout  & (((\registerArray[31][19]~q ) # (!\my_rf.rsel1[2]~input_o )))) # (!\Mux12~7_combout  & (\registerArray[23][19]~q  & ((\my_rf.rsel1[2]~input_o ))))

	.dataa(\registerArray[23][19]~q ),
	.datab(\Mux12~7_combout ),
	.datac(\registerArray[31][19]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux12~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~8 .lut_mask = 16'hE2CC;
defparam \Mux12~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N22
cycloneive_lcell_comb \Mux12~12 (
// Equation(s):
// \Mux12~12_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\registerArray[10][19]~q )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & (\registerArray[8][19]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[8][19]~q ),
	.datad(\registerArray[10][19]~q ),
	.cin(gnd),
	.combout(\Mux12~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~12 .lut_mask = 16'hBA98;
defparam \Mux12~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N14
cycloneive_lcell_comb \Mux12~13 (
// Equation(s):
// \Mux12~13_combout  = (\Mux12~12_combout  & (((\registerArray[11][19]~q ) # (!\my_rf.rsel1[0]~input_o )))) # (!\Mux12~12_combout  & (\registerArray[9][19]~q  & ((\my_rf.rsel1[0]~input_o ))))

	.dataa(\registerArray[9][19]~q ),
	.datab(\Mux12~12_combout ),
	.datac(\registerArray[11][19]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux12~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~13 .lut_mask = 16'hE2CC;
defparam \Mux12~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N30
cycloneive_lcell_comb \Mux12~14 (
// Equation(s):
// \Mux12~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][19]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][19]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[1][19]~q ),
	.datad(\registerArray[3][19]~q ),
	.cin(gnd),
	.combout(\Mux12~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~14 .lut_mask = 16'hA820;
defparam \Mux12~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N16
cycloneive_lcell_comb \Mux12~17 (
// Equation(s):
// \Mux12~17_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[13][19]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[12][19]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][19]~q ),
	.datad(\registerArray[13][19]~q ),
	.cin(gnd),
	.combout(\Mux12~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~17 .lut_mask = 16'hDC98;
defparam \Mux12~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N24
cycloneive_lcell_comb \Mux12~18 (
// Equation(s):
// \Mux12~18_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux12~17_combout  & ((\registerArray[15][19]~q ))) # (!\Mux12~17_combout  & (\registerArray[14][19]~q )))) # (!\my_rf.rsel1[1]~input_o  & (((\Mux12~17_combout ))))

	.dataa(\registerArray[14][19]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][19]~q ),
	.datad(\Mux12~17_combout ),
	.cin(gnd),
	.combout(\Mux12~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~18 .lut_mask = 16'hF388;
defparam \Mux12~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N26
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// \Mux11~0_combout  = (\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o ) # ((\registerArray[21][20]~q )))) # (!\my_rf.rsel1[2]~input_o  & (!\my_rf.rsel1[3]~input_o  & (\registerArray[17][20]~q )))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[17][20]~q ),
	.datad(\registerArray[21][20]~q ),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hBA98;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N24
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// \Mux11~1_combout  = (\Mux11~0_combout  & (((\registerArray[29][20]~q ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux11~0_combout  & (\registerArray[25][20]~q  & ((\my_rf.rsel1[3]~input_o ))))

	.dataa(\Mux11~0_combout ),
	.datab(\registerArray[25][20]~q ),
	.datac(\registerArray[29][20]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'hE4AA;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N8
cycloneive_lcell_comb \Mux11~2 (
// Equation(s):
// \Mux11~2_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[26][20]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[18][20]~q )))))

	.dataa(\registerArray[26][20]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][20]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~2 .lut_mask = 16'hEE30;
defparam \Mux11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N26
cycloneive_lcell_comb \Mux11~14 (
// Equation(s):
// \Mux11~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][20]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][20]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[1][20]~q ),
	.datad(\registerArray[3][20]~q ),
	.cin(gnd),
	.combout(\Mux11~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~14 .lut_mask = 16'hC840;
defparam \Mux11~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N22
cycloneive_lcell_comb \Mux11~17 (
// Equation(s):
// \Mux11~17_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[13][20]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[12][20]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][20]~q ),
	.datad(\registerArray[13][20]~q ),
	.cin(gnd),
	.combout(\Mux11~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~17 .lut_mask = 16'hDC98;
defparam \Mux11~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N28
cycloneive_lcell_comb \Mux10~7 (
// Equation(s):
// \Mux10~7_combout  = (\my_rf.rsel1[2]~input_o  & (\my_rf.rsel1[3]~input_o )) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & ((\registerArray[27][21]~q ))) # (!\my_rf.rsel1[3]~input_o  & (\registerArray[19][21]~q ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[19][21]~q ),
	.datad(\registerArray[27][21]~q ),
	.cin(gnd),
	.combout(\Mux10~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~7 .lut_mask = 16'hDC98;
defparam \Mux10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N18
cycloneive_lcell_comb \Mux10~8 (
// Equation(s):
// \Mux10~8_combout  = (\Mux10~7_combout  & (((\registerArray[31][21]~q ) # (!\my_rf.rsel1[2]~input_o )))) # (!\Mux10~7_combout  & (\registerArray[23][21]~q  & ((\my_rf.rsel1[2]~input_o ))))

	.dataa(\registerArray[23][21]~q ),
	.datab(\Mux10~7_combout ),
	.datac(\registerArray[31][21]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux10~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~8 .lut_mask = 16'hE2CC;
defparam \Mux10~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N8
cycloneive_lcell_comb \Mux10~10 (
// Equation(s):
// \Mux10~10_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[5][21]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[4][21]~q )))))

	.dataa(\registerArray[5][21]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[4][21]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux10~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~10 .lut_mask = 16'hEE30;
defparam \Mux10~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N26
cycloneive_lcell_comb \Mux10~12 (
// Equation(s):
// \Mux10~12_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\registerArray[10][21]~q )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & (\registerArray[8][21]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[8][21]~q ),
	.datad(\registerArray[10][21]~q ),
	.cin(gnd),
	.combout(\Mux10~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~12 .lut_mask = 16'hBA98;
defparam \Mux10~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N10
cycloneive_lcell_comb \Mux10~13 (
// Equation(s):
// \Mux10~13_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux10~12_combout  & (\registerArray[11][21]~q )) # (!\Mux10~12_combout  & ((\registerArray[9][21]~q ))))) # (!\my_rf.rsel1[0]~input_o  & (\Mux10~12_combout ))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux10~12_combout ),
	.datac(\registerArray[11][21]~q ),
	.datad(\registerArray[9][21]~q ),
	.cin(gnd),
	.combout(\Mux10~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~13 .lut_mask = 16'hE6C4;
defparam \Mux10~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N2
cycloneive_lcell_comb \Mux10~17 (
// Equation(s):
// \Mux10~17_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[13][21]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[12][21]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][21]~q ),
	.datad(\registerArray[13][21]~q ),
	.cin(gnd),
	.combout(\Mux10~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~17 .lut_mask = 16'hDC98;
defparam \Mux10~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N24
cycloneive_lcell_comb \Mux9~2 (
// Equation(s):
// \Mux9~2_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[26][22]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[18][22]~q )))))

	.dataa(\registerArray[26][22]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][22]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux9~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~2 .lut_mask = 16'hEE30;
defparam \Mux9~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N20
cycloneive_lcell_comb \Mux9~3 (
// Equation(s):
// \Mux9~3_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux9~2_combout  & ((\registerArray[30][22]~q ))) # (!\Mux9~2_combout  & (\registerArray[22][22]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux9~2_combout ))))

	.dataa(\registerArray[22][22]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[30][22]~q ),
	.datad(\Mux9~2_combout ),
	.cin(gnd),
	.combout(\Mux9~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~3 .lut_mask = 16'hF388;
defparam \Mux9~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N22
cycloneive_lcell_comb \Mux9~4 (
// Equation(s):
// \Mux9~4_combout  = (\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o ) # ((\registerArray[24][22]~q )))) # (!\my_rf.rsel1[3]~input_o  & (!\my_rf.rsel1[2]~input_o  & (\registerArray[16][22]~q )))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[16][22]~q ),
	.datad(\registerArray[24][22]~q ),
	.cin(gnd),
	.combout(\Mux9~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~4 .lut_mask = 16'hBA98;
defparam \Mux9~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N26
cycloneive_lcell_comb \Mux9~5 (
// Equation(s):
// \Mux9~5_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux9~4_combout  & ((\registerArray[28][22]~q ))) # (!\Mux9~4_combout  & (\registerArray[20][22]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux9~4_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[20][22]~q ),
	.datac(\registerArray[28][22]~q ),
	.datad(\Mux9~4_combout ),
	.cin(gnd),
	.combout(\Mux9~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~5 .lut_mask = 16'hF588;
defparam \Mux9~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N10
cycloneive_lcell_comb \Mux9~6 (
// Equation(s):
// \Mux9~6_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\Mux9~3_combout ))) # (!\my_rf.rsel1[1]~input_o  & (\Mux9~5_combout ))))

	.dataa(\Mux9~5_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\Mux9~3_combout ),
	.cin(gnd),
	.combout(\Mux9~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~6 .lut_mask = 16'hF2C2;
defparam \Mux9~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N26
cycloneive_lcell_comb \Mux9~7 (
// Equation(s):
// \Mux9~7_combout  = (\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o ) # ((\registerArray[23][22]~q )))) # (!\my_rf.rsel1[2]~input_o  & (!\my_rf.rsel1[3]~input_o  & (\registerArray[19][22]~q )))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[19][22]~q ),
	.datad(\registerArray[23][22]~q ),
	.cin(gnd),
	.combout(\Mux9~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~7 .lut_mask = 16'hBA98;
defparam \Mux9~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N4
cycloneive_lcell_comb \Mux9~12 (
// Equation(s):
// \Mux9~12_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[5][22]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[4][22]~q )))))

	.dataa(\registerArray[5][22]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[4][22]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux9~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~12 .lut_mask = 16'hEE30;
defparam \Mux9~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N10
cycloneive_lcell_comb \Mux9~14 (
// Equation(s):
// \Mux9~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][22]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][22]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[1][22]~q ),
	.datad(\registerArray[3][22]~q ),
	.cin(gnd),
	.combout(\Mux9~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~14 .lut_mask = 16'hC840;
defparam \Mux9~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N22
cycloneive_lcell_comb \Mux9~15 (
// Equation(s):
// \Mux9~15_combout  = (\Mux9~14_combout ) # ((\my_rf.rsel1[1]~input_o  & (\registerArray[2][22]~q  & !\my_rf.rsel1[0]~input_o )))

	.dataa(\Mux9~14_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[2][22]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux9~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~15 .lut_mask = 16'hAAEA;
defparam \Mux9~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N18
cycloneive_lcell_comb \Mux9~17 (
// Equation(s):
// \Mux9~17_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[13][22]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[12][22]~q )))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[13][22]~q ),
	.datac(\registerArray[12][22]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux9~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~17 .lut_mask = 16'hEE50;
defparam \Mux9~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N10
cycloneive_lcell_comb \Mux9~18 (
// Equation(s):
// \Mux9~18_combout  = (\Mux9~17_combout  & (((\registerArray[15][22]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux9~17_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[14][22]~q ))))

	.dataa(\Mux9~17_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][22]~q ),
	.datad(\registerArray[14][22]~q ),
	.cin(gnd),
	.combout(\Mux9~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~18 .lut_mask = 16'hE6A2;
defparam \Mux9~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N14
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// \Mux8~0_combout  = (\my_rf.rsel1[3]~input_o  & ((\registerArray[25][23]~q ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((\registerArray[17][23]~q  & !\my_rf.rsel1[2]~input_o ))))

	.dataa(\registerArray[25][23]~q ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[17][23]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hCCB8;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N20
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// \Mux8~1_combout  = (\Mux8~0_combout  & (((\registerArray[29][23]~q ) # (!\my_rf.rsel1[2]~input_o )))) # (!\Mux8~0_combout  & (\registerArray[21][23]~q  & ((\my_rf.rsel1[2]~input_o ))))

	.dataa(\Mux8~0_combout ),
	.datab(\registerArray[21][23]~q ),
	.datac(\registerArray[29][23]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'hE4AA;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N10
cycloneive_lcell_comb \Mux8~2 (
// Equation(s):
// \Mux8~2_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[22][23]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][23]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][23]~q ),
	.datad(\registerArray[22][23]~q ),
	.cin(gnd),
	.combout(\Mux8~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~2 .lut_mask = 16'hDC98;
defparam \Mux8~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N16
cycloneive_lcell_comb \Mux8~4 (
// Equation(s):
// \Mux8~4_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[20][23]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[16][23]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[16][23]~q ),
	.datad(\registerArray[20][23]~q ),
	.cin(gnd),
	.combout(\Mux8~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~4 .lut_mask = 16'hDC98;
defparam \Mux8~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N6
cycloneive_lcell_comb \Mux8~5 (
// Equation(s):
// \Mux8~5_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux8~4_combout  & (\registerArray[28][23]~q )) # (!\Mux8~4_combout  & ((\registerArray[24][23]~q ))))) # (!\my_rf.rsel1[3]~input_o  & (\Mux8~4_combout ))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux8~4_combout ),
	.datac(\registerArray[28][23]~q ),
	.datad(\registerArray[24][23]~q ),
	.cin(gnd),
	.combout(\Mux8~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~5 .lut_mask = 16'hE6C4;
defparam \Mux8~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N24
cycloneive_lcell_comb \Mux8~10 (
// Equation(s):
// \Mux8~10_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[5][23]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[4][23]~q )))))

	.dataa(\registerArray[5][23]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[4][23]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux8~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~10 .lut_mask = 16'hEE30;
defparam \Mux8~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y31_N14
cycloneive_lcell_comb \Mux8~11 (
// Equation(s):
// \Mux8~11_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux8~10_combout  & ((\registerArray[7][23]~q ))) # (!\Mux8~10_combout  & (\registerArray[6][23]~q )))) # (!\my_rf.rsel1[1]~input_o  & (((\Mux8~10_combout ))))

	.dataa(\registerArray[6][23]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[7][23]~q ),
	.datad(\Mux8~10_combout ),
	.cin(gnd),
	.combout(\Mux8~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~11 .lut_mask = 16'hF388;
defparam \Mux8~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N30
cycloneive_lcell_comb \Mux8~14 (
// Equation(s):
// \Mux8~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][23]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][23]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[1][23]~q ),
	.datad(\registerArray[3][23]~q ),
	.cin(gnd),
	.combout(\Mux8~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~14 .lut_mask = 16'hC840;
defparam \Mux8~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N30
cycloneive_lcell_comb \Mux8~15 (
// Equation(s):
// \Mux8~15_combout  = (\Mux8~14_combout ) # ((!\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o  & \registerArray[2][23]~q )))

	.dataa(\Mux8~14_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\registerArray[2][23]~q ),
	.cin(gnd),
	.combout(\Mux8~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~15 .lut_mask = 16'hBAAA;
defparam \Mux8~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N14
cycloneive_lcell_comb \Mux8~17 (
// Equation(s):
// \Mux8~17_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[13][23]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[12][23]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][23]~q ),
	.datad(\registerArray[13][23]~q ),
	.cin(gnd),
	.combout(\Mux8~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~17 .lut_mask = 16'hDC98;
defparam \Mux8~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N14
cycloneive_lcell_comb \Mux7~2 (
// Equation(s):
// \Mux7~2_combout  = (\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o ) # ((\registerArray[26][24]~q )))) # (!\my_rf.rsel1[3]~input_o  & (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][24]~q )))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][24]~q ),
	.datad(\registerArray[26][24]~q ),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~2 .lut_mask = 16'hBA98;
defparam \Mux7~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y37_N26
cycloneive_lcell_comb \Mux7~3 (
// Equation(s):
// \Mux7~3_combout  = (\Mux7~2_combout  & (((\registerArray[30][24]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux7~2_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[22][24]~q ))))

	.dataa(\Mux7~2_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[30][24]~q ),
	.datad(\registerArray[22][24]~q ),
	.cin(gnd),
	.combout(\Mux7~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~3 .lut_mask = 16'hE6A2;
defparam \Mux7~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N28
cycloneive_lcell_comb \Mux7~4 (
// Equation(s):
// \Mux7~4_combout  = (\my_rf.rsel1[3]~input_o  & ((\registerArray[24][24]~q ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((\registerArray[16][24]~q  & !\my_rf.rsel1[2]~input_o ))))

	.dataa(\registerArray[24][24]~q ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[16][24]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux7~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~4 .lut_mask = 16'hCCB8;
defparam \Mux7~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N16
cycloneive_lcell_comb \Mux7~5 (
// Equation(s):
// \Mux7~5_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux7~4_combout  & (\registerArray[28][24]~q )) # (!\Mux7~4_combout  & ((\registerArray[20][24]~q ))))) # (!\my_rf.rsel1[2]~input_o  & (\Mux7~4_combout ))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux7~4_combout ),
	.datac(\registerArray[28][24]~q ),
	.datad(\registerArray[20][24]~q ),
	.cin(gnd),
	.combout(\Mux7~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~5 .lut_mask = 16'hE6C4;
defparam \Mux7~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N30
cycloneive_lcell_comb \Mux7~6 (
// Equation(s):
// \Mux7~6_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o ) # (\Mux7~3_combout )))) # (!\my_rf.rsel1[1]~input_o  & (\Mux7~5_combout  & (!\my_rf.rsel1[0]~input_o )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\Mux7~5_combout ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\Mux7~3_combout ),
	.cin(gnd),
	.combout(\Mux7~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~6 .lut_mask = 16'hAEA4;
defparam \Mux7~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N14
cycloneive_lcell_comb \Mux7~7 (
// Equation(s):
// \Mux7~7_combout  = (\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o ) # ((\registerArray[23][24]~q )))) # (!\my_rf.rsel1[2]~input_o  & (!\my_rf.rsel1[3]~input_o  & (\registerArray[19][24]~q )))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[19][24]~q ),
	.datad(\registerArray[23][24]~q ),
	.cin(gnd),
	.combout(\Mux7~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~7 .lut_mask = 16'hBA98;
defparam \Mux7~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N26
cycloneive_lcell_comb \Mux7~10 (
// Equation(s):
// \Mux7~10_combout  = (\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o )) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[10][24]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[8][24]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[8][24]~q ),
	.datad(\registerArray[10][24]~q ),
	.cin(gnd),
	.combout(\Mux7~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~10 .lut_mask = 16'hDC98;
defparam \Mux7~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N20
cycloneive_lcell_comb \Mux7~12 (
// Equation(s):
// \Mux7~12_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[5][24]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[4][24]~q )))))

	.dataa(\registerArray[5][24]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[4][24]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux7~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~12 .lut_mask = 16'hEE30;
defparam \Mux7~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N18
cycloneive_lcell_comb \Mux7~17 (
// Equation(s):
// \Mux7~17_combout  = (\my_rf.rsel1[0]~input_o  & ((\registerArray[13][24]~q ) # ((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & (((\registerArray[12][24]~q  & !\my_rf.rsel1[1]~input_o ))))

	.dataa(\registerArray[13][24]~q ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][24]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux7~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~17 .lut_mask = 16'hCCB8;
defparam \Mux7~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N26
cycloneive_lcell_comb \Mux6~2 (
// Equation(s):
// \Mux6~2_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[22][25]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][25]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][25]~q ),
	.datad(\registerArray[22][25]~q ),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~2 .lut_mask = 16'hDC98;
defparam \Mux6~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N28
cycloneive_lcell_comb \Mux6~4 (
// Equation(s):
// \Mux6~4_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[20][25]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[16][25]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[16][25]~q ),
	.datad(\registerArray[20][25]~q ),
	.cin(gnd),
	.combout(\Mux6~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~4 .lut_mask = 16'hDC98;
defparam \Mux6~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N14
cycloneive_lcell_comb \Mux6~10 (
// Equation(s):
// \Mux6~10_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[5][25]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[4][25]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[4][25]~q ),
	.datad(\registerArray[5][25]~q ),
	.cin(gnd),
	.combout(\Mux6~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~10 .lut_mask = 16'hDC98;
defparam \Mux6~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N6
cycloneive_lcell_comb \Mux6~12 (
// Equation(s):
// \Mux6~12_combout  = (\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o )) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[10][25]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[8][25]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[8][25]~q ),
	.datad(\registerArray[10][25]~q ),
	.cin(gnd),
	.combout(\Mux6~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~12 .lut_mask = 16'hDC98;
defparam \Mux6~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N22
cycloneive_lcell_comb \Mux6~13 (
// Equation(s):
// \Mux6~13_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux6~12_combout  & (\registerArray[11][25]~q )) # (!\Mux6~12_combout  & ((\registerArray[9][25]~q ))))) # (!\my_rf.rsel1[0]~input_o  & (\Mux6~12_combout ))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux6~12_combout ),
	.datac(\registerArray[11][25]~q ),
	.datad(\registerArray[9][25]~q ),
	.cin(gnd),
	.combout(\Mux6~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~13 .lut_mask = 16'hE6C4;
defparam \Mux6~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N6
cycloneive_lcell_comb \Mux6~17 (
// Equation(s):
// \Mux6~17_combout  = (\my_rf.rsel1[0]~input_o  & ((\registerArray[13][25]~q ) # ((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & (((\registerArray[12][25]~q  & !\my_rf.rsel1[1]~input_o ))))

	.dataa(\registerArray[13][25]~q ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][25]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux6~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~17 .lut_mask = 16'hCCB8;
defparam \Mux6~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N2
cycloneive_lcell_comb \Mux6~18 (
// Equation(s):
// \Mux6~18_combout  = (\Mux6~17_combout  & (((\registerArray[15][25]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux6~17_combout  & (\registerArray[14][25]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux6~17_combout ),
	.datab(\registerArray[14][25]~q ),
	.datac(\registerArray[15][25]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux6~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~18 .lut_mask = 16'hE4AA;
defparam \Mux6~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N16
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// \Mux5~0_combout  = (\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o ) # ((\registerArray[21][26]~q )))) # (!\my_rf.rsel1[2]~input_o  & (!\my_rf.rsel1[3]~input_o  & (\registerArray[17][26]~q )))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[17][26]~q ),
	.datad(\registerArray[21][26]~q ),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'hBA98;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N26
cycloneive_lcell_comb \Mux5~1 (
// Equation(s):
// \Mux5~1_combout  = (\Mux5~0_combout  & (((\registerArray[29][26]~q ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux5~0_combout  & (\registerArray[25][26]~q  & ((\my_rf.rsel1[3]~input_o ))))

	.dataa(\registerArray[25][26]~q ),
	.datab(\Mux5~0_combout ),
	.datac(\registerArray[29][26]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~1 .lut_mask = 16'hE2CC;
defparam \Mux5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N30
cycloneive_lcell_comb \Mux5~2 (
// Equation(s):
// \Mux5~2_combout  = (\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o ) # ((\registerArray[26][26]~q )))) # (!\my_rf.rsel1[3]~input_o  & (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][26]~q )))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][26]~q ),
	.datad(\registerArray[26][26]~q ),
	.cin(gnd),
	.combout(\Mux5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~2 .lut_mask = 16'hBA98;
defparam \Mux5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N2
cycloneive_lcell_comb \Mux5~3 (
// Equation(s):
// \Mux5~3_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux5~2_combout  & ((\registerArray[30][26]~q ))) # (!\Mux5~2_combout  & (\registerArray[22][26]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux5~2_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[22][26]~q ),
	.datac(\registerArray[30][26]~q ),
	.datad(\Mux5~2_combout ),
	.cin(gnd),
	.combout(\Mux5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~3 .lut_mask = 16'hF588;
defparam \Mux5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N24
cycloneive_lcell_comb \Mux5~4 (
// Equation(s):
// \Mux5~4_combout  = (\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o ) # ((\registerArray[24][26]~q )))) # (!\my_rf.rsel1[3]~input_o  & (!\my_rf.rsel1[2]~input_o  & (\registerArray[16][26]~q )))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[16][26]~q ),
	.datad(\registerArray[24][26]~q ),
	.cin(gnd),
	.combout(\Mux5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~4 .lut_mask = 16'hBA98;
defparam \Mux5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N4
cycloneive_lcell_comb \Mux5~7 (
// Equation(s):
// \Mux5~7_combout  = (\my_rf.rsel1[2]~input_o  & ((\registerArray[23][26]~q ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\registerArray[19][26]~q  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[23][26]~q ),
	.datac(\registerArray[19][26]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux5~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~7 .lut_mask = 16'hAAD8;
defparam \Mux5~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N18
cycloneive_lcell_comb \Mux5~10 (
// Equation(s):
// \Mux5~10_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\registerArray[10][26]~q )) # (!\my_rf.rsel1[1]~input_o  & ((\registerArray[8][26]~q )))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\registerArray[10][26]~q ),
	.datac(\registerArray[8][26]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux5~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~10 .lut_mask = 16'hEE50;
defparam \Mux5~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N10
cycloneive_lcell_comb \Mux5~11 (
// Equation(s):
// \Mux5~11_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux5~10_combout  & ((\registerArray[11][26]~q ))) # (!\Mux5~10_combout  & (\registerArray[9][26]~q )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux5~10_combout ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\registerArray[9][26]~q ),
	.datac(\registerArray[11][26]~q ),
	.datad(\Mux5~10_combout ),
	.cin(gnd),
	.combout(\Mux5~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~11 .lut_mask = 16'hF588;
defparam \Mux5~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N26
cycloneive_lcell_comb \Mux5~12 (
// Equation(s):
// \Mux5~12_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[5][26]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[4][26]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[4][26]~q ),
	.datad(\registerArray[5][26]~q ),
	.cin(gnd),
	.combout(\Mux5~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~12 .lut_mask = 16'hDC98;
defparam \Mux5~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N26
cycloneive_lcell_comb \Mux5~17 (
// Equation(s):
// \Mux5~17_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[13][26]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[12][26]~q )))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[13][26]~q ),
	.datac(\registerArray[12][26]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux5~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~17 .lut_mask = 16'hEE50;
defparam \Mux5~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N10
cycloneive_lcell_comb \Mux4~2 (
// Equation(s):
// \Mux4~2_combout  = (\my_rf.rsel1[2]~input_o  & ((\registerArray[22][27]~q ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\registerArray[18][27]~q  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\registerArray[22][27]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][27]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~2 .lut_mask = 16'hCCB8;
defparam \Mux4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N28
cycloneive_lcell_comb \Mux4~3 (
// Equation(s):
// \Mux4~3_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux4~2_combout  & ((\registerArray[30][27]~q ))) # (!\Mux4~2_combout  & (\registerArray[26][27]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux4~2_combout ))))

	.dataa(\registerArray[26][27]~q ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[30][27]~q ),
	.datad(\Mux4~2_combout ),
	.cin(gnd),
	.combout(\Mux4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~3 .lut_mask = 16'hF388;
defparam \Mux4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N16
cycloneive_lcell_comb \Mux4~4 (
// Equation(s):
// \Mux4~4_combout  = (\my_rf.rsel1[2]~input_o  & ((\registerArray[20][27]~q ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\registerArray[16][27]~q  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\registerArray[20][27]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[16][27]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~4 .lut_mask = 16'hCCB8;
defparam \Mux4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N20
cycloneive_lcell_comb \Mux4~5 (
// Equation(s):
// \Mux4~5_combout  = (\Mux4~4_combout  & (((\registerArray[28][27]~q )) # (!\my_rf.rsel1[3]~input_o ))) # (!\Mux4~4_combout  & (\my_rf.rsel1[3]~input_o  & ((\registerArray[24][27]~q ))))

	.dataa(\Mux4~4_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[28][27]~q ),
	.datad(\registerArray[24][27]~q ),
	.cin(gnd),
	.combout(\Mux4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~5 .lut_mask = 16'hE6A2;
defparam \Mux4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N26
cycloneive_lcell_comb \Mux4~6 (
// Equation(s):
// \Mux4~6_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o ) # (\Mux4~3_combout )))) # (!\my_rf.rsel1[1]~input_o  & (\Mux4~5_combout  & (!\my_rf.rsel1[0]~input_o )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\Mux4~5_combout ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\Mux4~3_combout ),
	.cin(gnd),
	.combout(\Mux4~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~6 .lut_mask = 16'hAEA4;
defparam \Mux4~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N22
cycloneive_lcell_comb \Mux4~12 (
// Equation(s):
// \Mux4~12_combout  = (\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o )) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[10][27]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[8][27]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[8][27]~q ),
	.datad(\registerArray[10][27]~q ),
	.cin(gnd),
	.combout(\Mux4~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~12 .lut_mask = 16'hDC98;
defparam \Mux4~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N26
cycloneive_lcell_comb \Mux4~13 (
// Equation(s):
// \Mux4~13_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux4~12_combout  & (\registerArray[11][27]~q )) # (!\Mux4~12_combout  & ((\registerArray[9][27]~q ))))) # (!\my_rf.rsel1[0]~input_o  & (\Mux4~12_combout ))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux4~12_combout ),
	.datac(\registerArray[11][27]~q ),
	.datad(\registerArray[9][27]~q ),
	.cin(gnd),
	.combout(\Mux4~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~13 .lut_mask = 16'hE6C4;
defparam \Mux4~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N26
cycloneive_lcell_comb \Mux3~7 (
// Equation(s):
// \Mux3~7_combout  = (\my_rf.rsel1[2]~input_o  & ((\registerArray[23][28]~q ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\registerArray[19][28]~q  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[23][28]~q ),
	.datac(\registerArray[19][28]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux3~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~7 .lut_mask = 16'hAAD8;
defparam \Mux3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N14
cycloneive_lcell_comb \Mux3~8 (
// Equation(s):
// \Mux3~8_combout  = (\Mux3~7_combout  & (((\registerArray[31][28]~q )) # (!\my_rf.rsel1[3]~input_o ))) # (!\Mux3~7_combout  & (\my_rf.rsel1[3]~input_o  & ((\registerArray[27][28]~q ))))

	.dataa(\Mux3~7_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[31][28]~q ),
	.datad(\registerArray[27][28]~q ),
	.cin(gnd),
	.combout(\Mux3~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~8 .lut_mask = 16'hE6A2;
defparam \Mux3~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N2
cycloneive_lcell_comb \Mux3~10 (
// Equation(s):
// \Mux3~10_combout  = (\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o )) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[10][28]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[8][28]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[8][28]~q ),
	.datad(\registerArray[10][28]~q ),
	.cin(gnd),
	.combout(\Mux3~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~10 .lut_mask = 16'hDC98;
defparam \Mux3~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N0
cycloneive_lcell_comb \Mux3~12 (
// Equation(s):
// \Mux3~12_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[5][28]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[4][28]~q )))))

	.dataa(\registerArray[5][28]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[4][28]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux3~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~12 .lut_mask = 16'hEE30;
defparam \Mux3~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N14
cycloneive_lcell_comb \Mux3~13 (
// Equation(s):
// \Mux3~13_combout  = (\Mux3~12_combout  & (((\registerArray[7][28]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux3~12_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[6][28]~q ))))

	.dataa(\Mux3~12_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[7][28]~q ),
	.datad(\registerArray[6][28]~q ),
	.cin(gnd),
	.combout(\Mux3~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~13 .lut_mask = 16'hE6A2;
defparam \Mux3~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N18
cycloneive_lcell_comb \Mux3~14 (
// Equation(s):
// \Mux3~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\registerArray[3][28]~q )) # (!\my_rf.rsel1[1]~input_o  & ((\registerArray[1][28]~q )))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\registerArray[3][28]~q ),
	.datac(\registerArray[1][28]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux3~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~14 .lut_mask = 16'h88A0;
defparam \Mux3~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N10
cycloneive_lcell_comb \Mux3~17 (
// Equation(s):
// \Mux3~17_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[13][28]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[12][28]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][28]~q ),
	.datad(\registerArray[13][28]~q ),
	.cin(gnd),
	.combout(\Mux3~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~17 .lut_mask = 16'hDC98;
defparam \Mux3~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y34_N18
cycloneive_lcell_comb \Mux3~18 (
// Equation(s):
// \Mux3~18_combout  = (\Mux3~17_combout  & (((\registerArray[15][28]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux3~17_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[14][28]~q ))))

	.dataa(\Mux3~17_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][28]~q ),
	.datad(\registerArray[14][28]~q ),
	.cin(gnd),
	.combout(\Mux3~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~18 .lut_mask = 16'hE6A2;
defparam \Mux3~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N6
cycloneive_lcell_comb \Mux2~2 (
// Equation(s):
// \Mux2~2_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[22][29]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][29]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][29]~q ),
	.datad(\registerArray[22][29]~q ),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~2 .lut_mask = 16'hDC98;
defparam \Mux2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N4
cycloneive_lcell_comb \Mux2~3 (
// Equation(s):
// \Mux2~3_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux2~2_combout  & (\registerArray[30][29]~q )) # (!\Mux2~2_combout  & ((\registerArray[26][29]~q ))))) # (!\my_rf.rsel1[3]~input_o  & (\Mux2~2_combout ))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux2~2_combout ),
	.datac(\registerArray[30][29]~q ),
	.datad(\registerArray[26][29]~q ),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~3 .lut_mask = 16'hE6C4;
defparam \Mux2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N2
cycloneive_lcell_comb \Mux2~7 (
// Equation(s):
// \Mux2~7_combout  = (\my_rf.rsel1[2]~input_o  & (\my_rf.rsel1[3]~input_o )) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & ((\registerArray[27][29]~q ))) # (!\my_rf.rsel1[3]~input_o  & (\registerArray[19][29]~q ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[19][29]~q ),
	.datad(\registerArray[27][29]~q ),
	.cin(gnd),
	.combout(\Mux2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~7 .lut_mask = 16'hDC98;
defparam \Mux2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N4
cycloneive_lcell_comb \Mux2~8 (
// Equation(s):
// \Mux2~8_combout  = (\Mux2~7_combout  & (((\registerArray[31][29]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux2~7_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[23][29]~q ))))

	.dataa(\Mux2~7_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[31][29]~q ),
	.datad(\registerArray[23][29]~q ),
	.cin(gnd),
	.combout(\Mux2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~8 .lut_mask = 16'hE6A2;
defparam \Mux2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N10
cycloneive_lcell_comb \Mux2~10 (
// Equation(s):
// \Mux2~10_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[5][29]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[4][29]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[4][29]~q ),
	.datad(\registerArray[5][29]~q ),
	.cin(gnd),
	.combout(\Mux2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~10 .lut_mask = 16'hDC98;
defparam \Mux2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N14
cycloneive_lcell_comb \Mux2~12 (
// Equation(s):
// \Mux2~12_combout  = (\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o )) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[10][29]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[8][29]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[8][29]~q ),
	.datad(\registerArray[10][29]~q ),
	.cin(gnd),
	.combout(\Mux2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~12 .lut_mask = 16'hDC98;
defparam \Mux2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N20
cycloneive_lcell_comb \Mux2~13 (
// Equation(s):
// \Mux2~13_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux2~12_combout  & (\registerArray[11][29]~q )) # (!\Mux2~12_combout  & ((\registerArray[9][29]~q ))))) # (!\my_rf.rsel1[0]~input_o  & (\Mux2~12_combout ))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux2~12_combout ),
	.datac(\registerArray[11][29]~q ),
	.datad(\registerArray[9][29]~q ),
	.cin(gnd),
	.combout(\Mux2~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~13 .lut_mask = 16'hE6C4;
defparam \Mux2~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N30
cycloneive_lcell_comb \Mux2~17 (
// Equation(s):
// \Mux2~17_combout  = (\my_rf.rsel1[0]~input_o  & ((\registerArray[13][29]~q ) # ((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & (((\registerArray[12][29]~q  & !\my_rf.rsel1[1]~input_o ))))

	.dataa(\registerArray[13][29]~q ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][29]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux2~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~17 .lut_mask = 16'hCCB8;
defparam \Mux2~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N30
cycloneive_lcell_comb \Mux2~18 (
// Equation(s):
// \Mux2~18_combout  = (\Mux2~17_combout  & (((\registerArray[15][29]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux2~17_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[14][29]~q ))))

	.dataa(\Mux2~17_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][29]~q ),
	.datad(\registerArray[14][29]~q ),
	.cin(gnd),
	.combout(\Mux2~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~18 .lut_mask = 16'hE6A2;
defparam \Mux2~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N14
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// \Mux1~0_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[21][30]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[17][30]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[17][30]~q ),
	.datad(\registerArray[21][30]~q ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'hDC98;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N6
cycloneive_lcell_comb \Mux1~2 (
// Equation(s):
// \Mux1~2_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[26][30]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[18][30]~q )))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[26][30]~q ),
	.datac(\registerArray[18][30]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~2 .lut_mask = 16'hEE50;
defparam \Mux1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N24
cycloneive_lcell_comb \Mux1~3 (
// Equation(s):
// \Mux1~3_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux1~2_combout  & (\registerArray[30][30]~q )) # (!\Mux1~2_combout  & ((\registerArray[22][30]~q ))))) # (!\my_rf.rsel1[2]~input_o  & (\Mux1~2_combout ))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux1~2_combout ),
	.datac(\registerArray[30][30]~q ),
	.datad(\registerArray[22][30]~q ),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~3 .lut_mask = 16'hE6C4;
defparam \Mux1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N20
cycloneive_lcell_comb \Mux1~4 (
// Equation(s):
// \Mux1~4_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[24][30]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[16][30]~q )))))

	.dataa(\registerArray[24][30]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[16][30]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~4 .lut_mask = 16'hEE30;
defparam \Mux1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N10
cycloneive_lcell_comb \Mux1~5 (
// Equation(s):
// \Mux1~5_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux1~4_combout  & (\registerArray[28][30]~q )) # (!\Mux1~4_combout  & ((\registerArray[20][30]~q ))))) # (!\my_rf.rsel1[2]~input_o  & (\Mux1~4_combout ))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux1~4_combout ),
	.datac(\registerArray[28][30]~q ),
	.datad(\registerArray[20][30]~q ),
	.cin(gnd),
	.combout(\Mux1~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~5 .lut_mask = 16'hE6C4;
defparam \Mux1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N6
cycloneive_lcell_comb \Mux1~6 (
// Equation(s):
// \Mux1~6_combout  = (\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o )) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\Mux1~3_combout )) # (!\my_rf.rsel1[1]~input_o  & ((\Mux1~5_combout )))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\Mux1~3_combout ),
	.datad(\Mux1~5_combout ),
	.cin(gnd),
	.combout(\Mux1~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~6 .lut_mask = 16'hD9C8;
defparam \Mux1~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N14
cycloneive_lcell_comb \Mux1~10 (
// Equation(s):
// \Mux1~10_combout  = (\my_rf.rsel1[1]~input_o  & ((\registerArray[10][30]~q ) # ((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & (((\registerArray[8][30]~q  & !\my_rf.rsel1[0]~input_o ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[10][30]~q ),
	.datac(\registerArray[8][30]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~10 .lut_mask = 16'hAAD8;
defparam \Mux1~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N30
cycloneive_lcell_comb \Mux1~11 (
// Equation(s):
// \Mux1~11_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux1~10_combout  & ((\registerArray[11][30]~q ))) # (!\Mux1~10_combout  & (\registerArray[9][30]~q )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux1~10_combout ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\registerArray[9][30]~q ),
	.datac(\registerArray[11][30]~q ),
	.datad(\Mux1~10_combout ),
	.cin(gnd),
	.combout(\Mux1~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~11 .lut_mask = 16'hF588;
defparam \Mux1~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N12
cycloneive_lcell_comb \Mux1~12 (
// Equation(s):
// \Mux1~12_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[5][30]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[4][30]~q )))))

	.dataa(\registerArray[5][30]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[4][30]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux1~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~12 .lut_mask = 16'hEE30;
defparam \Mux1~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N2
cycloneive_lcell_comb \Mux1~14 (
// Equation(s):
// \Mux1~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][30]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][30]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[1][30]~q ),
	.datad(\registerArray[3][30]~q ),
	.cin(gnd),
	.combout(\Mux1~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~14 .lut_mask = 16'hC840;
defparam \Mux1~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N26
cycloneive_lcell_comb \Mux1~15 (
// Equation(s):
// \Mux1~15_combout  = (\Mux1~14_combout ) # ((!\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o  & \registerArray[2][30]~q )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\Mux1~14_combout ),
	.datad(\registerArray[2][30]~q ),
	.cin(gnd),
	.combout(\Mux1~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~15 .lut_mask = 16'hF4F0;
defparam \Mux1~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N14
cycloneive_lcell_comb \Mux1~17 (
// Equation(s):
// \Mux1~17_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[13][30]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[12][30]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][30]~q ),
	.datad(\registerArray[13][30]~q ),
	.cin(gnd),
	.combout(\Mux1~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~17 .lut_mask = 16'hDC98;
defparam \Mux1~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N8
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// \Mux0~0_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[25][31]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[17][31]~q )))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[25][31]~q ),
	.datac(\registerArray[17][31]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'hEE50;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N26
cycloneive_lcell_comb \Mux0~1 (
// Equation(s):
// \Mux0~1_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux0~0_combout  & (\registerArray[29][31]~q )) # (!\Mux0~0_combout  & ((\registerArray[21][31]~q ))))) # (!\my_rf.rsel1[2]~input_o  & (\Mux0~0_combout ))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux0~0_combout ),
	.datac(\registerArray[29][31]~q ),
	.datad(\registerArray[21][31]~q ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~1 .lut_mask = 16'hE6C4;
defparam \Mux0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N6
cycloneive_lcell_comb \Mux0~2 (
// Equation(s):
// \Mux0~2_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[22][31]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][31]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][31]~q ),
	.datad(\registerArray[22][31]~q ),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~2 .lut_mask = 16'hDC98;
defparam \Mux0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N8
cycloneive_lcell_comb \Mux0~3 (
// Equation(s):
// \Mux0~3_combout  = (\Mux0~2_combout  & (((\registerArray[30][31]~q ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux0~2_combout  & (\registerArray[26][31]~q  & ((\my_rf.rsel1[3]~input_o ))))

	.dataa(\Mux0~2_combout ),
	.datab(\registerArray[26][31]~q ),
	.datac(\registerArray[30][31]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~3 .lut_mask = 16'hE4AA;
defparam \Mux0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N6
cycloneive_lcell_comb \Mux0~7 (
// Equation(s):
// \Mux0~7_combout  = (\my_rf.rsel1[3]~input_o  & ((\registerArray[27][31]~q ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((\registerArray[19][31]~q  & !\my_rf.rsel1[2]~input_o ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[27][31]~q ),
	.datac(\registerArray[19][31]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~7 .lut_mask = 16'hAAD8;
defparam \Mux0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y37_N22
cycloneive_lcell_comb \Mux0~12 (
// Equation(s):
// \Mux0~12_combout  = (\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o )) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[10][31]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[8][31]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[8][31]~q ),
	.datad(\registerArray[10][31]~q ),
	.cin(gnd),
	.combout(\Mux0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~12 .lut_mask = 16'hDC98;
defparam \Mux0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y37_N22
cycloneive_lcell_comb \Mux0~13 (
// Equation(s):
// \Mux0~13_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux0~12_combout  & ((\registerArray[11][31]~q ))) # (!\Mux0~12_combout  & (\registerArray[9][31]~q )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux0~12_combout ))))

	.dataa(\registerArray[9][31]~q ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[11][31]~q ),
	.datad(\Mux0~12_combout ),
	.cin(gnd),
	.combout(\Mux0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~13 .lut_mask = 16'hF388;
defparam \Mux0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N30
cycloneive_lcell_comb \Mux0~14 (
// Equation(s):
// \Mux0~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][31]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][31]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[1][31]~q ),
	.datad(\registerArray[3][31]~q ),
	.cin(gnd),
	.combout(\Mux0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~14 .lut_mask = 16'hC840;
defparam \Mux0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y36_N2
cycloneive_lcell_comb \Mux0~17 (
// Equation(s):
// \Mux0~17_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[13][31]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[12][31]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][31]~q ),
	.datad(\registerArray[13][31]~q ),
	.cin(gnd),
	.combout(\Mux0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~17 .lut_mask = 16'hDC98;
defparam \Mux0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N12
cycloneive_lcell_comb \Mux0~18 (
// Equation(s):
// \Mux0~18_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux0~17_combout  & ((\registerArray[15][31]~q ))) # (!\Mux0~17_combout  & (\registerArray[14][31]~q )))) # (!\my_rf.rsel1[1]~input_o  & (((\Mux0~17_combout ))))

	.dataa(\registerArray[14][31]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][31]~q ),
	.datad(\Mux0~17_combout ),
	.cin(gnd),
	.combout(\Mux0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~18 .lut_mask = 16'hF388;
defparam \Mux0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N8
cycloneive_io_ibuf \clk~input (
	.i(clk),
	.ibar(gnd),
	.o(\clk~input_o ));
// synopsys translate_off
defparam \clk~input .bus_hold = "false";
defparam \clk~input .simulate_z_as = "z";
// synopsys translate_on

// Location: CLKCTRL_G2
cycloneive_clkctrl \clk~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\clk~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\clk~inputclkctrl_outclk ));
// synopsys translate_off
defparam \clk~inputclkctrl .clock_type = "global clock";
defparam \clk~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: IOOBUF_X52_Y73_N2
cycloneive_io_obuf \my_rf.rdat2[0]~output (
	.i(\Mux63~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [0]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[0]~output .bus_hold = "false";
defparam \my_rf.rdat2[0]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N16
cycloneive_io_obuf \my_rf.rdat2[1]~output (
	.i(\Mux62~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [1]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[1]~output .bus_hold = "false";
defparam \my_rf.rdat2[1]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N23
cycloneive_io_obuf \my_rf.rdat2[2]~output (
	.i(\Mux61~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [2]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[2]~output .bus_hold = "false";
defparam \my_rf.rdat2[2]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y43_N16
cycloneive_io_obuf \my_rf.rdat2[3]~output (
	.i(\Mux60~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [3]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[3]~output .bus_hold = "false";
defparam \my_rf.rdat2[3]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y0_N23
cycloneive_io_obuf \my_rf.rdat2[4]~output (
	.i(\Mux59~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [4]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[4]~output .bus_hold = "false";
defparam \my_rf.rdat2[4]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y27_N16
cycloneive_io_obuf \my_rf.rdat2[5]~output (
	.i(\Mux58~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [5]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[5]~output .bus_hold = "false";
defparam \my_rf.rdat2[5]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X58_Y73_N9
cycloneive_io_obuf \my_rf.rdat2[6]~output (
	.i(\Mux57~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [6]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[6]~output .bus_hold = "false";
defparam \my_rf.rdat2[6]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X58_Y73_N16
cycloneive_io_obuf \my_rf.rdat2[7]~output (
	.i(\Mux56~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [7]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[7]~output .bus_hold = "false";
defparam \my_rf.rdat2[7]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y73_N2
cycloneive_io_obuf \my_rf.rdat2[8]~output (
	.i(\Mux55~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [8]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[8]~output .bus_hold = "false";
defparam \my_rf.rdat2[8]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N2
cycloneive_io_obuf \my_rf.rdat2[9]~output (
	.i(\Mux54~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [9]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[9]~output .bus_hold = "false";
defparam \my_rf.rdat2[9]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y42_N9
cycloneive_io_obuf \my_rf.rdat2[10]~output (
	.i(\Mux53~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [10]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[10]~output .bus_hold = "false";
defparam \my_rf.rdat2[10]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y73_N9
cycloneive_io_obuf \my_rf.rdat2[11]~output (
	.i(\Mux52~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [11]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[11]~output .bus_hold = "false";
defparam \my_rf.rdat2[11]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N23
cycloneive_io_obuf \my_rf.rdat2[12]~output (
	.i(\Mux51~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [12]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[12]~output .bus_hold = "false";
defparam \my_rf.rdat2[12]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N2
cycloneive_io_obuf \my_rf.rdat2[13]~output (
	.i(\Mux50~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [13]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[13]~output .bus_hold = "false";
defparam \my_rf.rdat2[13]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X35_Y0_N23
cycloneive_io_obuf \my_rf.rdat2[14]~output (
	.i(\Mux49~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [14]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[14]~output .bus_hold = "false";
defparam \my_rf.rdat2[14]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X38_Y73_N23
cycloneive_io_obuf \my_rf.rdat2[15]~output (
	.i(\Mux48~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [15]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[15]~output .bus_hold = "false";
defparam \my_rf.rdat2[15]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y44_N2
cycloneive_io_obuf \my_rf.rdat2[16]~output (
	.i(\Mux47~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [16]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[16]~output .bus_hold = "false";
defparam \my_rf.rdat2[16]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X33_Y73_N9
cycloneive_io_obuf \my_rf.rdat2[17]~output (
	.i(\Mux46~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [17]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[17]~output .bus_hold = "false";
defparam \my_rf.rdat2[17]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X31_Y0_N9
cycloneive_io_obuf \my_rf.rdat2[18]~output (
	.i(\Mux45~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [18]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[18]~output .bus_hold = "false";
defparam \my_rf.rdat2[18]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y73_N16
cycloneive_io_obuf \my_rf.rdat2[19]~output (
	.i(\Mux44~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [19]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[19]~output .bus_hold = "false";
defparam \my_rf.rdat2[19]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y44_N9
cycloneive_io_obuf \my_rf.rdat2[20]~output (
	.i(\Mux43~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [20]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[20]~output .bus_hold = "false";
defparam \my_rf.rdat2[20]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y25_N23
cycloneive_io_obuf \my_rf.rdat2[21]~output (
	.i(\Mux42~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [21]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[21]~output .bus_hold = "false";
defparam \my_rf.rdat2[21]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X35_Y0_N16
cycloneive_io_obuf \my_rf.rdat2[22]~output (
	.i(\Mux41~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [22]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[22]~output .bus_hold = "false";
defparam \my_rf.rdat2[22]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y24_N9
cycloneive_io_obuf \my_rf.rdat2[23]~output (
	.i(\Mux40~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [23]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[23]~output .bus_hold = "false";
defparam \my_rf.rdat2[23]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N16
cycloneive_io_obuf \my_rf.rdat2[24]~output (
	.i(\Mux39~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [24]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[24]~output .bus_hold = "false";
defparam \my_rf.rdat2[24]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X33_Y0_N9
cycloneive_io_obuf \my_rf.rdat2[25]~output (
	.i(\Mux38~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [25]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[25]~output .bus_hold = "false";
defparam \my_rf.rdat2[25]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X38_Y73_N9
cycloneive_io_obuf \my_rf.rdat2[26]~output (
	.i(\Mux37~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [26]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[26]~output .bus_hold = "false";
defparam \my_rf.rdat2[26]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y30_N2
cycloneive_io_obuf \my_rf.rdat2[27]~output (
	.i(\Mux36~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [27]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[27]~output .bus_hold = "false";
defparam \my_rf.rdat2[27]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X38_Y73_N16
cycloneive_io_obuf \my_rf.rdat2[28]~output (
	.i(\Mux35~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [28]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[28]~output .bus_hold = "false";
defparam \my_rf.rdat2[28]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X42_Y73_N9
cycloneive_io_obuf \my_rf.rdat2[29]~output (
	.i(\Mux34~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [29]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[29]~output .bus_hold = "false";
defparam \my_rf.rdat2[29]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y46_N16
cycloneive_io_obuf \my_rf.rdat2[30]~output (
	.i(\Mux33~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [30]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[30]~output .bus_hold = "false";
defparam \my_rf.rdat2[30]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X40_Y73_N9
cycloneive_io_obuf \my_rf.rdat2[31]~output (
	.i(\Mux32~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat2 [31]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat2[31]~output .bus_hold = "false";
defparam \my_rf.rdat2[31]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X58_Y73_N2
cycloneive_io_obuf \my_rf.rdat1[0]~output (
	.i(\Mux31~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [0]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[0]~output .bus_hold = "false";
defparam \my_rf.rdat1[0]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y45_N16
cycloneive_io_obuf \my_rf.rdat1[1]~output (
	.i(\Mux30~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [1]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[1]~output .bus_hold = "false";
defparam \my_rf.rdat1[1]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y0_N16
cycloneive_io_obuf \my_rf.rdat1[2]~output (
	.i(\Mux29~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [2]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[2]~output .bus_hold = "false";
defparam \my_rf.rdat1[2]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X49_Y73_N16
cycloneive_io_obuf \my_rf.rdat1[3]~output (
	.i(\Mux28~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [3]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[3]~output .bus_hold = "false";
defparam \my_rf.rdat1[3]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X29_Y0_N16
cycloneive_io_obuf \my_rf.rdat1[4]~output (
	.i(\Mux27~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [4]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[4]~output .bus_hold = "false";
defparam \my_rf.rdat1[4]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y73_N9
cycloneive_io_obuf \my_rf.rdat1[5]~output (
	.i(\Mux26~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [5]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[5]~output .bus_hold = "false";
defparam \my_rf.rdat1[5]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N16
cycloneive_io_obuf \my_rf.rdat1[6]~output (
	.i(\Mux25~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [6]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[6]~output .bus_hold = "false";
defparam \my_rf.rdat1[6]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N9
cycloneive_io_obuf \my_rf.rdat1[7]~output (
	.i(\Mux24~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [7]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[7]~output .bus_hold = "false";
defparam \my_rf.rdat1[7]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X58_Y73_N23
cycloneive_io_obuf \my_rf.rdat1[8]~output (
	.i(\Mux23~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [8]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[8]~output .bus_hold = "false";
defparam \my_rf.rdat1[8]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N9
cycloneive_io_obuf \my_rf.rdat1[9]~output (
	.i(\Mux22~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [9]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[9]~output .bus_hold = "false";
defparam \my_rf.rdat1[9]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X49_Y73_N23
cycloneive_io_obuf \my_rf.rdat1[10]~output (
	.i(\Mux21~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [10]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[10]~output .bus_hold = "false";
defparam \my_rf.rdat1[10]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y36_N2
cycloneive_io_obuf \my_rf.rdat1[11]~output (
	.i(\Mux20~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [11]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[11]~output .bus_hold = "false";
defparam \my_rf.rdat1[11]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y30_N9
cycloneive_io_obuf \my_rf.rdat1[12]~output (
	.i(\Mux19~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [12]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[12]~output .bus_hold = "false";
defparam \my_rf.rdat1[12]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N9
cycloneive_io_obuf \my_rf.rdat1[13]~output (
	.i(\Mux18~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [13]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[13]~output .bus_hold = "false";
defparam \my_rf.rdat1[13]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y45_N23
cycloneive_io_obuf \my_rf.rdat1[14]~output (
	.i(\Mux17~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [14]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[14]~output .bus_hold = "false";
defparam \my_rf.rdat1[14]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X35_Y73_N23
cycloneive_io_obuf \my_rf.rdat1[15]~output (
	.i(\Mux16~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [15]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[15]~output .bus_hold = "false";
defparam \my_rf.rdat1[15]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y27_N23
cycloneive_io_obuf \my_rf.rdat1[16]~output (
	.i(\Mux15~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [16]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[16]~output .bus_hold = "false";
defparam \my_rf.rdat1[16]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X47_Y73_N2
cycloneive_io_obuf \my_rf.rdat1[17]~output (
	.i(\Mux14~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [17]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[17]~output .bus_hold = "false";
defparam \my_rf.rdat1[17]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X45_Y73_N2
cycloneive_io_obuf \my_rf.rdat1[18]~output (
	.i(\Mux13~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [18]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[18]~output .bus_hold = "false";
defparam \my_rf.rdat1[18]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y25_N16
cycloneive_io_obuf \my_rf.rdat1[19]~output (
	.i(\Mux12~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [19]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[19]~output .bus_hold = "false";
defparam \my_rf.rdat1[19]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X27_Y0_N23
cycloneive_io_obuf \my_rf.rdat1[20]~output (
	.i(\Mux11~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [20]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[20]~output .bus_hold = "false";
defparam \my_rf.rdat1[20]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X29_Y0_N23
cycloneive_io_obuf \my_rf.rdat1[21]~output (
	.i(\Mux10~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [21]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[21]~output .bus_hold = "false";
defparam \my_rf.rdat1[21]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y44_N23
cycloneive_io_obuf \my_rf.rdat1[22]~output (
	.i(\Mux9~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [22]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[22]~output .bus_hold = "false";
defparam \my_rf.rdat1[22]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y42_N2
cycloneive_io_obuf \my_rf.rdat1[23]~output (
	.i(\Mux8~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [23]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[23]~output .bus_hold = "false";
defparam \my_rf.rdat1[23]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y26_N16
cycloneive_io_obuf \my_rf.rdat1[24]~output (
	.i(\Mux7~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [24]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[24]~output .bus_hold = "false";
defparam \my_rf.rdat1[24]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X35_Y73_N16
cycloneive_io_obuf \my_rf.rdat1[25]~output (
	.i(\Mux6~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [25]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[25]~output .bus_hold = "false";
defparam \my_rf.rdat1[25]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y44_N16
cycloneive_io_obuf \my_rf.rdat1[26]~output (
	.i(\Mux5~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [26]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[26]~output .bus_hold = "false";
defparam \my_rf.rdat1[26]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X40_Y73_N2
cycloneive_io_obuf \my_rf.rdat1[27]~output (
	.i(\Mux4~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [27]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[27]~output .bus_hold = "false";
defparam \my_rf.rdat1[27]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X38_Y73_N2
cycloneive_io_obuf \my_rf.rdat1[28]~output (
	.i(\Mux3~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [28]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[28]~output .bus_hold = "false";
defparam \my_rf.rdat1[28]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X27_Y0_N9
cycloneive_io_obuf \my_rf.rdat1[29]~output (
	.i(\Mux2~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [29]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[29]~output .bus_hold = "false";
defparam \my_rf.rdat1[29]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N16
cycloneive_io_obuf \my_rf.rdat1[30]~output (
	.i(\Mux1~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [30]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[30]~output .bus_hold = "false";
defparam \my_rf.rdat1[30]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X42_Y73_N2
cycloneive_io_obuf \my_rf.rdat1[31]~output (
	.i(\Mux0~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\my_rf.rdat1 [31]),
	.obar());
// synopsys translate_off
defparam \my_rf.rdat1[31]~output .bus_hold = "false";
defparam \my_rf.rdat1[31]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOIBUF_X0_Y35_N8
cycloneive_io_ibuf \my_rf.rsel2[4]~input (
	.i(\my_rf.rsel2 [4]),
	.ibar(gnd),
	.o(\my_rf.rsel2[4]~input_o ));
// synopsys translate_off
defparam \my_rf.rsel2[4]~input .bus_hold = "false";
defparam \my_rf.rsel2[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y28_N15
cycloneive_io_ibuf \my_rf.rsel2[3]~input (
	.i(\my_rf.rsel2 [3]),
	.ibar(gnd),
	.o(\my_rf.rsel2[3]~input_o ));
// synopsys translate_off
defparam \my_rf.rsel2[3]~input .bus_hold = "false";
defparam \my_rf.rsel2[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N22
cycloneive_io_ibuf \my_rf.rsel2[0]~input (
	.i(\my_rf.rsel2 [0]),
	.ibar(gnd),
	.o(\my_rf.rsel2[0]~input_o ));
// synopsys translate_off
defparam \my_rf.rsel2[0]~input .bus_hold = "false";
defparam \my_rf.rsel2[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X56_Y0_N22
cycloneive_io_ibuf \my_rf.wdat[0]~input (
	.i(\my_rf.wdat [0]),
	.ibar(gnd),
	.o(\my_rf.wdat[0]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[0]~input .bus_hold = "false";
defparam \my_rf.wdat[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N15
cycloneive_io_ibuf \n_rst~input (
	.i(n_rst),
	.ibar(gnd),
	.o(\n_rst~input_o ));
// synopsys translate_off
defparam \n_rst~input .bus_hold = "false";
defparam \n_rst~input .simulate_z_as = "z";
// synopsys translate_on

// Location: CLKCTRL_G4
cycloneive_clkctrl \n_rst~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\n_rst~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\n_rst~inputclkctrl_outclk ));
// synopsys translate_off
defparam \n_rst~inputclkctrl .clock_type = "global clock";
defparam \n_rst~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: IOIBUF_X31_Y0_N1
cycloneive_io_ibuf \my_rf.wsel[3]~input (
	.i(\my_rf.wsel [3]),
	.ibar(gnd),
	.o(\my_rf.wsel[3]~input_o ));
// synopsys translate_off
defparam \my_rf.wsel[3]~input .bus_hold = "false";
defparam \my_rf.wsel[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y24_N15
cycloneive_io_ibuf \my_rf.wsel[1]~input (
	.i(\my_rf.wsel [1]),
	.ibar(gnd),
	.o(\my_rf.wsel[1]~input_o ));
// synopsys translate_off
defparam \my_rf.wsel[1]~input .bus_hold = "false";
defparam \my_rf.wsel[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y31_N15
cycloneive_io_ibuf \my_rf.wsel[0]~input (
	.i(\my_rf.wsel [0]),
	.ibar(gnd),
	.o(\my_rf.wsel[0]~input_o ));
// synopsys translate_off
defparam \my_rf.wsel[0]~input .bus_hold = "false";
defparam \my_rf.wsel[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X42_Y31_N6
cycloneive_lcell_comb \Decoder0~8 (
// Equation(s):
// \Decoder0~8_combout  = (\my_rf.WEN~input_o  & (\my_rf.wsel[3]~input_o  & (\my_rf.wsel[1]~input_o  & !\my_rf.wsel[0]~input_o )))

	.dataa(\my_rf.WEN~input_o ),
	.datab(\my_rf.wsel[3]~input_o ),
	.datac(\my_rf.wsel[1]~input_o ),
	.datad(\my_rf.wsel[0]~input_o ),
	.cin(gnd),
	.combout(\Decoder0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~8 .lut_mask = 16'h0080;
defparam \Decoder0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X0_Y28_N22
cycloneive_io_ibuf \my_rf.wsel[2]~input (
	.i(\my_rf.wsel [2]),
	.ibar(gnd),
	.o(\my_rf.wsel[2]~input_o ));
// synopsys translate_off
defparam \my_rf.wsel[2]~input .bus_hold = "false";
defparam \my_rf.wsel[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X33_Y0_N1
cycloneive_io_ibuf \my_rf.wsel[4]~input (
	.i(\my_rf.wsel [4]),
	.ibar(gnd),
	.o(\my_rf.wsel[4]~input_o ));
// synopsys translate_off
defparam \my_rf.wsel[4]~input .bus_hold = "false";
defparam \my_rf.wsel[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X41_Y32_N8
cycloneive_lcell_comb \Decoder0~25 (
// Equation(s):
// \Decoder0~25_combout  = (\Decoder0~8_combout  & (!\my_rf.wsel[2]~input_o  & !\my_rf.wsel[4]~input_o ))

	.dataa(gnd),
	.datab(\Decoder0~8_combout ),
	.datac(\my_rf.wsel[2]~input_o ),
	.datad(\my_rf.wsel[4]~input_o ),
	.cin(gnd),
	.combout(\Decoder0~25_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~25 .lut_mask = 16'h000C;
defparam \Decoder0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y31_N1
dffeas \registerArray[10][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][0] .is_wysiwyg = "true";
defparam \registerArray[10][0] .power_up = "low";
// synopsys translate_on

// Location: IOIBUF_X0_Y24_N1
cycloneive_io_ibuf \my_rf.WEN~input (
	.i(\my_rf.WEN ),
	.ibar(gnd),
	.o(\my_rf.WEN~input_o ));
// synopsys translate_off
defparam \my_rf.WEN~input .bus_hold = "false";
defparam \my_rf.WEN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X42_Y31_N12
cycloneive_lcell_comb \Decoder0~14 (
// Equation(s):
// \Decoder0~14_combout  = (!\my_rf.wsel[0]~input_o  & (\my_rf.wsel[3]~input_o  & (!\my_rf.wsel[1]~input_o  & !\my_rf.wsel[2]~input_o )))

	.dataa(\my_rf.wsel[0]~input_o ),
	.datab(\my_rf.wsel[3]~input_o ),
	.datac(\my_rf.wsel[1]~input_o ),
	.datad(\my_rf.wsel[2]~input_o ),
	.cin(gnd),
	.combout(\Decoder0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~14 .lut_mask = 16'h0004;
defparam \Decoder0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y31_N24
cycloneive_lcell_comb \Decoder0~26 (
// Equation(s):
// \Decoder0~26_combout  = (!\my_rf.wsel[4]~input_o  & (\my_rf.WEN~input_o  & \Decoder0~14_combout ))

	.dataa(\my_rf.wsel[4]~input_o ),
	.datab(gnd),
	.datac(\my_rf.WEN~input_o ),
	.datad(\Decoder0~14_combout ),
	.cin(gnd),
	.combout(\Decoder0~26_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~26 .lut_mask = 16'h5000;
defparam \Decoder0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y31_N11
dffeas \registerArray[8][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][0] .is_wysiwyg = "true";
defparam \registerArray[8][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N0
cycloneive_lcell_comb \Mux63~10 (
// Equation(s):
// \Mux63~10_combout  = (\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o ) # ((\registerArray[10][0]~q )))) # (!\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & ((\registerArray[8][0]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[10][0]~q ),
	.datad(\registerArray[8][0]~q ),
	.cin(gnd),
	.combout(\Mux63~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~10 .lut_mask = 16'hB9A8;
defparam \Mux63~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y31_N8
cycloneive_lcell_comb \Decoder0~0 (
// Equation(s):
// \Decoder0~0_combout  = (\my_rf.wsel[0]~input_o  & (\my_rf.WEN~input_o  & (!\my_rf.wsel[1]~input_o  & !\my_rf.wsel[2]~input_o )))

	.dataa(\my_rf.wsel[0]~input_o ),
	.datab(\my_rf.WEN~input_o ),
	.datac(\my_rf.wsel[1]~input_o ),
	.datad(\my_rf.wsel[2]~input_o ),
	.cin(gnd),
	.combout(\Decoder0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~0 .lut_mask = 16'h0008;
defparam \Decoder0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y31_N24
cycloneive_lcell_comb \Decoder0~24 (
// Equation(s):
// \Decoder0~24_combout  = (\my_rf.wsel[3]~input_o  & (!\my_rf.wsel[4]~input_o  & \Decoder0~0_combout ))

	.dataa(\my_rf.wsel[3]~input_o ),
	.datab(gnd),
	.datac(\my_rf.wsel[4]~input_o ),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~24_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~24 .lut_mask = 16'h0A00;
defparam \Decoder0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y31_N1
dffeas \registerArray[9][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][0] .is_wysiwyg = "true";
defparam \registerArray[9][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N0
cycloneive_lcell_comb \Mux63~11 (
// Equation(s):
// \Mux63~11_combout  = (\Mux63~10_combout  & ((\registerArray[11][0]~q ) # ((!\my_rf.rsel2[0]~input_o )))) # (!\Mux63~10_combout  & (((\registerArray[9][0]~q  & \my_rf.rsel2[0]~input_o ))))

	.dataa(\registerArray[11][0]~q ),
	.datab(\Mux63~10_combout ),
	.datac(\registerArray[9][0]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux63~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~11 .lut_mask = 16'hB8CC;
defparam \Mux63~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X0_Y29_N15
cycloneive_io_ibuf \my_rf.rsel2[1]~input (
	.i(\my_rf.rsel2 [1]),
	.ibar(gnd),
	.o(\my_rf.rsel2[1]~input_o ));
// synopsys translate_off
defparam \my_rf.rsel2[1]~input .bus_hold = "false";
defparam \my_rf.rsel2[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X41_Y32_N22
cycloneive_lcell_comb \Decoder0~35 (
// Equation(s):
// \Decoder0~35_combout  = (\Decoder0~8_combout  & (\my_rf.wsel[2]~input_o  & !\my_rf.wsel[4]~input_o ))

	.dataa(gnd),
	.datab(\Decoder0~8_combout ),
	.datac(\my_rf.wsel[2]~input_o ),
	.datad(\my_rf.wsel[4]~input_o ),
	.cin(gnd),
	.combout(\Decoder0~35_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~35 .lut_mask = 16'h00C0;
defparam \Decoder0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N9
dffeas \registerArray[14][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][0] .is_wysiwyg = "true";
defparam \registerArray[14][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y31_N16
cycloneive_lcell_comb \Decoder0~12 (
// Equation(s):
// \Decoder0~12_combout  = (\my_rf.WEN~input_o  & (!\my_rf.wsel[1]~input_o  & \my_rf.wsel[2]~input_o ))

	.dataa(gnd),
	.datab(\my_rf.WEN~input_o ),
	.datac(\my_rf.wsel[1]~input_o ),
	.datad(\my_rf.wsel[2]~input_o ),
	.cin(gnd),
	.combout(\Decoder0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~12 .lut_mask = 16'h0C00;
defparam \Decoder0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y31_N20
cycloneive_lcell_comb \Decoder0~37 (
// Equation(s):
// \Decoder0~37_combout  = (!\my_rf.wsel[4]~input_o  & (\my_rf.wsel[3]~input_o  & (!\my_rf.wsel[0]~input_o  & \Decoder0~12_combout )))

	.dataa(\my_rf.wsel[4]~input_o ),
	.datab(\my_rf.wsel[3]~input_o ),
	.datac(\my_rf.wsel[0]~input_o ),
	.datad(\Decoder0~12_combout ),
	.cin(gnd),
	.combout(\Decoder0~37_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~37 .lut_mask = 16'h0400;
defparam \Decoder0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N3
dffeas \registerArray[12][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][0] .is_wysiwyg = "true";
defparam \registerArray[12][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y31_N2
cycloneive_lcell_comb \Decoder0~2 (
// Equation(s):
// \Decoder0~2_combout  = (\my_rf.wsel[0]~input_o  & (\my_rf.WEN~input_o  & (!\my_rf.wsel[1]~input_o  & \my_rf.wsel[2]~input_o )))

	.dataa(\my_rf.wsel[0]~input_o ),
	.datab(\my_rf.WEN~input_o ),
	.datac(\my_rf.wsel[1]~input_o ),
	.datad(\my_rf.wsel[2]~input_o ),
	.cin(gnd),
	.combout(\Decoder0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~2 .lut_mask = 16'h0800;
defparam \Decoder0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y31_N20
cycloneive_lcell_comb \Decoder0~36 (
// Equation(s):
// \Decoder0~36_combout  = (\my_rf.wsel[3]~input_o  & (!\my_rf.wsel[4]~input_o  & \Decoder0~2_combout ))

	.dataa(\my_rf.wsel[3]~input_o ),
	.datab(gnd),
	.datac(\my_rf.wsel[4]~input_o ),
	.datad(\Decoder0~2_combout ),
	.cin(gnd),
	.combout(\Decoder0~36_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~36 .lut_mask = 16'h0A00;
defparam \Decoder0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N25
dffeas \registerArray[13][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][0] .is_wysiwyg = "true";
defparam \registerArray[13][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N24
cycloneive_lcell_comb \Mux63~17 (
// Equation(s):
// \Mux63~17_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & ((\registerArray[13][0]~q ))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[12][0]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[12][0]~q ),
	.datac(\registerArray[13][0]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux63~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~17 .lut_mask = 16'hFA44;
defparam \Mux63~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N8
cycloneive_lcell_comb \Mux63~18 (
// Equation(s):
// \Mux63~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux63~17_combout  & (\registerArray[15][0]~q )) # (!\Mux63~17_combout  & ((\registerArray[14][0]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux63~17_combout ))))

	.dataa(\registerArray[15][0]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][0]~q ),
	.datad(\Mux63~17_combout ),
	.cin(gnd),
	.combout(\Mux63~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~18 .lut_mask = 16'hBBC0;
defparam \Mux63~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N4
cycloneive_lcell_comb \Mux63~19 (
// Equation(s):
// \Mux63~19_combout  = (\Mux63~16_combout  & (((\Mux63~18_combout )) # (!\my_rf.rsel2[3]~input_o ))) # (!\Mux63~16_combout  & (\my_rf.rsel2[3]~input_o  & (\Mux63~11_combout )))

	.dataa(\Mux63~16_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux63~11_combout ),
	.datad(\Mux63~18_combout ),
	.cin(gnd),
	.combout(\Mux63~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~19 .lut_mask = 16'hEA62;
defparam \Mux63~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N15
cycloneive_io_ibuf \my_rf.rsel2[2]~input (
	.i(\my_rf.rsel2 [2]),
	.ibar(gnd),
	.o(\my_rf.rsel2[2]~input_o ));
// synopsys translate_off
defparam \my_rf.rsel2[2]~input .bus_hold = "false";
defparam \my_rf.rsel2[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X42_Y31_N4
cycloneive_lcell_comb \Decoder0~6 (
// Equation(s):
// \Decoder0~6_combout  = (\my_rf.WEN~input_o  & (!\my_rf.wsel[3]~input_o  & (\my_rf.wsel[1]~input_o  & !\my_rf.wsel[0]~input_o )))

	.dataa(\my_rf.WEN~input_o ),
	.datab(\my_rf.wsel[3]~input_o ),
	.datac(\my_rf.wsel[1]~input_o ),
	.datad(\my_rf.wsel[0]~input_o ),
	.cin(gnd),
	.combout(\Decoder0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~6 .lut_mask = 16'h0020;
defparam \Decoder0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y32_N24
cycloneive_lcell_comb \Decoder0~7 (
// Equation(s):
// \Decoder0~7_combout  = (\my_rf.wsel[4]~input_o  & (\my_rf.wsel[2]~input_o  & \Decoder0~6_combout ))

	.dataa(gnd),
	.datab(\my_rf.wsel[4]~input_o ),
	.datac(\my_rf.wsel[2]~input_o ),
	.datad(\Decoder0~6_combout ),
	.cin(gnd),
	.combout(\Decoder0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~7 .lut_mask = 16'hC000;
defparam \Decoder0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N1
dffeas \registerArray[22][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][0] .is_wysiwyg = "true";
defparam \registerArray[22][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y32_N30
cycloneive_lcell_comb \Decoder0~11 (
// Equation(s):
// \Decoder0~11_combout  = (\Decoder0~8_combout  & (\my_rf.wsel[2]~input_o  & \my_rf.wsel[4]~input_o ))

	.dataa(gnd),
	.datab(\Decoder0~8_combout ),
	.datac(\my_rf.wsel[2]~input_o ),
	.datad(\my_rf.wsel[4]~input_o ),
	.cin(gnd),
	.combout(\Decoder0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~11 .lut_mask = 16'hC000;
defparam \Decoder0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y38_N17
dffeas \registerArray[30][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][0] .is_wysiwyg = "true";
defparam \registerArray[30][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N0
cycloneive_lcell_comb \Mux63~3 (
// Equation(s):
// \Mux63~3_combout  = (\Mux63~2_combout  & (((\registerArray[30][0]~q )) # (!\my_rf.rsel2[2]~input_o ))) # (!\Mux63~2_combout  & (\my_rf.rsel2[2]~input_o  & (\registerArray[22][0]~q )))

	.dataa(\Mux63~2_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][0]~q ),
	.datad(\registerArray[30][0]~q ),
	.cin(gnd),
	.combout(\Mux63~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~3 .lut_mask = 16'hEA62;
defparam \Mux63~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y31_N18
cycloneive_lcell_comb \Decoder0~13 (
// Equation(s):
// \Decoder0~13_combout  = (\my_rf.wsel[4]~input_o  & (!\my_rf.wsel[3]~input_o  & (!\my_rf.wsel[0]~input_o  & \Decoder0~12_combout )))

	.dataa(\my_rf.wsel[4]~input_o ),
	.datab(\my_rf.wsel[3]~input_o ),
	.datac(\my_rf.wsel[0]~input_o ),
	.datad(\Decoder0~12_combout ),
	.cin(gnd),
	.combout(\Decoder0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~13 .lut_mask = 16'h0200;
defparam \Decoder0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y35_N9
dffeas \registerArray[20][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][0] .is_wysiwyg = "true";
defparam \registerArray[20][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y31_N28
cycloneive_lcell_comb \Decoder0~18 (
// Equation(s):
// \Decoder0~18_combout  = (\my_rf.wsel[4]~input_o  & (\my_rf.wsel[3]~input_o  & (!\my_rf.wsel[0]~input_o  & \Decoder0~12_combout )))

	.dataa(\my_rf.wsel[4]~input_o ),
	.datab(\my_rf.wsel[3]~input_o ),
	.datac(\my_rf.wsel[0]~input_o ),
	.datad(\Decoder0~12_combout ),
	.cin(gnd),
	.combout(\Decoder0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~18 .lut_mask = 16'h0800;
defparam \Decoder0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y35_N9
dffeas \registerArray[28][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][0] .is_wysiwyg = "true";
defparam \registerArray[28][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N8
cycloneive_lcell_comb \Mux63~5 (
// Equation(s):
// \Mux63~5_combout  = (\Mux63~4_combout  & (((\registerArray[28][0]~q )) # (!\my_rf.rsel2[2]~input_o ))) # (!\Mux63~4_combout  & (\my_rf.rsel2[2]~input_o  & (\registerArray[20][0]~q )))

	.dataa(\Mux63~4_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[20][0]~q ),
	.datad(\registerArray[28][0]~q ),
	.cin(gnd),
	.combout(\Mux63~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~5 .lut_mask = 16'hEA62;
defparam \Mux63~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N14
cycloneive_lcell_comb \Mux63~6 (
// Equation(s):
// \Mux63~6_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux63~3_combout ) # ((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (((!\my_rf.rsel2[0]~input_o  & \Mux63~5_combout ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux63~3_combout ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux63~5_combout ),
	.cin(gnd),
	.combout(\Mux63~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~6 .lut_mask = 16'hADA8;
defparam \Mux63~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y31_N14
cycloneive_lcell_comb \Decoder0~5 (
// Equation(s):
// \Decoder0~5_combout  = (\my_rf.wsel[3]~input_o  & (\my_rf.wsel[4]~input_o  & \Decoder0~2_combout ))

	.dataa(\my_rf.wsel[3]~input_o ),
	.datab(gnd),
	.datac(\my_rf.wsel[4]~input_o ),
	.datad(\Decoder0~2_combout ),
	.cin(gnd),
	.combout(\Decoder0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~5 .lut_mask = 16'hA000;
defparam \Decoder0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y32_N25
dffeas \registerArray[29][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][0] .is_wysiwyg = "true";
defparam \registerArray[29][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y31_N2
cycloneive_lcell_comb \Decoder0~3 (
// Equation(s):
// \Decoder0~3_combout  = (!\my_rf.wsel[3]~input_o  & (\my_rf.wsel[4]~input_o  & \Decoder0~2_combout ))

	.dataa(\my_rf.wsel[3]~input_o ),
	.datab(gnd),
	.datac(\my_rf.wsel[4]~input_o ),
	.datad(\Decoder0~2_combout ),
	.cin(gnd),
	.combout(\Decoder0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~3 .lut_mask = 16'h5000;
defparam \Decoder0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N1
dffeas \registerArray[21][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][0] .is_wysiwyg = "true";
defparam \registerArray[21][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y31_N28
cycloneive_lcell_comb \Decoder0~4 (
// Equation(s):
// \Decoder0~4_combout  = (!\my_rf.wsel[3]~input_o  & (\my_rf.wsel[4]~input_o  & \Decoder0~0_combout ))

	.dataa(\my_rf.wsel[3]~input_o ),
	.datab(gnd),
	.datac(\my_rf.wsel[4]~input_o ),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~4 .lut_mask = 16'h5000;
defparam \Decoder0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N3
dffeas \registerArray[17][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][0] .is_wysiwyg = "true";
defparam \registerArray[17][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N0
cycloneive_lcell_comb \Mux63~0 (
// Equation(s):
// \Mux63~0_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[21][0]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[17][0]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[21][0]~q ),
	.datad(\registerArray[17][0]~q ),
	.cin(gnd),
	.combout(\Mux63~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~0 .lut_mask = 16'hB9A8;
defparam \Mux63~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N20
cycloneive_lcell_comb \Mux63~1 (
// Equation(s):
// \Mux63~1_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux63~0_combout  & ((\registerArray[29][0]~q ))) # (!\Mux63~0_combout  & (\registerArray[25][0]~q )))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux63~0_combout ))))

	.dataa(\registerArray[25][0]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[29][0]~q ),
	.datad(\Mux63~0_combout ),
	.cin(gnd),
	.combout(\Mux63~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~1 .lut_mask = 16'hF388;
defparam \Mux63~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N16
cycloneive_lcell_comb \Mux63~9 (
// Equation(s):
// \Mux63~9_combout  = (\Mux63~6_combout  & ((\Mux63~8_combout ) # ((!\my_rf.rsel2[0]~input_o )))) # (!\Mux63~6_combout  & (((\my_rf.rsel2[0]~input_o  & \Mux63~1_combout ))))

	.dataa(\Mux63~8_combout ),
	.datab(\Mux63~6_combout ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux63~1_combout ),
	.cin(gnd),
	.combout(\Mux63~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~9 .lut_mask = 16'hBC8C;
defparam \Mux63~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N22
cycloneive_lcell_comb \Mux63~20 (
// Equation(s):
// \Mux63~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux63~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux63~19_combout ))

	.dataa(gnd),
	.datab(\my_rf.rsel2[4]~input_o ),
	.datac(\Mux63~19_combout ),
	.datad(\Mux63~9_combout ),
	.cin(gnd),
	.combout(\Mux63~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~20 .lut_mask = 16'hFC30;
defparam \Mux63~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N22
cycloneive_io_ibuf \my_rf.wdat[1]~input (
	.i(\my_rf.wdat [1]),
	.ibar(gnd),
	.o(\my_rf.wdat[1]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[1]~input .bus_hold = "false";
defparam \my_rf.wdat[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X53_Y33_N13
dffeas \registerArray[14][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][1] .is_wysiwyg = "true";
defparam \registerArray[14][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N29
dffeas \registerArray[13][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][1] .is_wysiwyg = "true";
defparam \registerArray[13][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N28
cycloneive_lcell_comb \Mux62~17 (
// Equation(s):
// \Mux62~17_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & ((\registerArray[13][1]~q ))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[12][1]~q ))))

	.dataa(\registerArray[12][1]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[13][1]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux62~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~17 .lut_mask = 16'hFC22;
defparam \Mux62~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N12
cycloneive_lcell_comb \Mux62~18 (
// Equation(s):
// \Mux62~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux62~17_combout  & (\registerArray[15][1]~q )) # (!\Mux62~17_combout  & ((\registerArray[14][1]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux62~17_combout ))))

	.dataa(\registerArray[15][1]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][1]~q ),
	.datad(\Mux62~17_combout ),
	.cin(gnd),
	.combout(\Mux62~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~18 .lut_mask = 16'hBBC0;
defparam \Mux62~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y32_N26
cycloneive_lcell_comb \Decoder0~28 (
// Equation(s):
// \Decoder0~28_combout  = (!\my_rf.wsel[4]~input_o  & (\my_rf.wsel[2]~input_o  & \Decoder0~6_combout ))

	.dataa(gnd),
	.datab(\my_rf.wsel[4]~input_o ),
	.datac(\my_rf.wsel[2]~input_o ),
	.datad(\Decoder0~6_combout ),
	.cin(gnd),
	.combout(\Decoder0~28_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~28 .lut_mask = 16'h3000;
defparam \Decoder0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y29_N13
dffeas \registerArray[6][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][1] .is_wysiwyg = "true";
defparam \registerArray[6][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y31_N4
cycloneive_lcell_comb \Decoder0~29 (
// Equation(s):
// \Decoder0~29_combout  = (!\my_rf.wsel[3]~input_o  & (!\my_rf.wsel[4]~input_o  & \Decoder0~2_combout ))

	.dataa(\my_rf.wsel[3]~input_o ),
	.datab(gnd),
	.datac(\my_rf.wsel[4]~input_o ),
	.datad(\Decoder0~2_combout ),
	.cin(gnd),
	.combout(\Decoder0~29_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~29 .lut_mask = 16'h0500;
defparam \Decoder0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y29_N21
dffeas \registerArray[5][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][1] .is_wysiwyg = "true";
defparam \registerArray[5][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N20
cycloneive_lcell_comb \Mux62~10 (
// Equation(s):
// \Mux62~10_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[5][1]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][1]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[4][1]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][1]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux62~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~10 .lut_mask = 16'hCCE2;
defparam \Mux62~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N12
cycloneive_lcell_comb \Mux62~11 (
// Equation(s):
// \Mux62~11_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux62~10_combout  & (\registerArray[7][1]~q )) # (!\Mux62~10_combout  & ((\registerArray[6][1]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux62~10_combout ))))

	.dataa(\registerArray[7][1]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[6][1]~q ),
	.datad(\Mux62~10_combout ),
	.cin(gnd),
	.combout(\Mux62~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~11 .lut_mask = 16'hBBC0;
defparam \Mux62~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N6
cycloneive_lcell_comb \Mux62~19 (
// Equation(s):
// \Mux62~19_combout  = (\Mux62~16_combout  & ((\Mux62~18_combout ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux62~16_combout  & (((\my_rf.rsel2[2]~input_o  & \Mux62~11_combout ))))

	.dataa(\Mux62~16_combout ),
	.datab(\Mux62~18_combout ),
	.datac(\my_rf.rsel2[2]~input_o ),
	.datad(\Mux62~11_combout ),
	.cin(gnd),
	.combout(\Mux62~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~19 .lut_mask = 16'hDA8A;
defparam \Mux62~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y31_N14
cycloneive_lcell_comb \Decoder0~19 (
// Equation(s):
// \Decoder0~19_combout  = (\my_rf.WEN~input_o  & (\my_rf.wsel[1]~input_o  & \my_rf.wsel[0]~input_o ))

	.dataa(gnd),
	.datab(\my_rf.WEN~input_o ),
	.datac(\my_rf.wsel[1]~input_o ),
	.datad(\my_rf.wsel[0]~input_o ),
	.cin(gnd),
	.combout(\Decoder0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~19 .lut_mask = 16'hC000;
defparam \Decoder0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y31_N10
cycloneive_lcell_comb \Decoder0~21 (
// Equation(s):
// \Decoder0~21_combout  = (!\my_rf.wsel[3]~input_o  & (\my_rf.wsel[2]~input_o  & (\my_rf.wsel[4]~input_o  & \Decoder0~19_combout )))

	.dataa(\my_rf.wsel[3]~input_o ),
	.datab(\my_rf.wsel[2]~input_o ),
	.datac(\my_rf.wsel[4]~input_o ),
	.datad(\Decoder0~19_combout ),
	.cin(gnd),
	.combout(\Decoder0~21_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~21 .lut_mask = 16'h4000;
defparam \Decoder0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y28_N21
dffeas \registerArray[23][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][1] .is_wysiwyg = "true";
defparam \registerArray[23][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y31_N22
cycloneive_lcell_comb \Decoder0~23 (
// Equation(s):
// \Decoder0~23_combout  = (\my_rf.wsel[3]~input_o  & (\my_rf.wsel[2]~input_o  & (\my_rf.wsel[4]~input_o  & \Decoder0~19_combout )))

	.dataa(\my_rf.wsel[3]~input_o ),
	.datab(\my_rf.wsel[2]~input_o ),
	.datac(\my_rf.wsel[4]~input_o ),
	.datad(\Decoder0~19_combout ),
	.cin(gnd),
	.combout(\Decoder0~23_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~23 .lut_mask = 16'h8000;
defparam \Decoder0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y28_N31
dffeas \registerArray[31][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][1] .is_wysiwyg = "true";
defparam \registerArray[31][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N20
cycloneive_lcell_comb \Mux62~8 (
// Equation(s):
// \Mux62~8_combout  = (\Mux62~7_combout  & (((\registerArray[31][1]~q )) # (!\my_rf.rsel2[2]~input_o ))) # (!\Mux62~7_combout  & (\my_rf.rsel2[2]~input_o  & (\registerArray[23][1]~q )))

	.dataa(\Mux62~7_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[23][1]~q ),
	.datad(\registerArray[31][1]~q ),
	.cin(gnd),
	.combout(\Mux62~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~8 .lut_mask = 16'hEA62;
defparam \Mux62~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y36_N1
dffeas \registerArray[20][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][1] .is_wysiwyg = "true";
defparam \registerArray[20][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y31_N0
cycloneive_lcell_comb \Decoder0~16 (
// Equation(s):
// \Decoder0~16_combout  = (\my_rf.wsel[4]~input_o  & (\my_rf.WEN~input_o  & (!\my_rf.wsel[1]~input_o  & !\my_rf.wsel[2]~input_o )))

	.dataa(\my_rf.wsel[4]~input_o ),
	.datab(\my_rf.WEN~input_o ),
	.datac(\my_rf.wsel[1]~input_o ),
	.datad(\my_rf.wsel[2]~input_o ),
	.cin(gnd),
	.combout(\Decoder0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~16 .lut_mask = 16'h0008;
defparam \Decoder0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y31_N26
cycloneive_lcell_comb \Decoder0~17 (
// Equation(s):
// \Decoder0~17_combout  = (!\my_rf.wsel[0]~input_o  & (!\my_rf.wsel[3]~input_o  & \Decoder0~16_combout ))

	.dataa(\my_rf.wsel[0]~input_o ),
	.datab(\my_rf.wsel[3]~input_o ),
	.datac(gnd),
	.datad(\Decoder0~16_combout ),
	.cin(gnd),
	.combout(\Decoder0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~17 .lut_mask = 16'h1100;
defparam \Decoder0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y36_N3
dffeas \registerArray[16][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][1] .is_wysiwyg = "true";
defparam \registerArray[16][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N0
cycloneive_lcell_comb \Mux62~4 (
// Equation(s):
// \Mux62~4_combout  = (\my_rf.rsel2[3]~input_o  & (\my_rf.rsel2[2]~input_o )) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\registerArray[20][1]~q )) # (!\my_rf.rsel2[2]~input_o  & ((\registerArray[16][1]~q )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[20][1]~q ),
	.datad(\registerArray[16][1]~q ),
	.cin(gnd),
	.combout(\Mux62~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~4 .lut_mask = 16'hD9C8;
defparam \Mux62~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y31_N22
cycloneive_lcell_comb \Decoder0~15 (
// Equation(s):
// \Decoder0~15_combout  = (\my_rf.wsel[4]~input_o  & (\my_rf.WEN~input_o  & \Decoder0~14_combout ))

	.dataa(\my_rf.wsel[4]~input_o ),
	.datab(gnd),
	.datac(\my_rf.WEN~input_o ),
	.datad(\Decoder0~14_combout ),
	.cin(gnd),
	.combout(\Decoder0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~15 .lut_mask = 16'hA000;
defparam \Decoder0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N17
dffeas \registerArray[24][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][1] .is_wysiwyg = "true";
defparam \registerArray[24][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N19
dffeas \registerArray[28][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][1] .is_wysiwyg = "true";
defparam \registerArray[28][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N16
cycloneive_lcell_comb \Mux62~5 (
// Equation(s):
// \Mux62~5_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux62~4_combout  & ((\registerArray[28][1]~q ))) # (!\Mux62~4_combout  & (\registerArray[24][1]~q )))) # (!\my_rf.rsel2[3]~input_o  & (\Mux62~4_combout ))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux62~4_combout ),
	.datac(\registerArray[24][1]~q ),
	.datad(\registerArray[28][1]~q ),
	.cin(gnd),
	.combout(\Mux62~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~5 .lut_mask = 16'hEC64;
defparam \Mux62~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y32_N18
cycloneive_lcell_comb \Decoder0~9 (
// Equation(s):
// \Decoder0~9_combout  = (\Decoder0~8_combout  & (!\my_rf.wsel[2]~input_o  & \my_rf.wsel[4]~input_o ))

	.dataa(gnd),
	.datab(\Decoder0~8_combout ),
	.datac(\my_rf.wsel[2]~input_o ),
	.datad(\my_rf.wsel[4]~input_o ),
	.cin(gnd),
	.combout(\Decoder0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~9 .lut_mask = 16'h0C00;
defparam \Decoder0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y32_N1
dffeas \registerArray[26][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][1] .is_wysiwyg = "true";
defparam \registerArray[26][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y36_N17
dffeas \registerArray[22][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][1] .is_wysiwyg = "true";
defparam \registerArray[22][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N16
cycloneive_lcell_comb \Mux62~2 (
// Equation(s):
// \Mux62~2_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[22][1]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[18][1]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[18][1]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][1]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux62~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~2 .lut_mask = 16'hCCE2;
defparam \Mux62~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N0
cycloneive_lcell_comb \Mux62~3 (
// Equation(s):
// \Mux62~3_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux62~2_combout  & (\registerArray[30][1]~q )) # (!\Mux62~2_combout  & ((\registerArray[26][1]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux62~2_combout ))))

	.dataa(\registerArray[30][1]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[26][1]~q ),
	.datad(\Mux62~2_combout ),
	.cin(gnd),
	.combout(\Mux62~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~3 .lut_mask = 16'hBBC0;
defparam \Mux62~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N24
cycloneive_lcell_comb \Mux62~6 (
// Equation(s):
// \Mux62~6_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o ) # (\Mux62~3_combout )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux62~5_combout  & (!\my_rf.rsel2[0]~input_o )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux62~5_combout ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux62~3_combout ),
	.cin(gnd),
	.combout(\Mux62~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~6 .lut_mask = 16'hAEA4;
defparam \Mux62~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N10
cycloneive_lcell_comb \Mux62~9 (
// Equation(s):
// \Mux62~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux62~6_combout  & ((\Mux62~8_combout ))) # (!\Mux62~6_combout  & (\Mux62~1_combout )))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux62~6_combout ))))

	.dataa(\Mux62~1_combout ),
	.datab(\Mux62~8_combout ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux62~6_combout ),
	.cin(gnd),
	.combout(\Mux62~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~9 .lut_mask = 16'hCFA0;
defparam \Mux62~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N8
cycloneive_lcell_comb \Mux62~20 (
// Equation(s):
// \Mux62~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux62~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux62~19_combout ))

	.dataa(\Mux62~19_combout ),
	.datab(gnd),
	.datac(\my_rf.rsel2[4]~input_o ),
	.datad(\Mux62~9_combout ),
	.cin(gnd),
	.combout(\Mux62~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~20 .lut_mask = 16'hFA0A;
defparam \Mux62~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N22
cycloneive_io_ibuf \my_rf.wdat[2]~input (
	.i(\my_rf.wdat [2]),
	.ibar(gnd),
	.o(\my_rf.wdat[2]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[2]~input .bus_hold = "false";
defparam \my_rf.wdat[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X53_Y33_N25
dffeas \registerArray[14][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][2] .is_wysiwyg = "true";
defparam \registerArray[14][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y31_N30
cycloneive_lcell_comb \Decoder0~38 (
// Equation(s):
// \Decoder0~38_combout  = (\my_rf.wsel[3]~input_o  & (\my_rf.wsel[2]~input_o  & (!\my_rf.wsel[4]~input_o  & \Decoder0~19_combout )))

	.dataa(\my_rf.wsel[3]~input_o ),
	.datab(\my_rf.wsel[2]~input_o ),
	.datac(\my_rf.wsel[4]~input_o ),
	.datad(\Decoder0~19_combout ),
	.cin(gnd),
	.combout(\Decoder0~38_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~38 .lut_mask = 16'h0800;
defparam \Decoder0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N19
dffeas \registerArray[15][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][2] .is_wysiwyg = "true";
defparam \registerArray[15][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N24
cycloneive_lcell_comb \Mux61~18 (
// Equation(s):
// \Mux61~18_combout  = (\Mux61~17_combout  & (((\registerArray[15][2]~q )) # (!\my_rf.rsel2[1]~input_o ))) # (!\Mux61~17_combout  & (\my_rf.rsel2[1]~input_o  & (\registerArray[14][2]~q )))

	.dataa(\Mux61~17_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][2]~q ),
	.datad(\registerArray[15][2]~q ),
	.cin(gnd),
	.combout(\Mux61~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~18 .lut_mask = 16'hEA62;
defparam \Mux61~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y29_N1
dffeas \registerArray[6][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][2] .is_wysiwyg = "true";
defparam \registerArray[6][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y29_N1
dffeas \registerArray[5][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][2] .is_wysiwyg = "true";
defparam \registerArray[5][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N0
cycloneive_lcell_comb \Mux61~12 (
// Equation(s):
// \Mux61~12_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[5][2]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][2]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[4][2]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][2]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux61~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~12 .lut_mask = 16'hCCE2;
defparam \Mux61~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N0
cycloneive_lcell_comb \Mux61~13 (
// Equation(s):
// \Mux61~13_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux61~12_combout  & (\registerArray[7][2]~q )) # (!\Mux61~12_combout  & ((\registerArray[6][2]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux61~12_combout ))))

	.dataa(\registerArray[7][2]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[6][2]~q ),
	.datad(\Mux61~12_combout ),
	.cin(gnd),
	.combout(\Mux61~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~13 .lut_mask = 16'hBBC0;
defparam \Mux61~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y32_N28
cycloneive_lcell_comb \Decoder0~34 (
// Equation(s):
// \Decoder0~34_combout  = (!\my_rf.wsel[4]~input_o  & (!\my_rf.wsel[2]~input_o  & \Decoder0~6_combout ))

	.dataa(gnd),
	.datab(\my_rf.wsel[4]~input_o ),
	.datac(\my_rf.wsel[2]~input_o ),
	.datad(\Decoder0~6_combout ),
	.cin(gnd),
	.combout(\Decoder0~34_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~34 .lut_mask = 16'h0300;
defparam \Decoder0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N27
dffeas \registerArray[2][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][2] .is_wysiwyg = "true";
defparam \registerArray[2][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y31_N8
cycloneive_lcell_comb \Decoder0~32 (
// Equation(s):
// \Decoder0~32_combout  = (!\my_rf.wsel[3]~input_o  & (!\my_rf.wsel[2]~input_o  & (!\my_rf.wsel[4]~input_o  & \Decoder0~19_combout )))

	.dataa(\my_rf.wsel[3]~input_o ),
	.datab(\my_rf.wsel[2]~input_o ),
	.datac(\my_rf.wsel[4]~input_o ),
	.datad(\Decoder0~19_combout ),
	.cin(gnd),
	.combout(\Decoder0~32_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~32 .lut_mask = 16'h0100;
defparam \Decoder0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y31_N25
dffeas \registerArray[3][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][2] .is_wysiwyg = "true";
defparam \registerArray[3][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N24
cycloneive_lcell_comb \Mux61~14 (
// Equation(s):
// \Mux61~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[3][2]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[1][2]~q ))))

	.dataa(\registerArray[1][2]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][2]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux61~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~14 .lut_mask = 16'hC088;
defparam \Mux61~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N26
cycloneive_lcell_comb \Mux61~15 (
// Equation(s):
// \Mux61~15_combout  = (\Mux61~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][2]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][2]~q ),
	.datad(\Mux61~14_combout ),
	.cin(gnd),
	.combout(\Mux61~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~15 .lut_mask = 16'hFF20;
defparam \Mux61~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N6
cycloneive_lcell_comb \Mux61~16 (
// Equation(s):
// \Mux61~16_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\Mux61~13_combout )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\Mux61~15_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux61~13_combout ),
	.datad(\Mux61~15_combout ),
	.cin(gnd),
	.combout(\Mux61~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~16 .lut_mask = 16'hB9A8;
defparam \Mux61~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N8
cycloneive_lcell_comb \Mux61~19 (
// Equation(s):
// \Mux61~19_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux61~16_combout  & ((\Mux61~18_combout ))) # (!\Mux61~16_combout  & (\Mux61~11_combout )))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux61~16_combout ))))

	.dataa(\Mux61~11_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux61~18_combout ),
	.datad(\Mux61~16_combout ),
	.cin(gnd),
	.combout(\Mux61~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~19 .lut_mask = 16'hF388;
defparam \Mux61~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y28_N19
dffeas \registerArray[31][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][2] .is_wysiwyg = "true";
defparam \registerArray[31][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y31_N16
cycloneive_lcell_comb \Decoder0~20 (
// Equation(s):
// \Decoder0~20_combout  = (\my_rf.wsel[3]~input_o  & (!\my_rf.wsel[2]~input_o  & (\my_rf.wsel[4]~input_o  & \Decoder0~19_combout )))

	.dataa(\my_rf.wsel[3]~input_o ),
	.datab(\my_rf.wsel[2]~input_o ),
	.datac(\my_rf.wsel[4]~input_o ),
	.datad(\Decoder0~19_combout ),
	.cin(gnd),
	.combout(\Decoder0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~20 .lut_mask = 16'h2000;
defparam \Decoder0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y28_N9
dffeas \registerArray[27][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][2] .is_wysiwyg = "true";
defparam \registerArray[27][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N25
dffeas \registerArray[23][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][2] .is_wysiwyg = "true";
defparam \registerArray[23][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y31_N12
cycloneive_lcell_comb \Decoder0~22 (
// Equation(s):
// \Decoder0~22_combout  = (!\my_rf.wsel[3]~input_o  & (!\my_rf.wsel[2]~input_o  & (\my_rf.wsel[4]~input_o  & \Decoder0~19_combout )))

	.dataa(\my_rf.wsel[3]~input_o ),
	.datab(\my_rf.wsel[2]~input_o ),
	.datac(\my_rf.wsel[4]~input_o ),
	.datad(\Decoder0~19_combout ),
	.cin(gnd),
	.combout(\Decoder0~22_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~22 .lut_mask = 16'h1000;
defparam \Decoder0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y28_N19
dffeas \registerArray[19][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][2] .is_wysiwyg = "true";
defparam \registerArray[19][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N24
cycloneive_lcell_comb \Mux61~7 (
// Equation(s):
// \Mux61~7_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[23][2]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[19][2]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[23][2]~q ),
	.datad(\registerArray[19][2]~q ),
	.cin(gnd),
	.combout(\Mux61~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~7 .lut_mask = 16'hB9A8;
defparam \Mux61~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N8
cycloneive_lcell_comb \Mux61~8 (
// Equation(s):
// \Mux61~8_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux61~7_combout  & (\registerArray[31][2]~q )) # (!\Mux61~7_combout  & ((\registerArray[27][2]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux61~7_combout ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[31][2]~q ),
	.datac(\registerArray[27][2]~q ),
	.datad(\Mux61~7_combout ),
	.cin(gnd),
	.combout(\Mux61~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~8 .lut_mask = 16'hDDA0;
defparam \Mux61~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N27
dffeas \registerArray[29][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][2] .is_wysiwyg = "true";
defparam \registerArray[29][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N19
dffeas \registerArray[21][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][2] .is_wysiwyg = "true";
defparam \registerArray[21][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N29
dffeas \registerArray[17][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][2] .is_wysiwyg = "true";
defparam \registerArray[17][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N18
cycloneive_lcell_comb \Mux61~0 (
// Equation(s):
// \Mux61~0_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[21][2]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[17][2]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[21][2]~q ),
	.datad(\registerArray[17][2]~q ),
	.cin(gnd),
	.combout(\Mux61~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~0 .lut_mask = 16'hB9A8;
defparam \Mux61~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N0
cycloneive_lcell_comb \Mux61~1 (
// Equation(s):
// \Mux61~1_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux61~0_combout  & ((\registerArray[29][2]~q ))) # (!\Mux61~0_combout  & (\registerArray[25][2]~q )))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux61~0_combout ))))

	.dataa(\registerArray[25][2]~q ),
	.datab(\registerArray[29][2]~q ),
	.datac(\my_rf.rsel2[3]~input_o ),
	.datad(\Mux61~0_combout ),
	.cin(gnd),
	.combout(\Mux61~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~1 .lut_mask = 16'hCFA0;
defparam \Mux61~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N12
cycloneive_lcell_comb \Mux61~9 (
// Equation(s):
// \Mux61~9_combout  = (\Mux61~6_combout  & (((\Mux61~8_combout )) # (!\my_rf.rsel2[0]~input_o ))) # (!\Mux61~6_combout  & (\my_rf.rsel2[0]~input_o  & ((\Mux61~1_combout ))))

	.dataa(\Mux61~6_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux61~8_combout ),
	.datad(\Mux61~1_combout ),
	.cin(gnd),
	.combout(\Mux61~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~9 .lut_mask = 16'hE6A2;
defparam \Mux61~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N18
cycloneive_lcell_comb \Mux61~20 (
// Equation(s):
// \Mux61~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux61~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux61~19_combout ))

	.dataa(gnd),
	.datab(\my_rf.rsel2[4]~input_o ),
	.datac(\Mux61~19_combout ),
	.datad(\Mux61~9_combout ),
	.cin(gnd),
	.combout(\Mux61~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~20 .lut_mask = 16'hFC30;
defparam \Mux61~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N15
cycloneive_io_ibuf \my_rf.wdat[3]~input (
	.i(\my_rf.wdat [3]),
	.ibar(gnd),
	.o(\my_rf.wdat[3]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[3]~input .bus_hold = "false";
defparam \my_rf.wdat[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X43_Y31_N6
cycloneive_lcell_comb \Decoder0~31 (
// Equation(s):
// \Decoder0~31_combout  = (!\my_rf.wsel[3]~input_o  & (\my_rf.wsel[2]~input_o  & (!\my_rf.wsel[4]~input_o  & \Decoder0~19_combout )))

	.dataa(\my_rf.wsel[3]~input_o ),
	.datab(\my_rf.wsel[2]~input_o ),
	.datac(\my_rf.wsel[4]~input_o ),
	.datad(\Decoder0~19_combout ),
	.cin(gnd),
	.combout(\Decoder0~31_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~31 .lut_mask = 16'h0400;
defparam \Decoder0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y29_N15
dffeas \registerArray[7][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][3] .is_wysiwyg = "true";
defparam \registerArray[7][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y29_N29
dffeas \registerArray[6][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][3] .is_wysiwyg = "true";
defparam \registerArray[6][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N28
cycloneive_lcell_comb \Mux60~11 (
// Equation(s):
// \Mux60~11_combout  = (\Mux60~10_combout  & ((\registerArray[7][3]~q ) # ((!\my_rf.rsel2[1]~input_o )))) # (!\Mux60~10_combout  & (((\registerArray[6][3]~q  & \my_rf.rsel2[1]~input_o ))))

	.dataa(\Mux60~10_combout ),
	.datab(\registerArray[7][3]~q ),
	.datac(\registerArray[6][3]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux60~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~11 .lut_mask = 16'hD8AA;
defparam \Mux60~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y31_N5
dffeas \registerArray[9][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][3] .is_wysiwyg = "true";
defparam \registerArray[9][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y31_N5
dffeas \registerArray[10][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][3] .is_wysiwyg = "true";
defparam \registerArray[10][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N4
cycloneive_lcell_comb \Mux60~12 (
// Equation(s):
// \Mux60~12_combout  = (\my_rf.rsel2[0]~input_o  & (((\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[10][3]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[8][3]~q ))))

	.dataa(\registerArray[8][3]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[10][3]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux60~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~12 .lut_mask = 16'hFC22;
defparam \Mux60~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N4
cycloneive_lcell_comb \Mux60~13 (
// Equation(s):
// \Mux60~13_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux60~12_combout  & (\registerArray[11][3]~q )) # (!\Mux60~12_combout  & ((\registerArray[9][3]~q ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux60~12_combout ))))

	.dataa(\registerArray[11][3]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[9][3]~q ),
	.datad(\Mux60~12_combout ),
	.cin(gnd),
	.combout(\Mux60~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~13 .lut_mask = 16'hBBC0;
defparam \Mux60~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N21
dffeas \registerArray[2][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][3] .is_wysiwyg = "true";
defparam \registerArray[2][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N13
dffeas \registerArray[3][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][3] .is_wysiwyg = "true";
defparam \registerArray[3][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N12
cycloneive_lcell_comb \Mux60~14 (
// Equation(s):
// \Mux60~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[3][3]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[1][3]~q ))))

	.dataa(\registerArray[1][3]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][3]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux60~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~14 .lut_mask = 16'hC088;
defparam \Mux60~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N20
cycloneive_lcell_comb \Mux60~15 (
// Equation(s):
// \Mux60~15_combout  = (\Mux60~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][3]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][3]~q ),
	.datad(\Mux60~14_combout ),
	.cin(gnd),
	.combout(\Mux60~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~15 .lut_mask = 16'hFF20;
defparam \Mux60~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N26
cycloneive_lcell_comb \Mux60~16 (
// Equation(s):
// \Mux60~16_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\Mux60~13_combout )) # (!\my_rf.rsel2[3]~input_o  & ((\Mux60~15_combout )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux60~13_combout ),
	.datac(\my_rf.rsel2[3]~input_o ),
	.datad(\Mux60~15_combout ),
	.cin(gnd),
	.combout(\Mux60~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~16 .lut_mask = 16'hE5E0;
defparam \Mux60~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N21
dffeas \registerArray[14][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][3] .is_wysiwyg = "true";
defparam \registerArray[14][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N15
dffeas \registerArray[12][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][3] .is_wysiwyg = "true";
defparam \registerArray[12][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N21
dffeas \registerArray[13][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][3] .is_wysiwyg = "true";
defparam \registerArray[13][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N20
cycloneive_lcell_comb \Mux60~17 (
// Equation(s):
// \Mux60~17_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & ((\registerArray[13][3]~q ))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[12][3]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[12][3]~q ),
	.datac(\registerArray[13][3]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux60~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~17 .lut_mask = 16'hFA44;
defparam \Mux60~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N20
cycloneive_lcell_comb \Mux60~18 (
// Equation(s):
// \Mux60~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux60~17_combout  & (\registerArray[15][3]~q )) # (!\Mux60~17_combout  & ((\registerArray[14][3]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux60~17_combout ))))

	.dataa(\registerArray[15][3]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][3]~q ),
	.datad(\Mux60~17_combout ),
	.cin(gnd),
	.combout(\Mux60~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~18 .lut_mask = 16'hBBC0;
defparam \Mux60~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N28
cycloneive_lcell_comb \Mux60~19 (
// Equation(s):
// \Mux60~19_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux60~16_combout  & ((\Mux60~18_combout ))) # (!\Mux60~16_combout  & (\Mux60~11_combout )))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux60~16_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux60~11_combout ),
	.datac(\Mux60~16_combout ),
	.datad(\Mux60~18_combout ),
	.cin(gnd),
	.combout(\Mux60~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~19 .lut_mask = 16'hF858;
defparam \Mux60~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N9
dffeas \registerArray[29][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][3] .is_wysiwyg = "true";
defparam \registerArray[29][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y0_N17
dffeas \registerArray[21][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[3]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][3] .is_wysiwyg = "true";
defparam \registerArray[21][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y31_N0
cycloneive_lcell_comb \Decoder0~1 (
// Equation(s):
// \Decoder0~1_combout  = (\my_rf.wsel[3]~input_o  & (\my_rf.wsel[4]~input_o  & \Decoder0~0_combout ))

	.dataa(\my_rf.wsel[3]~input_o ),
	.datab(gnd),
	.datac(\my_rf.wsel[4]~input_o ),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~1 .lut_mask = 16'hA000;
defparam \Decoder0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N5
dffeas \registerArray[25][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][3] .is_wysiwyg = "true";
defparam \registerArray[25][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N4
cycloneive_lcell_comb \Mux60~0 (
// Equation(s):
// \Mux60~0_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & ((\registerArray[25][3]~q ))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[17][3]~q ))))

	.dataa(\registerArray[17][3]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[25][3]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux60~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~0 .lut_mask = 16'hFC22;
defparam \Mux60~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N4
cycloneive_lcell_comb \Mux60~1 (
// Equation(s):
// \Mux60~1_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux60~0_combout  & (\registerArray[29][3]~q )) # (!\Mux60~0_combout  & ((\registerArray[21][3]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux60~0_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[29][3]~q ),
	.datac(\registerArray[21][3]~q ),
	.datad(\Mux60~0_combout ),
	.cin(gnd),
	.combout(\Mux60~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~1 .lut_mask = 16'hDDA0;
defparam \Mux60~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y28_N29
dffeas \registerArray[23][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][3] .is_wysiwyg = "true";
defparam \registerArray[23][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y28_N29
dffeas \registerArray[27][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][3] .is_wysiwyg = "true";
defparam \registerArray[27][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N31
dffeas \registerArray[19][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][3] .is_wysiwyg = "true";
defparam \registerArray[19][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N28
cycloneive_lcell_comb \Mux60~7 (
// Equation(s):
// \Mux60~7_combout  = (\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o ) # ((\registerArray[27][3]~q )))) # (!\my_rf.rsel2[3]~input_o  & (!\my_rf.rsel2[2]~input_o  & ((\registerArray[19][3]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[27][3]~q ),
	.datad(\registerArray[19][3]~q ),
	.cin(gnd),
	.combout(\Mux60~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~7 .lut_mask = 16'hB9A8;
defparam \Mux60~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N28
cycloneive_lcell_comb \Mux60~8 (
// Equation(s):
// \Mux60~8_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux60~7_combout  & (\registerArray[31][3]~q )) # (!\Mux60~7_combout  & ((\registerArray[23][3]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux60~7_combout ))))

	.dataa(\registerArray[31][3]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[23][3]~q ),
	.datad(\Mux60~7_combout ),
	.cin(gnd),
	.combout(\Mux60~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~8 .lut_mask = 16'hBBC0;
defparam \Mux60~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N16
cycloneive_lcell_comb \Mux60~9 (
// Equation(s):
// \Mux60~9_combout  = (\Mux60~6_combout  & (((\Mux60~8_combout )) # (!\my_rf.rsel2[0]~input_o ))) # (!\Mux60~6_combout  & (\my_rf.rsel2[0]~input_o  & (\Mux60~1_combout )))

	.dataa(\Mux60~6_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux60~1_combout ),
	.datad(\Mux60~8_combout ),
	.cin(gnd),
	.combout(\Mux60~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~9 .lut_mask = 16'hEA62;
defparam \Mux60~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N14
cycloneive_lcell_comb \Mux60~20 (
// Equation(s):
// \Mux60~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux60~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux60~19_combout ))

	.dataa(gnd),
	.datab(\Mux60~19_combout ),
	.datac(\my_rf.rsel2[4]~input_o ),
	.datad(\Mux60~9_combout ),
	.cin(gnd),
	.combout(\Mux60~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~20 .lut_mask = 16'hFC0C;
defparam \Mux60~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N22
cycloneive_io_ibuf \my_rf.wdat[4]~input (
	.i(\my_rf.wdat [4]),
	.ibar(gnd),
	.o(\my_rf.wdat[4]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[4]~input .bus_hold = "false";
defparam \my_rf.wdat[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X45_Y33_N1
dffeas \registerArray[21][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][4] .is_wysiwyg = "true";
defparam \registerArray[21][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N11
dffeas \registerArray[17][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][4] .is_wysiwyg = "true";
defparam \registerArray[17][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N0
cycloneive_lcell_comb \Mux59~0 (
// Equation(s):
// \Mux59~0_combout  = (\my_rf.rsel2[3]~input_o  & (\my_rf.rsel2[2]~input_o )) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\registerArray[21][4]~q )) # (!\my_rf.rsel2[2]~input_o  & ((\registerArray[17][4]~q )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[21][4]~q ),
	.datad(\registerArray[17][4]~q ),
	.cin(gnd),
	.combout(\Mux59~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~0 .lut_mask = 16'hD9C8;
defparam \Mux59~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y0_N24
dffeas \registerArray[25][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[4]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][4] .is_wysiwyg = "true";
defparam \registerArray[25][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N0
cycloneive_lcell_comb \Mux59~1 (
// Equation(s):
// \Mux59~1_combout  = (\Mux59~0_combout  & ((\registerArray[29][4]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux59~0_combout  & (((\my_rf.rsel2[3]~input_o  & \registerArray[25][4]~q ))))

	.dataa(\registerArray[29][4]~q ),
	.datab(\Mux59~0_combout ),
	.datac(\my_rf.rsel2[3]~input_o ),
	.datad(\registerArray[25][4]~q ),
	.cin(gnd),
	.combout(\Mux59~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~1 .lut_mask = 16'hBC8C;
defparam \Mux59~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y32_N25
dffeas \registerArray[27][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][4] .is_wysiwyg = "true";
defparam \registerArray[27][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y32_N19
dffeas \registerArray[31][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][4] .is_wysiwyg = "true";
defparam \registerArray[31][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N24
cycloneive_lcell_comb \Mux59~8 (
// Equation(s):
// \Mux59~8_combout  = (\Mux59~7_combout  & (((\registerArray[31][4]~q )) # (!\my_rf.rsel2[3]~input_o ))) # (!\Mux59~7_combout  & (\my_rf.rsel2[3]~input_o  & (\registerArray[27][4]~q )))

	.dataa(\Mux59~7_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][4]~q ),
	.datad(\registerArray[31][4]~q ),
	.cin(gnd),
	.combout(\Mux59~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~8 .lut_mask = 16'hEA62;
defparam \Mux59~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N27
dffeas \registerArray[28][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][4] .is_wysiwyg = "true";
defparam \registerArray[28][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N29
dffeas \registerArray[20][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][4] .is_wysiwyg = "true";
defparam \registerArray[20][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y31_N3
dffeas \registerArray[24][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][4] .is_wysiwyg = "true";
defparam \registerArray[24][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y31_N29
dffeas \registerArray[16][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][4] .is_wysiwyg = "true";
defparam \registerArray[16][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N2
cycloneive_lcell_comb \Mux59~4 (
// Equation(s):
// \Mux59~4_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[24][4]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][4]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][4]~q ),
	.datad(\registerArray[16][4]~q ),
	.cin(gnd),
	.combout(\Mux59~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~4 .lut_mask = 16'hD9C8;
defparam \Mux59~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N28
cycloneive_lcell_comb \Mux59~5 (
// Equation(s):
// \Mux59~5_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux59~4_combout  & (\registerArray[28][4]~q )) # (!\Mux59~4_combout  & ((\registerArray[20][4]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux59~4_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[28][4]~q ),
	.datac(\registerArray[20][4]~q ),
	.datad(\Mux59~4_combout ),
	.cin(gnd),
	.combout(\Mux59~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~5 .lut_mask = 16'hDDA0;
defparam \Mux59~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N6
cycloneive_lcell_comb \Mux59~6 (
// Equation(s):
// \Mux59~6_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux59~3_combout ) # ((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (((!\my_rf.rsel2[0]~input_o  & \Mux59~5_combout ))))

	.dataa(\Mux59~3_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux59~5_combout ),
	.cin(gnd),
	.combout(\Mux59~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~6 .lut_mask = 16'hCBC8;
defparam \Mux59~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N8
cycloneive_lcell_comb \Mux59~9 (
// Equation(s):
// \Mux59~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux59~6_combout  & ((\Mux59~8_combout ))) # (!\Mux59~6_combout  & (\Mux59~1_combout )))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux59~6_combout ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\Mux59~1_combout ),
	.datac(\Mux59~8_combout ),
	.datad(\Mux59~6_combout ),
	.cin(gnd),
	.combout(\Mux59~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~9 .lut_mask = 16'hF588;
defparam \Mux59~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y31_N9
dffeas \registerArray[10][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][4] .is_wysiwyg = "true";
defparam \registerArray[10][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N8
cycloneive_lcell_comb \Mux59~10 (
// Equation(s):
// \Mux59~10_combout  = (\my_rf.rsel2[0]~input_o  & (((\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[10][4]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[8][4]~q ))))

	.dataa(\registerArray[8][4]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[10][4]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux59~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~10 .lut_mask = 16'hFC22;
defparam \Mux59~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y31_N17
dffeas \registerArray[9][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][4] .is_wysiwyg = "true";
defparam \registerArray[9][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N16
cycloneive_lcell_comb \Mux59~11 (
// Equation(s):
// \Mux59~11_combout  = (\Mux59~10_combout  & ((\registerArray[11][4]~q ) # ((!\my_rf.rsel2[0]~input_o )))) # (!\Mux59~10_combout  & (((\registerArray[9][4]~q  & \my_rf.rsel2[0]~input_o ))))

	.dataa(\registerArray[11][4]~q ),
	.datab(\Mux59~10_combout ),
	.datac(\registerArray[9][4]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux59~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~11 .lut_mask = 16'hB8CC;
defparam \Mux59~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N19
dffeas \registerArray[12][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][4] .is_wysiwyg = "true";
defparam \registerArray[12][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N9
dffeas \registerArray[13][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][4] .is_wysiwyg = "true";
defparam \registerArray[13][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N8
cycloneive_lcell_comb \Mux59~17 (
// Equation(s):
// \Mux59~17_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & ((\registerArray[13][4]~q ))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[12][4]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[12][4]~q ),
	.datac(\registerArray[13][4]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux59~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~17 .lut_mask = 16'hFA44;
defparam \Mux59~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N17
dffeas \registerArray[14][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][4] .is_wysiwyg = "true";
defparam \registerArray[14][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N3
dffeas \registerArray[15][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][4] .is_wysiwyg = "true";
defparam \registerArray[15][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N16
cycloneive_lcell_comb \Mux59~18 (
// Equation(s):
// \Mux59~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux59~17_combout  & ((\registerArray[15][4]~q ))) # (!\Mux59~17_combout  & (\registerArray[14][4]~q )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux59~17_combout ))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux59~17_combout ),
	.datac(\registerArray[14][4]~q ),
	.datad(\registerArray[15][4]~q ),
	.cin(gnd),
	.combout(\Mux59~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~18 .lut_mask = 16'hEC64;
defparam \Mux59~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N20
cycloneive_lcell_comb \Mux59~19 (
// Equation(s):
// \Mux59~19_combout  = (\Mux59~16_combout  & (((\Mux59~18_combout ) # (!\my_rf.rsel2[3]~input_o )))) # (!\Mux59~16_combout  & (\Mux59~11_combout  & (\my_rf.rsel2[3]~input_o )))

	.dataa(\Mux59~16_combout ),
	.datab(\Mux59~11_combout ),
	.datac(\my_rf.rsel2[3]~input_o ),
	.datad(\Mux59~18_combout ),
	.cin(gnd),
	.combout(\Mux59~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~19 .lut_mask = 16'hEA4A;
defparam \Mux59~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N14
cycloneive_lcell_comb \Mux59~20 (
// Equation(s):
// \Mux59~20_combout  = (\my_rf.rsel2[4]~input_o  & (\Mux59~9_combout )) # (!\my_rf.rsel2[4]~input_o  & ((\Mux59~19_combout )))

	.dataa(gnd),
	.datab(\my_rf.rsel2[4]~input_o ),
	.datac(\Mux59~9_combout ),
	.datad(\Mux59~19_combout ),
	.cin(gnd),
	.combout(\Mux59~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~20 .lut_mask = 16'hF3C0;
defparam \Mux59~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N1
cycloneive_io_ibuf \my_rf.wdat[5]~input (
	.i(\my_rf.wdat [5]),
	.ibar(gnd),
	.o(\my_rf.wdat[5]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[5]~input .bus_hold = "false";
defparam \my_rf.wdat[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X53_Y35_N9
dffeas \registerArray[2][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][5] .is_wysiwyg = "true";
defparam \registerArray[2][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N8
cycloneive_lcell_comb \Mux58~15 (
// Equation(s):
// \Mux58~15_combout  = (\Mux58~14_combout ) # ((!\my_rf.rsel2[0]~input_o  & (\registerArray[2][5]~q  & \my_rf.rsel2[1]~input_o )))

	.dataa(\Mux58~14_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][5]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux58~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~15 .lut_mask = 16'hBAAA;
defparam \Mux58~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N18
cycloneive_lcell_comb \Mux58~16 (
// Equation(s):
// \Mux58~16_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux58~13_combout ) # ((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux58~15_combout  & !\my_rf.rsel2[2]~input_o ))))

	.dataa(\Mux58~13_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux58~15_combout ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux58~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~16 .lut_mask = 16'hCCB8;
defparam \Mux58~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N29
dffeas \registerArray[14][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][5] .is_wysiwyg = "true";
defparam \registerArray[14][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N1
dffeas \registerArray[12][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][5] .is_wysiwyg = "true";
defparam \registerArray[12][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N23
dffeas \registerArray[13][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][5] .is_wysiwyg = "true";
defparam \registerArray[13][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N22
cycloneive_lcell_comb \Mux58~17 (
// Equation(s):
// \Mux58~17_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & ((\registerArray[13][5]~q ))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[12][5]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[12][5]~q ),
	.datac(\registerArray[13][5]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux58~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~17 .lut_mask = 16'hFA44;
defparam \Mux58~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N28
cycloneive_lcell_comb \Mux58~18 (
// Equation(s):
// \Mux58~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux58~17_combout  & (\registerArray[15][5]~q )) # (!\Mux58~17_combout  & ((\registerArray[14][5]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux58~17_combout ))))

	.dataa(\registerArray[15][5]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][5]~q ),
	.datad(\Mux58~17_combout ),
	.cin(gnd),
	.combout(\Mux58~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~18 .lut_mask = 16'hBBC0;
defparam \Mux58~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N12
cycloneive_lcell_comb \Mux58~19 (
// Equation(s):
// \Mux58~19_combout  = (\Mux58~16_combout  & (((\Mux58~18_combout ) # (!\my_rf.rsel2[2]~input_o )))) # (!\Mux58~16_combout  & (\Mux58~11_combout  & ((\my_rf.rsel2[2]~input_o ))))

	.dataa(\Mux58~11_combout ),
	.datab(\Mux58~16_combout ),
	.datac(\Mux58~18_combout ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux58~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~19 .lut_mask = 16'hE2CC;
defparam \Mux58~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N9
dffeas \registerArray[25][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][5] .is_wysiwyg = "true";
defparam \registerArray[25][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N8
cycloneive_lcell_comb \Mux58~0 (
// Equation(s):
// \Mux58~0_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & ((\registerArray[25][5]~q ))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[17][5]~q ))))

	.dataa(\registerArray[17][5]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[25][5]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux58~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~0 .lut_mask = 16'hFC22;
defparam \Mux58~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N13
dffeas \registerArray[29][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][5] .is_wysiwyg = "true";
defparam \registerArray[29][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N20
cycloneive_lcell_comb \Mux58~1 (
// Equation(s):
// \Mux58~1_combout  = (\Mux58~0_combout  & (((\registerArray[29][5]~q ) # (!\my_rf.rsel2[2]~input_o )))) # (!\Mux58~0_combout  & (\registerArray[21][5]~q  & (\my_rf.rsel2[2]~input_o )))

	.dataa(\registerArray[21][5]~q ),
	.datab(\Mux58~0_combout ),
	.datac(\my_rf.rsel2[2]~input_o ),
	.datad(\registerArray[29][5]~q ),
	.cin(gnd),
	.combout(\Mux58~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~1 .lut_mask = 16'hEC2C;
defparam \Mux58~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y32_N29
dffeas \registerArray[27][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][5] .is_wysiwyg = "true";
defparam \registerArray[27][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N28
cycloneive_lcell_comb \Mux58~7 (
// Equation(s):
// \Mux58~7_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & ((\registerArray[27][5]~q ))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[19][5]~q ))))

	.dataa(\registerArray[19][5]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[27][5]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux58~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~7 .lut_mask = 16'hFC22;
defparam \Mux58~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y32_N25
dffeas \registerArray[23][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][5] .is_wysiwyg = "true";
defparam \registerArray[23][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N24
cycloneive_lcell_comb \Mux58~8 (
// Equation(s):
// \Mux58~8_combout  = (\Mux58~7_combout  & ((\registerArray[31][5]~q ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux58~7_combout  & (((\registerArray[23][5]~q  & \my_rf.rsel2[2]~input_o ))))

	.dataa(\registerArray[31][5]~q ),
	.datab(\Mux58~7_combout ),
	.datac(\registerArray[23][5]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux58~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~8 .lut_mask = 16'hB8CC;
defparam \Mux58~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y38_N9
dffeas \registerArray[30][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][5] .is_wysiwyg = "true";
defparam \registerArray[30][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y37_N9
dffeas \registerArray[26][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][5] .is_wysiwyg = "true";
defparam \registerArray[26][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y36_N21
dffeas \registerArray[22][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][5] .is_wysiwyg = "true";
defparam \registerArray[22][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N20
cycloneive_lcell_comb \Mux58~2 (
// Equation(s):
// \Mux58~2_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[22][5]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[18][5]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[18][5]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][5]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux58~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~2 .lut_mask = 16'hCCE2;
defparam \Mux58~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y37_N8
cycloneive_lcell_comb \Mux58~3 (
// Equation(s):
// \Mux58~3_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux58~2_combout  & (\registerArray[30][5]~q )) # (!\Mux58~2_combout  & ((\registerArray[26][5]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux58~2_combout ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[30][5]~q ),
	.datac(\registerArray[26][5]~q ),
	.datad(\Mux58~2_combout ),
	.cin(gnd),
	.combout(\Mux58~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~3 .lut_mask = 16'hDDA0;
defparam \Mux58~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y36_N25
dffeas \registerArray[20][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][5] .is_wysiwyg = "true";
defparam \registerArray[20][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N19
dffeas \registerArray[16][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][5] .is_wysiwyg = "true";
defparam \registerArray[16][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N24
cycloneive_lcell_comb \Mux58~4 (
// Equation(s):
// \Mux58~4_combout  = (\my_rf.rsel2[3]~input_o  & (\my_rf.rsel2[2]~input_o )) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\registerArray[20][5]~q )) # (!\my_rf.rsel2[2]~input_o  & ((\registerArray[16][5]~q )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[20][5]~q ),
	.datad(\registerArray[16][5]~q ),
	.cin(gnd),
	.combout(\Mux58~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~4 .lut_mask = 16'hD9C8;
defparam \Mux58~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N5
dffeas \registerArray[24][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][5] .is_wysiwyg = "true";
defparam \registerArray[24][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N4
cycloneive_lcell_comb \Mux58~5 (
// Equation(s):
// \Mux58~5_combout  = (\Mux58~4_combout  & ((\registerArray[28][5]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux58~4_combout  & (((\registerArray[24][5]~q  & \my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[28][5]~q ),
	.datab(\Mux58~4_combout ),
	.datac(\registerArray[24][5]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux58~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~5 .lut_mask = 16'hB8CC;
defparam \Mux58~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N4
cycloneive_lcell_comb \Mux58~6 (
// Equation(s):
// \Mux58~6_combout  = (\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o ) # ((\Mux58~3_combout )))) # (!\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & ((\Mux58~5_combout ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux58~3_combout ),
	.datad(\Mux58~5_combout ),
	.cin(gnd),
	.combout(\Mux58~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~6 .lut_mask = 16'hB9A8;
defparam \Mux58~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N16
cycloneive_lcell_comb \Mux58~9 (
// Equation(s):
// \Mux58~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux58~6_combout  & ((\Mux58~8_combout ))) # (!\Mux58~6_combout  & (\Mux58~1_combout )))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux58~6_combout ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\Mux58~1_combout ),
	.datac(\Mux58~8_combout ),
	.datad(\Mux58~6_combout ),
	.cin(gnd),
	.combout(\Mux58~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~9 .lut_mask = 16'hF588;
defparam \Mux58~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N30
cycloneive_lcell_comb \Mux58~20 (
// Equation(s):
// \Mux58~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux58~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux58~19_combout ))

	.dataa(\Mux58~19_combout ),
	.datab(gnd),
	.datac(\my_rf.rsel2[4]~input_o ),
	.datad(\Mux58~9_combout ),
	.cin(gnd),
	.combout(\Mux58~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~20 .lut_mask = 16'hFA0A;
defparam \Mux58~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X56_Y0_N1
cycloneive_io_ibuf \my_rf.wdat[6]~input (
	.i(\my_rf.wdat [6]),
	.ibar(gnd),
	.o(\my_rf.wdat[6]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[6]~input .bus_hold = "false";
defparam \my_rf.wdat[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X49_Y31_N1
dffeas \registerArray[9][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][6] .is_wysiwyg = "true";
defparam \registerArray[9][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y31_N17
dffeas \registerArray[10][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][6] .is_wysiwyg = "true";
defparam \registerArray[10][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y31_N19
dffeas \registerArray[8][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][6] .is_wysiwyg = "true";
defparam \registerArray[8][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N16
cycloneive_lcell_comb \Mux57~10 (
// Equation(s):
// \Mux57~10_combout  = (\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o ) # ((\registerArray[10][6]~q )))) # (!\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & ((\registerArray[8][6]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[10][6]~q ),
	.datad(\registerArray[8][6]~q ),
	.cin(gnd),
	.combout(\Mux57~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~10 .lut_mask = 16'hB9A8;
defparam \Mux57~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N0
cycloneive_lcell_comb \Mux57~11 (
// Equation(s):
// \Mux57~11_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux57~10_combout  & (\registerArray[11][6]~q )) # (!\Mux57~10_combout  & ((\registerArray[9][6]~q ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux57~10_combout ))))

	.dataa(\registerArray[11][6]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[9][6]~q ),
	.datad(\Mux57~10_combout ),
	.cin(gnd),
	.combout(\Mux57~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~11 .lut_mask = 16'hBBC0;
defparam \Mux57~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N9
dffeas \registerArray[6][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][6] .is_wysiwyg = "true";
defparam \registerArray[6][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N25
dffeas \registerArray[7][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][6] .is_wysiwyg = "true";
defparam \registerArray[7][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N8
cycloneive_lcell_comb \Mux57~13 (
// Equation(s):
// \Mux57~13_combout  = (\Mux57~12_combout  & (((\registerArray[7][6]~q )) # (!\my_rf.rsel2[1]~input_o ))) # (!\Mux57~12_combout  & (\my_rf.rsel2[1]~input_o  & (\registerArray[6][6]~q )))

	.dataa(\Mux57~12_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[6][6]~q ),
	.datad(\registerArray[7][6]~q ),
	.cin(gnd),
	.combout(\Mux57~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~13 .lut_mask = 16'hEA62;
defparam \Mux57~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N18
cycloneive_lcell_comb \Mux57~16 (
// Equation(s):
// \Mux57~16_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o ) # (\Mux57~13_combout )))) # (!\my_rf.rsel2[2]~input_o  & (\Mux57~15_combout  & (!\my_rf.rsel2[3]~input_o )))

	.dataa(\Mux57~15_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\my_rf.rsel2[3]~input_o ),
	.datad(\Mux57~13_combout ),
	.cin(gnd),
	.combout(\Mux57~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~16 .lut_mask = 16'hCEC2;
defparam \Mux57~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N6
cycloneive_lcell_comb \Mux57~19 (
// Equation(s):
// \Mux57~19_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux57~16_combout  & (\Mux57~18_combout )) # (!\Mux57~16_combout  & ((\Mux57~11_combout ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux57~16_combout ))))

	.dataa(\Mux57~18_combout ),
	.datab(\Mux57~11_combout ),
	.datac(\my_rf.rsel2[3]~input_o ),
	.datad(\Mux57~16_combout ),
	.cin(gnd),
	.combout(\Mux57~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~19 .lut_mask = 16'hAFC0;
defparam \Mux57~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y32_N11
dffeas \registerArray[23][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][6] .is_wysiwyg = "true";
defparam \registerArray[23][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y33_N9
dffeas \registerArray[19][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][6] .is_wysiwyg = "true";
defparam \registerArray[19][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N10
cycloneive_lcell_comb \Mux57~7 (
// Equation(s):
// \Mux57~7_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[23][6]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[19][6]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[23][6]~q ),
	.datad(\registerArray[19][6]~q ),
	.cin(gnd),
	.combout(\Mux57~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~7 .lut_mask = 16'hB9A8;
defparam \Mux57~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y32_N1
dffeas \registerArray[27][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][6] .is_wysiwyg = "true";
defparam \registerArray[27][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N0
cycloneive_lcell_comb \Mux57~8 (
// Equation(s):
// \Mux57~8_combout  = (\Mux57~7_combout  & ((\registerArray[31][6]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux57~7_combout  & (((\registerArray[27][6]~q  & \my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[31][6]~q ),
	.datab(\Mux57~7_combout ),
	.datac(\registerArray[27][6]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux57~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~8 .lut_mask = 16'hB8CC;
defparam \Mux57~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y36_N29
dffeas \registerArray[20][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][6] .is_wysiwyg = "true";
defparam \registerArray[20][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N1
dffeas \registerArray[24][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][6] .is_wysiwyg = "true";
defparam \registerArray[24][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N0
cycloneive_lcell_comb \Mux57~4 (
// Equation(s):
// \Mux57~4_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & ((\registerArray[24][6]~q ))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[16][6]~q ))))

	.dataa(\registerArray[16][6]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[24][6]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux57~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~4 .lut_mask = 16'hFC22;
defparam \Mux57~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N28
cycloneive_lcell_comb \Mux57~5 (
// Equation(s):
// \Mux57~5_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux57~4_combout  & (\registerArray[28][6]~q )) # (!\Mux57~4_combout  & ((\registerArray[20][6]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux57~4_combout ))))

	.dataa(\registerArray[28][6]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[20][6]~q ),
	.datad(\Mux57~4_combout ),
	.cin(gnd),
	.combout(\Mux57~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~5 .lut_mask = 16'hBBC0;
defparam \Mux57~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N12
cycloneive_lcell_comb \Mux57~6 (
// Equation(s):
// \Mux57~6_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux57~3_combout ) # ((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux57~5_combout  & !\my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux57~3_combout ),
	.datab(\Mux57~5_combout ),
	.datac(\my_rf.rsel2[1]~input_o ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux57~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~6 .lut_mask = 16'hF0AC;
defparam \Mux57~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N30
cycloneive_lcell_comb \Mux57~9 (
// Equation(s):
// \Mux57~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux57~6_combout  & ((\Mux57~8_combout ))) # (!\Mux57~6_combout  & (\Mux57~1_combout )))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux57~6_combout ))))

	.dataa(\Mux57~1_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux57~8_combout ),
	.datad(\Mux57~6_combout ),
	.cin(gnd),
	.combout(\Mux57~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~9 .lut_mask = 16'hF388;
defparam \Mux57~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N0
cycloneive_lcell_comb \Mux57~20 (
// Equation(s):
// \Mux57~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux57~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux57~19_combout ))

	.dataa(\Mux57~19_combout ),
	.datab(\my_rf.rsel2[4]~input_o ),
	.datac(gnd),
	.datad(\Mux57~9_combout ),
	.cin(gnd),
	.combout(\Mux57~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~20 .lut_mask = 16'hEE22;
defparam \Mux57~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N8
cycloneive_io_ibuf \my_rf.wdat[7]~input (
	.i(\my_rf.wdat [7]),
	.ibar(gnd),
	.o(\my_rf.wdat[7]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[7]~input .bus_hold = "false";
defparam \my_rf.wdat[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X46_Y36_N15
dffeas \registerArray[30][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][7] .is_wysiwyg = "true";
defparam \registerArray[30][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y36_N21
dffeas \registerArray[26][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][7] .is_wysiwyg = "true";
defparam \registerArray[26][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y36_N5
dffeas \registerArray[22][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][7] .is_wysiwyg = "true";
defparam \registerArray[22][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y32_N4
cycloneive_lcell_comb \Decoder0~10 (
// Equation(s):
// \Decoder0~10_combout  = (\my_rf.wsel[4]~input_o  & (!\my_rf.wsel[2]~input_o  & \Decoder0~6_combout ))

	.dataa(gnd),
	.datab(\my_rf.wsel[4]~input_o ),
	.datac(\my_rf.wsel[2]~input_o ),
	.datad(\Decoder0~6_combout ),
	.cin(gnd),
	.combout(\Decoder0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~10 .lut_mask = 16'h0C00;
defparam \Decoder0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N7
dffeas \registerArray[18][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][7] .is_wysiwyg = "true";
defparam \registerArray[18][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N4
cycloneive_lcell_comb \Mux56~2 (
// Equation(s):
// \Mux56~2_combout  = (\my_rf.rsel2[3]~input_o  & (\my_rf.rsel2[2]~input_o )) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\registerArray[22][7]~q )) # (!\my_rf.rsel2[2]~input_o  & ((\registerArray[18][7]~q )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][7]~q ),
	.datad(\registerArray[18][7]~q ),
	.cin(gnd),
	.combout(\Mux56~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~2 .lut_mask = 16'hD9C8;
defparam \Mux56~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N20
cycloneive_lcell_comb \Mux56~3 (
// Equation(s):
// \Mux56~3_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux56~2_combout  & (\registerArray[30][7]~q )) # (!\Mux56~2_combout  & ((\registerArray[26][7]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux56~2_combout ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[30][7]~q ),
	.datac(\registerArray[26][7]~q ),
	.datad(\Mux56~2_combout ),
	.cin(gnd),
	.combout(\Mux56~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~3 .lut_mask = 16'hDDA0;
defparam \Mux56~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y36_N17
dffeas \registerArray[20][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][7] .is_wysiwyg = "true";
defparam \registerArray[20][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N11
dffeas \registerArray[16][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][7] .is_wysiwyg = "true";
defparam \registerArray[16][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N16
cycloneive_lcell_comb \Mux56~4 (
// Equation(s):
// \Mux56~4_combout  = (\my_rf.rsel2[3]~input_o  & (\my_rf.rsel2[2]~input_o )) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\registerArray[20][7]~q )) # (!\my_rf.rsel2[2]~input_o  & ((\registerArray[16][7]~q )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[20][7]~q ),
	.datad(\registerArray[16][7]~q ),
	.cin(gnd),
	.combout(\Mux56~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~4 .lut_mask = 16'hD9C8;
defparam \Mux56~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N21
dffeas \registerArray[24][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][7] .is_wysiwyg = "true";
defparam \registerArray[24][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N20
cycloneive_lcell_comb \Mux56~5 (
// Equation(s):
// \Mux56~5_combout  = (\Mux56~4_combout  & ((\registerArray[28][7]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux56~4_combout  & (((\registerArray[24][7]~q  & \my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[28][7]~q ),
	.datab(\Mux56~4_combout ),
	.datac(\registerArray[24][7]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux56~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~5 .lut_mask = 16'hB8CC;
defparam \Mux56~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N14
cycloneive_lcell_comb \Mux56~6 (
// Equation(s):
// \Mux56~6_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux56~3_combout ) # ((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux56~5_combout  & !\my_rf.rsel2[0]~input_o ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux56~3_combout ),
	.datac(\Mux56~5_combout ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux56~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~6 .lut_mask = 16'hAAD8;
defparam \Mux56~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y33_N1
dffeas \registerArray[23][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][7] .is_wysiwyg = "true";
defparam \registerArray[23][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N19
dffeas \registerArray[31][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][7] .is_wysiwyg = "true";
defparam \registerArray[31][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N0
cycloneive_lcell_comb \Mux56~8 (
// Equation(s):
// \Mux56~8_combout  = (\Mux56~7_combout  & (((\registerArray[31][7]~q )) # (!\my_rf.rsel2[2]~input_o ))) # (!\Mux56~7_combout  & (\my_rf.rsel2[2]~input_o  & (\registerArray[23][7]~q )))

	.dataa(\Mux56~7_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[23][7]~q ),
	.datad(\registerArray[31][7]~q ),
	.cin(gnd),
	.combout(\Mux56~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~8 .lut_mask = 16'hEA62;
defparam \Mux56~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N0
cycloneive_lcell_comb \Mux56~9 (
// Equation(s):
// \Mux56~9_combout  = (\Mux56~6_combout  & (((\Mux56~8_combout ) # (!\my_rf.rsel2[0]~input_o )))) # (!\Mux56~6_combout  & (\Mux56~1_combout  & ((\my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux56~1_combout ),
	.datab(\Mux56~6_combout ),
	.datac(\Mux56~8_combout ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux56~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~9 .lut_mask = 16'hE2CC;
defparam \Mux56~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N1
dffeas \registerArray[3][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][7] .is_wysiwyg = "true";
defparam \registerArray[3][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y31_N26
cycloneive_lcell_comb \Decoder0~33 (
// Equation(s):
// \Decoder0~33_combout  = (!\my_rf.wsel[3]~input_o  & (!\my_rf.wsel[4]~input_o  & \Decoder0~0_combout ))

	.dataa(\my_rf.wsel[3]~input_o ),
	.datab(gnd),
	.datac(\my_rf.wsel[4]~input_o ),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~33_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~33 .lut_mask = 16'h0500;
defparam \Decoder0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N27
dffeas \registerArray[1][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][7] .is_wysiwyg = "true";
defparam \registerArray[1][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N0
cycloneive_lcell_comb \Mux56~14 (
// Equation(s):
// \Mux56~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][7]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][7]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][7]~q ),
	.datad(\registerArray[1][7]~q ),
	.cin(gnd),
	.combout(\Mux56~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~14 .lut_mask = 16'hC480;
defparam \Mux56~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N31
dffeas \registerArray[2][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][7] .is_wysiwyg = "true";
defparam \registerArray[2][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N30
cycloneive_lcell_comb \Mux56~15 (
// Equation(s):
// \Mux56~15_combout  = (\Mux56~14_combout ) # ((!\my_rf.rsel2[0]~input_o  & (\registerArray[2][7]~q  & \my_rf.rsel2[1]~input_o )))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\Mux56~14_combout ),
	.datac(\registerArray[2][7]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux56~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~15 .lut_mask = 16'hDCCC;
defparam \Mux56~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N26
cycloneive_lcell_comb \Mux56~16 (
// Equation(s):
// \Mux56~16_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux56~13_combout ) # ((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux56~15_combout  & !\my_rf.rsel2[2]~input_o ))))

	.dataa(\Mux56~13_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux56~15_combout ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux56~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~16 .lut_mask = 16'hCCB8;
defparam \Mux56~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y29_N25
dffeas \registerArray[6][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][7] .is_wysiwyg = "true";
defparam \registerArray[6][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N5
dffeas \registerArray[5][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][7] .is_wysiwyg = "true";
defparam \registerArray[5][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N4
cycloneive_lcell_comb \Mux56~10 (
// Equation(s):
// \Mux56~10_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[5][7]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][7]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[4][7]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][7]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux56~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~10 .lut_mask = 16'hCCE2;
defparam \Mux56~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N24
cycloneive_lcell_comb \Mux56~11 (
// Equation(s):
// \Mux56~11_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux56~10_combout  & (\registerArray[7][7]~q )) # (!\Mux56~10_combout  & ((\registerArray[6][7]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux56~10_combout ))))

	.dataa(\registerArray[7][7]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[6][7]~q ),
	.datad(\Mux56~10_combout ),
	.cin(gnd),
	.combout(\Mux56~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~11 .lut_mask = 16'hBBC0;
defparam \Mux56~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N20
cycloneive_lcell_comb \Mux56~19 (
// Equation(s):
// \Mux56~19_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux56~16_combout  & (\Mux56~18_combout )) # (!\Mux56~16_combout  & ((\Mux56~11_combout ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux56~16_combout ))))

	.dataa(\Mux56~18_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\Mux56~16_combout ),
	.datad(\Mux56~11_combout ),
	.cin(gnd),
	.combout(\Mux56~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~19 .lut_mask = 16'hBCB0;
defparam \Mux56~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N6
cycloneive_lcell_comb \Mux56~20 (
// Equation(s):
// \Mux56~20_combout  = (\my_rf.rsel2[4]~input_o  & (\Mux56~9_combout )) # (!\my_rf.rsel2[4]~input_o  & ((\Mux56~19_combout )))

	.dataa(\my_rf.rsel2[4]~input_o ),
	.datab(\Mux56~9_combout ),
	.datac(gnd),
	.datad(\Mux56~19_combout ),
	.cin(gnd),
	.combout(\Mux56~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~20 .lut_mask = 16'hDD88;
defparam \Mux56~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X56_Y0_N8
cycloneive_io_ibuf \my_rf.wdat[8]~input (
	.i(\my_rf.wdat [8]),
	.ibar(gnd),
	.o(\my_rf.wdat[8]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[8]~input .bus_hold = "false";
defparam \my_rf.wdat[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X50_Y36_N1
dffeas \registerArray[13][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][8] .is_wysiwyg = "true";
defparam \registerArray[13][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N11
dffeas \registerArray[12][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][8] .is_wysiwyg = "true";
defparam \registerArray[12][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N0
cycloneive_lcell_comb \Mux55~17 (
// Equation(s):
// \Mux55~17_combout  = (\my_rf.rsel2[1]~input_o  & (\my_rf.rsel2[0]~input_o )) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & (\registerArray[13][8]~q )) # (!\my_rf.rsel2[0]~input_o  & ((\registerArray[12][8]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[13][8]~q ),
	.datad(\registerArray[12][8]~q ),
	.cin(gnd),
	.combout(\Mux55~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~17 .lut_mask = 16'hD9C8;
defparam \Mux55~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N3
dffeas \registerArray[14][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][8] .is_wysiwyg = "true";
defparam \registerArray[14][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N21
dffeas \registerArray[15][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][8] .is_wysiwyg = "true";
defparam \registerArray[15][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N2
cycloneive_lcell_comb \Mux55~18 (
// Equation(s):
// \Mux55~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux55~17_combout  & ((\registerArray[15][8]~q ))) # (!\Mux55~17_combout  & (\registerArray[14][8]~q )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux55~17_combout ))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux55~17_combout ),
	.datac(\registerArray[14][8]~q ),
	.datad(\registerArray[15][8]~q ),
	.cin(gnd),
	.combout(\Mux55~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~18 .lut_mask = 16'hEC64;
defparam \Mux55~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N11
dffeas \registerArray[2][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][8] .is_wysiwyg = "true";
defparam \registerArray[2][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N10
cycloneive_lcell_comb \Mux55~15 (
// Equation(s):
// \Mux55~15_combout  = (\Mux55~14_combout ) # ((!\my_rf.rsel2[0]~input_o  & (\registerArray[2][8]~q  & \my_rf.rsel2[1]~input_o )))

	.dataa(\Mux55~14_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][8]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux55~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~15 .lut_mask = 16'hBAAA;
defparam \Mux55~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N1
dffeas \registerArray[5][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][8] .is_wysiwyg = "true";
defparam \registerArray[5][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N0
cycloneive_lcell_comb \Mux55~12 (
// Equation(s):
// \Mux55~12_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[5][8]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][8]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[4][8]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][8]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux55~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~12 .lut_mask = 16'hCCE2;
defparam \Mux55~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N3
dffeas \registerArray[6][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][8] .is_wysiwyg = "true";
defparam \registerArray[6][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N29
dffeas \registerArray[7][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][8] .is_wysiwyg = "true";
defparam \registerArray[7][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N2
cycloneive_lcell_comb \Mux55~13 (
// Equation(s):
// \Mux55~13_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux55~12_combout  & ((\registerArray[7][8]~q ))) # (!\Mux55~12_combout  & (\registerArray[6][8]~q )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux55~12_combout ))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux55~12_combout ),
	.datac(\registerArray[6][8]~q ),
	.datad(\registerArray[7][8]~q ),
	.cin(gnd),
	.combout(\Mux55~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~13 .lut_mask = 16'hEC64;
defparam \Mux55~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N4
cycloneive_lcell_comb \Mux55~16 (
// Equation(s):
// \Mux55~16_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\Mux55~13_combout )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & (\Mux55~15_combout )))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux55~15_combout ),
	.datad(\Mux55~13_combout ),
	.cin(gnd),
	.combout(\Mux55~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~16 .lut_mask = 16'hBA98;
defparam \Mux55~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y37_N1
dffeas \registerArray[9][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][8] .is_wysiwyg = "true";
defparam \registerArray[9][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y37_N25
dffeas \registerArray[10][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][8] .is_wysiwyg = "true";
defparam \registerArray[10][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y37_N24
cycloneive_lcell_comb \Mux55~10 (
// Equation(s):
// \Mux55~10_combout  = (\my_rf.rsel2[0]~input_o  & (((\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[10][8]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[8][8]~q ))))

	.dataa(\registerArray[8][8]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[10][8]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux55~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~10 .lut_mask = 16'hFC22;
defparam \Mux55~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y37_N0
cycloneive_lcell_comb \Mux55~11 (
// Equation(s):
// \Mux55~11_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux55~10_combout  & (\registerArray[11][8]~q )) # (!\Mux55~10_combout  & ((\registerArray[9][8]~q ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux55~10_combout ))))

	.dataa(\registerArray[11][8]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[9][8]~q ),
	.datad(\Mux55~10_combout ),
	.cin(gnd),
	.combout(\Mux55~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~11 .lut_mask = 16'hBBC0;
defparam \Mux55~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N22
cycloneive_lcell_comb \Mux55~19 (
// Equation(s):
// \Mux55~19_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux55~16_combout  & (\Mux55~18_combout )) # (!\Mux55~16_combout  & ((\Mux55~11_combout ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux55~16_combout ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux55~18_combout ),
	.datac(\Mux55~16_combout ),
	.datad(\Mux55~11_combout ),
	.cin(gnd),
	.combout(\Mux55~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~19 .lut_mask = 16'hDAD0;
defparam \Mux55~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y32_N5
dffeas \registerArray[21][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][8] .is_wysiwyg = "true";
defparam \registerArray[21][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N11
dffeas \registerArray[17][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][8] .is_wysiwyg = "true";
defparam \registerArray[17][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N4
cycloneive_lcell_comb \Mux55~0 (
// Equation(s):
// \Mux55~0_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[21][8]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[17][8]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[21][8]~q ),
	.datad(\registerArray[17][8]~q ),
	.cin(gnd),
	.combout(\Mux55~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~0 .lut_mask = 16'hB9A8;
defparam \Mux55~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y0_N10
dffeas \registerArray[25][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[8]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][8] .is_wysiwyg = "true";
defparam \registerArray[25][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y36_N27
dffeas \registerArray[29][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][8] .is_wysiwyg = "true";
defparam \registerArray[29][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N22
cycloneive_lcell_comb \Mux55~1 (
// Equation(s):
// \Mux55~1_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux55~0_combout  & ((\registerArray[29][8]~q ))) # (!\Mux55~0_combout  & (\registerArray[25][8]~q )))) # (!\my_rf.rsel2[3]~input_o  & (\Mux55~0_combout ))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux55~0_combout ),
	.datac(\registerArray[25][8]~q ),
	.datad(\registerArray[29][8]~q ),
	.cin(gnd),
	.combout(\Mux55~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~1 .lut_mask = 16'hEC64;
defparam \Mux55~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N25
dffeas \registerArray[20][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][8] .is_wysiwyg = "true";
defparam \registerArray[20][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y37_N3
dffeas \registerArray[28][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][8] .is_wysiwyg = "true";
defparam \registerArray[28][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N24
cycloneive_lcell_comb \Mux55~5 (
// Equation(s):
// \Mux55~5_combout  = (\Mux55~4_combout  & (((\registerArray[28][8]~q )) # (!\my_rf.rsel2[2]~input_o ))) # (!\Mux55~4_combout  & (\my_rf.rsel2[2]~input_o  & (\registerArray[20][8]~q )))

	.dataa(\Mux55~4_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[20][8]~q ),
	.datad(\registerArray[28][8]~q ),
	.cin(gnd),
	.combout(\Mux55~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~5 .lut_mask = 16'hEA62;
defparam \Mux55~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N9
dffeas \registerArray[22][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][8] .is_wysiwyg = "true";
defparam \registerArray[22][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y36_N27
dffeas \registerArray[30][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][8] .is_wysiwyg = "true";
defparam \registerArray[30][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N8
cycloneive_lcell_comb \Mux55~3 (
// Equation(s):
// \Mux55~3_combout  = (\Mux55~2_combout  & (((\registerArray[30][8]~q )) # (!\my_rf.rsel2[2]~input_o ))) # (!\Mux55~2_combout  & (\my_rf.rsel2[2]~input_o  & (\registerArray[22][8]~q )))

	.dataa(\Mux55~2_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][8]~q ),
	.datad(\registerArray[30][8]~q ),
	.cin(gnd),
	.combout(\Mux55~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~3 .lut_mask = 16'hEA62;
defparam \Mux55~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N16
cycloneive_lcell_comb \Mux55~6 (
// Equation(s):
// \Mux55~6_combout  = (\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o ) # ((\Mux55~3_combout )))) # (!\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & (\Mux55~5_combout )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux55~5_combout ),
	.datad(\Mux55~3_combout ),
	.cin(gnd),
	.combout(\Mux55~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~6 .lut_mask = 16'hBA98;
defparam \Mux55~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N2
cycloneive_lcell_comb \Mux55~9 (
// Equation(s):
// \Mux55~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux55~6_combout  & (\Mux55~8_combout )) # (!\Mux55~6_combout  & ((\Mux55~1_combout ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux55~6_combout ))))

	.dataa(\Mux55~8_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux55~1_combout ),
	.datad(\Mux55~6_combout ),
	.cin(gnd),
	.combout(\Mux55~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~9 .lut_mask = 16'hBBC0;
defparam \Mux55~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N8
cycloneive_lcell_comb \Mux55~20 (
// Equation(s):
// \Mux55~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux55~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux55~19_combout ))

	.dataa(\my_rf.rsel2[4]~input_o ),
	.datab(gnd),
	.datac(\Mux55~19_combout ),
	.datad(\Mux55~9_combout ),
	.cin(gnd),
	.combout(\Mux55~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~20 .lut_mask = 16'hFA50;
defparam \Mux55~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N1
cycloneive_io_ibuf \my_rf.wdat[9]~input (
	.i(\my_rf.wdat [9]),
	.ibar(gnd),
	.o(\my_rf.wdat[9]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[9]~input .bus_hold = "false";
defparam \my_rf.wdat[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X53_Y35_N7
dffeas \registerArray[2][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][9] .is_wysiwyg = "true";
defparam \registerArray[2][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N6
cycloneive_lcell_comb \Mux54~15 (
// Equation(s):
// \Mux54~15_combout  = (\Mux54~14_combout ) # ((!\my_rf.rsel2[0]~input_o  & (\registerArray[2][9]~q  & \my_rf.rsel2[1]~input_o )))

	.dataa(\Mux54~14_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][9]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux54~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~15 .lut_mask = 16'hBAAA;
defparam \Mux54~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N4
cycloneive_lcell_comb \Mux54~16 (
// Equation(s):
// \Mux54~16_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\Mux54~13_combout )) # (!\my_rf.rsel2[3]~input_o  & ((\Mux54~15_combout )))))

	.dataa(\Mux54~13_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\my_rf.rsel2[3]~input_o ),
	.datad(\Mux54~15_combout ),
	.cin(gnd),
	.combout(\Mux54~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~16 .lut_mask = 16'hE3E0;
defparam \Mux54~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N3
dffeas \registerArray[6][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][9] .is_wysiwyg = "true";
defparam \registerArray[6][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N23
dffeas \registerArray[7][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][9] .is_wysiwyg = "true";
defparam \registerArray[7][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N2
cycloneive_lcell_comb \Mux54~11 (
// Equation(s):
// \Mux54~11_combout  = (\Mux54~10_combout  & (((\registerArray[7][9]~q )) # (!\my_rf.rsel2[1]~input_o ))) # (!\Mux54~10_combout  & (\my_rf.rsel2[1]~input_o  & (\registerArray[6][9]~q )))

	.dataa(\Mux54~10_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[6][9]~q ),
	.datad(\registerArray[7][9]~q ),
	.cin(gnd),
	.combout(\Mux54~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~11 .lut_mask = 16'hEA62;
defparam \Mux54~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N14
cycloneive_lcell_comb \Mux54~19 (
// Equation(s):
// \Mux54~19_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux54~16_combout  & (\Mux54~18_combout )) # (!\Mux54~16_combout  & ((\Mux54~11_combout ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux54~16_combout ))))

	.dataa(\Mux54~18_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\Mux54~16_combout ),
	.datad(\Mux54~11_combout ),
	.cin(gnd),
	.combout(\Mux54~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~19 .lut_mask = 16'hBCB0;
defparam \Mux54~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y33_N17
dffeas \registerArray[23][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][9] .is_wysiwyg = "true";
defparam \registerArray[23][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N13
dffeas \registerArray[27][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][9] .is_wysiwyg = "true";
defparam \registerArray[27][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N12
cycloneive_lcell_comb \Mux54~7 (
// Equation(s):
// \Mux54~7_combout  = (\my_rf.rsel2[3]~input_o  & (((\registerArray[27][9]~q ) # (\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[19][9]~q  & ((!\my_rf.rsel2[2]~input_o ))))

	.dataa(\registerArray[19][9]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][9]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux54~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~7 .lut_mask = 16'hCCE2;
defparam \Mux54~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N16
cycloneive_lcell_comb \Mux54~8 (
// Equation(s):
// \Mux54~8_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux54~7_combout  & (\registerArray[31][9]~q )) # (!\Mux54~7_combout  & ((\registerArray[23][9]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux54~7_combout ))))

	.dataa(\registerArray[31][9]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[23][9]~q ),
	.datad(\Mux54~7_combout ),
	.cin(gnd),
	.combout(\Mux54~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~8 .lut_mask = 16'hBBC0;
defparam \Mux54~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y36_N13
dffeas \registerArray[20][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][9] .is_wysiwyg = "true";
defparam \registerArray[20][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N12
cycloneive_lcell_comb \Mux54~4 (
// Equation(s):
// \Mux54~4_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[20][9]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[16][9]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[16][9]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[20][9]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux54~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~4 .lut_mask = 16'hCCE2;
defparam \Mux54~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N17
dffeas \registerArray[24][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][9] .is_wysiwyg = "true";
defparam \registerArray[24][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N16
cycloneive_lcell_comb \Mux54~5 (
// Equation(s):
// \Mux54~5_combout  = (\Mux54~4_combout  & ((\registerArray[28][9]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux54~4_combout  & (((\registerArray[24][9]~q  & \my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[28][9]~q ),
	.datab(\Mux54~4_combout ),
	.datac(\registerArray[24][9]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux54~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~5 .lut_mask = 16'hB8CC;
defparam \Mux54~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y36_N29
dffeas \registerArray[26][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][9] .is_wysiwyg = "true";
defparam \registerArray[26][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y36_N17
dffeas \registerArray[22][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][9] .is_wysiwyg = "true";
defparam \registerArray[22][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y36_N3
dffeas \registerArray[18][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][9] .is_wysiwyg = "true";
defparam \registerArray[18][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N16
cycloneive_lcell_comb \Mux54~2 (
// Equation(s):
// \Mux54~2_combout  = (\my_rf.rsel2[3]~input_o  & (\my_rf.rsel2[2]~input_o )) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\registerArray[22][9]~q )) # (!\my_rf.rsel2[2]~input_o  & ((\registerArray[18][9]~q )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][9]~q ),
	.datad(\registerArray[18][9]~q ),
	.cin(gnd),
	.combout(\Mux54~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~2 .lut_mask = 16'hD9C8;
defparam \Mux54~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N28
cycloneive_lcell_comb \Mux54~3 (
// Equation(s):
// \Mux54~3_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux54~2_combout  & (\registerArray[30][9]~q )) # (!\Mux54~2_combout  & ((\registerArray[26][9]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux54~2_combout ))))

	.dataa(\registerArray[30][9]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[26][9]~q ),
	.datad(\Mux54~2_combout ),
	.cin(gnd),
	.combout(\Mux54~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~3 .lut_mask = 16'hBBC0;
defparam \Mux54~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N22
cycloneive_lcell_comb \Mux54~6 (
// Equation(s):
// \Mux54~6_combout  = (\my_rf.rsel2[0]~input_o  & (\my_rf.rsel2[1]~input_o )) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\Mux54~3_combout ))) # (!\my_rf.rsel2[1]~input_o  & (\Mux54~5_combout ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\Mux54~5_combout ),
	.datad(\Mux54~3_combout ),
	.cin(gnd),
	.combout(\Mux54~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~6 .lut_mask = 16'hDC98;
defparam \Mux54~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N23
dffeas \registerArray[29][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][9] .is_wysiwyg = "true";
defparam \registerArray[29][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y0_N3
dffeas \registerArray[21][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[9]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][9] .is_wysiwyg = "true";
defparam \registerArray[21][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N0
cycloneive_lcell_comb \Mux54~1 (
// Equation(s):
// \Mux54~1_combout  = (\Mux54~0_combout  & ((\registerArray[29][9]~q ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux54~0_combout  & (((\registerArray[21][9]~q  & \my_rf.rsel2[2]~input_o ))))

	.dataa(\Mux54~0_combout ),
	.datab(\registerArray[29][9]~q ),
	.datac(\registerArray[21][9]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux54~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~1 .lut_mask = 16'hD8AA;
defparam \Mux54~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N16
cycloneive_lcell_comb \Mux54~9 (
// Equation(s):
// \Mux54~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux54~6_combout  & (\Mux54~8_combout )) # (!\Mux54~6_combout  & ((\Mux54~1_combout ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux54~6_combout ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\Mux54~8_combout ),
	.datac(\Mux54~6_combout ),
	.datad(\Mux54~1_combout ),
	.cin(gnd),
	.combout(\Mux54~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~9 .lut_mask = 16'hDAD0;
defparam \Mux54~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N24
cycloneive_lcell_comb \Mux54~20 (
// Equation(s):
// \Mux54~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux54~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux54~19_combout ))

	.dataa(gnd),
	.datab(\my_rf.rsel2[4]~input_o ),
	.datac(\Mux54~19_combout ),
	.datad(\Mux54~9_combout ),
	.cin(gnd),
	.combout(\Mux54~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~20 .lut_mask = 16'hFC30;
defparam \Mux54~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X47_Y0_N1
cycloneive_io_ibuf \my_rf.wdat[10]~input (
	.i(\my_rf.wdat [10]),
	.ibar(gnd),
	.o(\my_rf.wdat[10]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[10]~input .bus_hold = "false";
defparam \my_rf.wdat[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X54_Y37_N1
dffeas \registerArray[5][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][10] .is_wysiwyg = "true";
defparam \registerArray[5][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y31_N10
cycloneive_lcell_comb \Decoder0~30 (
// Equation(s):
// \Decoder0~30_combout  = (!\my_rf.wsel[4]~input_o  & (!\my_rf.wsel[3]~input_o  & (!\my_rf.wsel[0]~input_o  & \Decoder0~12_combout )))

	.dataa(\my_rf.wsel[4]~input_o ),
	.datab(\my_rf.wsel[3]~input_o ),
	.datac(\my_rf.wsel[0]~input_o ),
	.datad(\Decoder0~12_combout ),
	.cin(gnd),
	.combout(\Decoder0~30_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~30 .lut_mask = 16'h0100;
defparam \Decoder0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N3
dffeas \registerArray[4][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][10] .is_wysiwyg = "true";
defparam \registerArray[4][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N0
cycloneive_lcell_comb \Mux53~12 (
// Equation(s):
// \Mux53~12_combout  = (\my_rf.rsel2[1]~input_o  & (\my_rf.rsel2[0]~input_o )) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & (\registerArray[5][10]~q )) # (!\my_rf.rsel2[0]~input_o  & ((\registerArray[4][10]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][10]~q ),
	.datad(\registerArray[4][10]~q ),
	.cin(gnd),
	.combout(\Mux53~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~12 .lut_mask = 16'hD9C8;
defparam \Mux53~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N17
dffeas \registerArray[6][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][10] .is_wysiwyg = "true";
defparam \registerArray[6][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N11
dffeas \registerArray[7][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][10] .is_wysiwyg = "true";
defparam \registerArray[7][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N16
cycloneive_lcell_comb \Mux53~13 (
// Equation(s):
// \Mux53~13_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux53~12_combout  & ((\registerArray[7][10]~q ))) # (!\Mux53~12_combout  & (\registerArray[6][10]~q )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux53~12_combout ))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux53~12_combout ),
	.datac(\registerArray[6][10]~q ),
	.datad(\registerArray[7][10]~q ),
	.cin(gnd),
	.combout(\Mux53~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~13 .lut_mask = 16'hEC64;
defparam \Mux53~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N17
dffeas \registerArray[2][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][10] .is_wysiwyg = "true";
defparam \registerArray[2][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N13
dffeas \registerArray[3][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][10] .is_wysiwyg = "true";
defparam \registerArray[3][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N7
dffeas \registerArray[1][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][10] .is_wysiwyg = "true";
defparam \registerArray[1][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N12
cycloneive_lcell_comb \Mux53~14 (
// Equation(s):
// \Mux53~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][10]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][10]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][10]~q ),
	.datad(\registerArray[1][10]~q ),
	.cin(gnd),
	.combout(\Mux53~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~14 .lut_mask = 16'hC480;
defparam \Mux53~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N16
cycloneive_lcell_comb \Mux53~15 (
// Equation(s):
// \Mux53~15_combout  = (\Mux53~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][10]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][10]~q ),
	.datad(\Mux53~14_combout ),
	.cin(gnd),
	.combout(\Mux53~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~15 .lut_mask = 16'hFF20;
defparam \Mux53~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N2
cycloneive_lcell_comb \Mux53~16 (
// Equation(s):
// \Mux53~16_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\Mux53~13_combout )) # (!\my_rf.rsel2[2]~input_o  & ((\Mux53~15_combout )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux53~13_combout ),
	.datac(\Mux53~15_combout ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux53~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~16 .lut_mask = 16'hEE50;
defparam \Mux53~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N15
dffeas \registerArray[15][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][10] .is_wysiwyg = "true";
defparam \registerArray[15][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N13
dffeas \registerArray[14][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][10] .is_wysiwyg = "true";
defparam \registerArray[14][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N13
dffeas \registerArray[13][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][10] .is_wysiwyg = "true";
defparam \registerArray[13][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N12
cycloneive_lcell_comb \Mux53~17 (
// Equation(s):
// \Mux53~17_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[13][10]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[12][10]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[12][10]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[13][10]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux53~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~17 .lut_mask = 16'hCCE2;
defparam \Mux53~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N12
cycloneive_lcell_comb \Mux53~18 (
// Equation(s):
// \Mux53~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux53~17_combout  & (\registerArray[15][10]~q )) # (!\Mux53~17_combout  & ((\registerArray[14][10]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux53~17_combout ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[15][10]~q ),
	.datac(\registerArray[14][10]~q ),
	.datad(\Mux53~17_combout ),
	.cin(gnd),
	.combout(\Mux53~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~18 .lut_mask = 16'hDDA0;
defparam \Mux53~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N12
cycloneive_lcell_comb \Mux53~19 (
// Equation(s):
// \Mux53~19_combout  = (\Mux53~16_combout  & (((\Mux53~18_combout ) # (!\my_rf.rsel2[3]~input_o )))) # (!\Mux53~16_combout  & (\Mux53~11_combout  & (\my_rf.rsel2[3]~input_o )))

	.dataa(\Mux53~11_combout ),
	.datab(\Mux53~16_combout ),
	.datac(\my_rf.rsel2[3]~input_o ),
	.datad(\Mux53~18_combout ),
	.cin(gnd),
	.combout(\Mux53~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~19 .lut_mask = 16'hEC2C;
defparam \Mux53~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y33_N23
dffeas \registerArray[31][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][10] .is_wysiwyg = "true";
defparam \registerArray[31][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N23
dffeas \registerArray[27][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][10] .is_wysiwyg = "true";
defparam \registerArray[27][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N29
dffeas \registerArray[23][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][10] .is_wysiwyg = "true";
defparam \registerArray[23][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y33_N23
dffeas \registerArray[19][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][10] .is_wysiwyg = "true";
defparam \registerArray[19][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N28
cycloneive_lcell_comb \Mux53~7 (
// Equation(s):
// \Mux53~7_combout  = (\my_rf.rsel2[3]~input_o  & (\my_rf.rsel2[2]~input_o )) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\registerArray[23][10]~q )) # (!\my_rf.rsel2[2]~input_o  & ((\registerArray[19][10]~q )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[23][10]~q ),
	.datad(\registerArray[19][10]~q ),
	.cin(gnd),
	.combout(\Mux53~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~7 .lut_mask = 16'hD9C8;
defparam \Mux53~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N22
cycloneive_lcell_comb \Mux53~8 (
// Equation(s):
// \Mux53~8_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux53~7_combout  & (\registerArray[31][10]~q )) # (!\Mux53~7_combout  & ((\registerArray[27][10]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux53~7_combout ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[31][10]~q ),
	.datac(\registerArray[27][10]~q ),
	.datad(\Mux53~7_combout ),
	.cin(gnd),
	.combout(\Mux53~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~8 .lut_mask = 16'hDDA0;
defparam \Mux53~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y36_N9
dffeas \registerArray[20][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][10] .is_wysiwyg = "true";
defparam \registerArray[20][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N15
dffeas \registerArray[16][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][10] .is_wysiwyg = "true";
defparam \registerArray[16][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N13
dffeas \registerArray[24][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][10] .is_wysiwyg = "true";
defparam \registerArray[24][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N12
cycloneive_lcell_comb \Mux53~4 (
// Equation(s):
// \Mux53~4_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & ((\registerArray[24][10]~q ))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[16][10]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[16][10]~q ),
	.datac(\registerArray[24][10]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux53~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~4 .lut_mask = 16'hFA44;
defparam \Mux53~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N8
cycloneive_lcell_comb \Mux53~5 (
// Equation(s):
// \Mux53~5_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux53~4_combout  & (\registerArray[28][10]~q )) # (!\Mux53~4_combout  & ((\registerArray[20][10]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux53~4_combout ))))

	.dataa(\registerArray[28][10]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[20][10]~q ),
	.datad(\Mux53~4_combout ),
	.cin(gnd),
	.combout(\Mux53~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~5 .lut_mask = 16'hBBC0;
defparam \Mux53~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N20
cycloneive_lcell_comb \Mux53~6 (
// Equation(s):
// \Mux53~6_combout  = (\my_rf.rsel2[0]~input_o  & (((\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\Mux53~3_combout )) # (!\my_rf.rsel2[1]~input_o  & ((\Mux53~5_combout )))))

	.dataa(\Mux53~3_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux53~5_combout ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux53~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~6 .lut_mask = 16'hEE30;
defparam \Mux53~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N16
cycloneive_lcell_comb \Mux53~9 (
// Equation(s):
// \Mux53~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux53~6_combout  & ((\Mux53~8_combout ))) # (!\Mux53~6_combout  & (\Mux53~1_combout )))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux53~6_combout ))))

	.dataa(\Mux53~1_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux53~8_combout ),
	.datad(\Mux53~6_combout ),
	.cin(gnd),
	.combout(\Mux53~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~9 .lut_mask = 16'hF388;
defparam \Mux53~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N14
cycloneive_lcell_comb \Mux53~20 (
// Equation(s):
// \Mux53~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux53~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux53~19_combout ))

	.dataa(\Mux53~19_combout ),
	.datab(\my_rf.rsel2[4]~input_o ),
	.datac(gnd),
	.datad(\Mux53~9_combout ),
	.cin(gnd),
	.combout(\Mux53~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~20 .lut_mask = 16'hEE22;
defparam \Mux53~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X0_Y34_N8
cycloneive_io_ibuf \my_rf.wdat[11]~input (
	.i(\my_rf.wdat [11]),
	.ibar(gnd),
	.o(\my_rf.wdat[11]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[11]~input .bus_hold = "false";
defparam \my_rf.wdat[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X46_Y36_N13
dffeas \registerArray[26][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][11] .is_wysiwyg = "true";
defparam \registerArray[26][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y36_N9
dffeas \registerArray[22][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][11] .is_wysiwyg = "true";
defparam \registerArray[22][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N8
cycloneive_lcell_comb \Mux52~2 (
// Equation(s):
// \Mux52~2_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[22][11]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[18][11]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[18][11]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][11]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux52~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~2 .lut_mask = 16'hCCE2;
defparam \Mux52~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N12
cycloneive_lcell_comb \Mux52~3 (
// Equation(s):
// \Mux52~3_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux52~2_combout  & (\registerArray[30][11]~q )) # (!\Mux52~2_combout  & ((\registerArray[26][11]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux52~2_combout ))))

	.dataa(\registerArray[30][11]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[26][11]~q ),
	.datad(\Mux52~2_combout ),
	.cin(gnd),
	.combout(\Mux52~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~3 .lut_mask = 16'hBBC0;
defparam \Mux52~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N24
cycloneive_lcell_comb \Mux52~6 (
// Equation(s):
// \Mux52~6_combout  = (\my_rf.rsel2[0]~input_o  & (((\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\Mux52~3_combout ))) # (!\my_rf.rsel2[1]~input_o  & (\Mux52~5_combout ))))

	.dataa(\Mux52~5_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\my_rf.rsel2[1]~input_o ),
	.datad(\Mux52~3_combout ),
	.cin(gnd),
	.combout(\Mux52~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~6 .lut_mask = 16'hF2C2;
defparam \Mux52~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y33_N25
dffeas \registerArray[23][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][11] .is_wysiwyg = "true";
defparam \registerArray[23][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N27
dffeas \registerArray[19][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][11] .is_wysiwyg = "true";
defparam \registerArray[19][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N1
dffeas \registerArray[27][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][11] .is_wysiwyg = "true";
defparam \registerArray[27][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N0
cycloneive_lcell_comb \Mux52~7 (
// Equation(s):
// \Mux52~7_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & ((\registerArray[27][11]~q ))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[19][11]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[19][11]~q ),
	.datac(\registerArray[27][11]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux52~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~7 .lut_mask = 16'hFA44;
defparam \Mux52~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N24
cycloneive_lcell_comb \Mux52~8 (
// Equation(s):
// \Mux52~8_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux52~7_combout  & (\registerArray[31][11]~q )) # (!\Mux52~7_combout  & ((\registerArray[23][11]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux52~7_combout ))))

	.dataa(\registerArray[31][11]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[23][11]~q ),
	.datad(\Mux52~7_combout ),
	.cin(gnd),
	.combout(\Mux52~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~8 .lut_mask = 16'hBBC0;
defparam \Mux52~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N18
cycloneive_lcell_comb \Mux52~9 (
// Equation(s):
// \Mux52~9_combout  = (\Mux52~6_combout  & (((\Mux52~8_combout ) # (!\my_rf.rsel2[0]~input_o )))) # (!\Mux52~6_combout  & (\Mux52~1_combout  & ((\my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux52~1_combout ),
	.datab(\Mux52~6_combout ),
	.datac(\Mux52~8_combout ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux52~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~9 .lut_mask = 16'hE2CC;
defparam \Mux52~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N11
dffeas \registerArray[2][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][11] .is_wysiwyg = "true";
defparam \registerArray[2][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N25
dffeas \registerArray[3][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][11] .is_wysiwyg = "true";
defparam \registerArray[3][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N19
dffeas \registerArray[1][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][11] .is_wysiwyg = "true";
defparam \registerArray[1][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N24
cycloneive_lcell_comb \Mux52~14 (
// Equation(s):
// \Mux52~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][11]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][11]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][11]~q ),
	.datad(\registerArray[1][11]~q ),
	.cin(gnd),
	.combout(\Mux52~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~14 .lut_mask = 16'hC480;
defparam \Mux52~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N10
cycloneive_lcell_comb \Mux52~15 (
// Equation(s):
// \Mux52~15_combout  = (\Mux52~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][11]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][11]~q ),
	.datad(\Mux52~14_combout ),
	.cin(gnd),
	.combout(\Mux52~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~15 .lut_mask = 16'hFF20;
defparam \Mux52~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y31_N18
cycloneive_lcell_comb \Decoder0~27 (
// Equation(s):
// \Decoder0~27_combout  = (\my_rf.wsel[3]~input_o  & (!\my_rf.wsel[2]~input_o  & (!\my_rf.wsel[4]~input_o  & \Decoder0~19_combout )))

	.dataa(\my_rf.wsel[3]~input_o ),
	.datab(\my_rf.wsel[2]~input_o ),
	.datac(\my_rf.wsel[4]~input_o ),
	.datad(\Decoder0~19_combout ),
	.cin(gnd),
	.combout(\Decoder0~27_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~27 .lut_mask = 16'h0200;
defparam \Decoder0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y37_N15
dffeas \registerArray[11][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][11] .is_wysiwyg = "true";
defparam \registerArray[11][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y37_N21
dffeas \registerArray[9][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][11] .is_wysiwyg = "true";
defparam \registerArray[9][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y37_N20
cycloneive_lcell_comb \Mux52~13 (
// Equation(s):
// \Mux52~13_combout  = (\Mux52~12_combout  & ((\registerArray[11][11]~q ) # ((!\my_rf.rsel2[0]~input_o )))) # (!\Mux52~12_combout  & (((\registerArray[9][11]~q  & \my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux52~12_combout ),
	.datab(\registerArray[11][11]~q ),
	.datac(\registerArray[9][11]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux52~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~13 .lut_mask = 16'hD8AA;
defparam \Mux52~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y37_N24
cycloneive_lcell_comb \Mux52~16 (
// Equation(s):
// \Mux52~16_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o ) # (\Mux52~13_combout )))) # (!\my_rf.rsel2[3]~input_o  & (\Mux52~15_combout  & (!\my_rf.rsel2[2]~input_o )))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux52~15_combout ),
	.datac(\my_rf.rsel2[2]~input_o ),
	.datad(\Mux52~13_combout ),
	.cin(gnd),
	.combout(\Mux52~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~16 .lut_mask = 16'hAEA4;
defparam \Mux52~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N13
dffeas \registerArray[5][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][11] .is_wysiwyg = "true";
defparam \registerArray[5][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N31
dffeas \registerArray[4][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][11] .is_wysiwyg = "true";
defparam \registerArray[4][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N12
cycloneive_lcell_comb \Mux52~10 (
// Equation(s):
// \Mux52~10_combout  = (\my_rf.rsel2[1]~input_o  & (\my_rf.rsel2[0]~input_o )) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & (\registerArray[5][11]~q )) # (!\my_rf.rsel2[0]~input_o  & ((\registerArray[4][11]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][11]~q ),
	.datad(\registerArray[4][11]~q ),
	.cin(gnd),
	.combout(\Mux52~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~10 .lut_mask = 16'hD9C8;
defparam \Mux52~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N13
dffeas \registerArray[6][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][11] .is_wysiwyg = "true";
defparam \registerArray[6][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N7
dffeas \registerArray[7][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][11] .is_wysiwyg = "true";
defparam \registerArray[7][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N12
cycloneive_lcell_comb \Mux52~11 (
// Equation(s):
// \Mux52~11_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux52~10_combout  & ((\registerArray[7][11]~q ))) # (!\Mux52~10_combout  & (\registerArray[6][11]~q )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux52~10_combout ))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux52~10_combout ),
	.datac(\registerArray[6][11]~q ),
	.datad(\registerArray[7][11]~q ),
	.cin(gnd),
	.combout(\Mux52~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~11 .lut_mask = 16'hEC64;
defparam \Mux52~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N0
cycloneive_lcell_comb \Mux52~19 (
// Equation(s):
// \Mux52~19_combout  = (\Mux52~16_combout  & ((\Mux52~18_combout ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux52~16_combout  & (((\my_rf.rsel2[2]~input_o  & \Mux52~11_combout ))))

	.dataa(\Mux52~18_combout ),
	.datab(\Mux52~16_combout ),
	.datac(\my_rf.rsel2[2]~input_o ),
	.datad(\Mux52~11_combout ),
	.cin(gnd),
	.combout(\Mux52~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~19 .lut_mask = 16'hBC8C;
defparam \Mux52~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N10
cycloneive_lcell_comb \Mux52~20 (
// Equation(s):
// \Mux52~20_combout  = (\my_rf.rsel2[4]~input_o  & (\Mux52~9_combout )) # (!\my_rf.rsel2[4]~input_o  & ((\Mux52~19_combout )))

	.dataa(gnd),
	.datab(\Mux52~9_combout ),
	.datac(\my_rf.rsel2[4]~input_o ),
	.datad(\Mux52~19_combout ),
	.cin(gnd),
	.combout(\Mux52~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~20 .lut_mask = 16'hCFC0;
defparam \Mux52~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X0_Y34_N1
cycloneive_io_ibuf \my_rf.wdat[12]~input (
	.i(\my_rf.wdat [12]),
	.ibar(gnd),
	.o(\my_rf.wdat[12]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[12]~input .bus_hold = "false";
defparam \my_rf.wdat[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X0_Y34_N3
dffeas \registerArray[25][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[12]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][12] .is_wysiwyg = "true";
defparam \registerArray[25][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y32_N27
dffeas \registerArray[29][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][12] .is_wysiwyg = "true";
defparam \registerArray[29][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N24
cycloneive_lcell_comb \Mux51~1 (
// Equation(s):
// \Mux51~1_combout  = (\Mux51~0_combout  & (((\registerArray[29][12]~q ) # (!\my_rf.rsel2[3]~input_o )))) # (!\Mux51~0_combout  & (\registerArray[25][12]~q  & (\my_rf.rsel2[3]~input_o )))

	.dataa(\Mux51~0_combout ),
	.datab(\registerArray[25][12]~q ),
	.datac(\my_rf.rsel2[3]~input_o ),
	.datad(\registerArray[29][12]~q ),
	.cin(gnd),
	.combout(\Mux51~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~1 .lut_mask = 16'hEA4A;
defparam \Mux51~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N15
dffeas \registerArray[28][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][12] .is_wysiwyg = "true";
defparam \registerArray[28][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y37_N29
dffeas \registerArray[20][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][12] .is_wysiwyg = "true";
defparam \registerArray[20][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N21
dffeas \registerArray[24][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][12] .is_wysiwyg = "true";
defparam \registerArray[24][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N7
dffeas \registerArray[16][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][12] .is_wysiwyg = "true";
defparam \registerArray[16][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N20
cycloneive_lcell_comb \Mux51~4 (
// Equation(s):
// \Mux51~4_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[24][12]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][12]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][12]~q ),
	.datad(\registerArray[16][12]~q ),
	.cin(gnd),
	.combout(\Mux51~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~4 .lut_mask = 16'hD9C8;
defparam \Mux51~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N28
cycloneive_lcell_comb \Mux51~5 (
// Equation(s):
// \Mux51~5_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux51~4_combout  & (\registerArray[28][12]~q )) # (!\Mux51~4_combout  & ((\registerArray[20][12]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux51~4_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[28][12]~q ),
	.datac(\registerArray[20][12]~q ),
	.datad(\Mux51~4_combout ),
	.cin(gnd),
	.combout(\Mux51~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~5 .lut_mask = 16'hDDA0;
defparam \Mux51~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N26
cycloneive_lcell_comb \Mux51~6 (
// Equation(s):
// \Mux51~6_combout  = (\my_rf.rsel2[0]~input_o  & (((\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\Mux51~3_combout )) # (!\my_rf.rsel2[1]~input_o  & ((\Mux51~5_combout )))))

	.dataa(\Mux51~3_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\my_rf.rsel2[1]~input_o ),
	.datad(\Mux51~5_combout ),
	.cin(gnd),
	.combout(\Mux51~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~6 .lut_mask = 16'hE3E0;
defparam \Mux51~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N28
cycloneive_lcell_comb \Mux51~9 (
// Equation(s):
// \Mux51~9_combout  = (\Mux51~6_combout  & ((\Mux51~8_combout ) # ((!\my_rf.rsel2[0]~input_o )))) # (!\Mux51~6_combout  & (((\Mux51~1_combout  & \my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux51~8_combout ),
	.datab(\Mux51~1_combout ),
	.datac(\Mux51~6_combout ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux51~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~9 .lut_mask = 16'hACF0;
defparam \Mux51~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y34_N17
dffeas \registerArray[11][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][12] .is_wysiwyg = "true";
defparam \registerArray[11][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N23
dffeas \registerArray[9][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][12] .is_wysiwyg = "true";
defparam \registerArray[9][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N22
cycloneive_lcell_comb \Mux51~11 (
// Equation(s):
// \Mux51~11_combout  = (\Mux51~10_combout  & ((\registerArray[11][12]~q ) # ((!\my_rf.rsel2[0]~input_o )))) # (!\Mux51~10_combout  & (((\registerArray[9][12]~q  & \my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux51~10_combout ),
	.datab(\registerArray[11][12]~q ),
	.datac(\registerArray[9][12]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux51~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~11 .lut_mask = 16'hD8AA;
defparam \Mux51~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N1
dffeas \registerArray[15][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][12] .is_wysiwyg = "true";
defparam \registerArray[15][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N31
dffeas \registerArray[14][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][12] .is_wysiwyg = "true";
defparam \registerArray[14][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N21
dffeas \registerArray[13][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][12] .is_wysiwyg = "true";
defparam \registerArray[13][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N31
dffeas \registerArray[12][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][12] .is_wysiwyg = "true";
defparam \registerArray[12][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N20
cycloneive_lcell_comb \Mux51~17 (
// Equation(s):
// \Mux51~17_combout  = (\my_rf.rsel2[1]~input_o  & (\my_rf.rsel2[0]~input_o )) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & (\registerArray[13][12]~q )) # (!\my_rf.rsel2[0]~input_o  & ((\registerArray[12][12]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[13][12]~q ),
	.datad(\registerArray[12][12]~q ),
	.cin(gnd),
	.combout(\Mux51~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~17 .lut_mask = 16'hD9C8;
defparam \Mux51~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N30
cycloneive_lcell_comb \Mux51~18 (
// Equation(s):
// \Mux51~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux51~17_combout  & (\registerArray[15][12]~q )) # (!\Mux51~17_combout  & ((\registerArray[14][12]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux51~17_combout ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[15][12]~q ),
	.datac(\registerArray[14][12]~q ),
	.datad(\Mux51~17_combout ),
	.cin(gnd),
	.combout(\Mux51~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~18 .lut_mask = 16'hDDA0;
defparam \Mux51~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N25
dffeas \registerArray[5][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][12] .is_wysiwyg = "true";
defparam \registerArray[5][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N11
dffeas \registerArray[4][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][12] .is_wysiwyg = "true";
defparam \registerArray[4][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N24
cycloneive_lcell_comb \Mux51~12 (
// Equation(s):
// \Mux51~12_combout  = (\my_rf.rsel2[1]~input_o  & (\my_rf.rsel2[0]~input_o )) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & (\registerArray[5][12]~q )) # (!\my_rf.rsel2[0]~input_o  & ((\registerArray[4][12]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][12]~q ),
	.datad(\registerArray[4][12]~q ),
	.cin(gnd),
	.combout(\Mux51~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~12 .lut_mask = 16'hD9C8;
defparam \Mux51~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N9
dffeas \registerArray[6][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][12] .is_wysiwyg = "true";
defparam \registerArray[6][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N8
cycloneive_lcell_comb \Mux51~13 (
// Equation(s):
// \Mux51~13_combout  = (\Mux51~12_combout  & ((\registerArray[7][12]~q ) # ((!\my_rf.rsel2[1]~input_o )))) # (!\Mux51~12_combout  & (((\registerArray[6][12]~q  & \my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[7][12]~q ),
	.datab(\Mux51~12_combout ),
	.datac(\registerArray[6][12]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux51~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~13 .lut_mask = 16'hB8CC;
defparam \Mux51~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N10
cycloneive_lcell_comb \Mux51~16 (
// Equation(s):
// \Mux51~16_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & ((\Mux51~13_combout ))) # (!\my_rf.rsel2[2]~input_o  & (\Mux51~15_combout ))))

	.dataa(\Mux51~15_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\my_rf.rsel2[2]~input_o ),
	.datad(\Mux51~13_combout ),
	.cin(gnd),
	.combout(\Mux51~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~16 .lut_mask = 16'hF2C2;
defparam \Mux51~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N4
cycloneive_lcell_comb \Mux51~19 (
// Equation(s):
// \Mux51~19_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux51~16_combout  & ((\Mux51~18_combout ))) # (!\Mux51~16_combout  & (\Mux51~11_combout )))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux51~16_combout ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux51~11_combout ),
	.datac(\Mux51~18_combout ),
	.datad(\Mux51~16_combout ),
	.cin(gnd),
	.combout(\Mux51~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~19 .lut_mask = 16'hF588;
defparam \Mux51~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N30
cycloneive_lcell_comb \Mux51~20 (
// Equation(s):
// \Mux51~20_combout  = (\my_rf.rsel2[4]~input_o  & (\Mux51~9_combout )) # (!\my_rf.rsel2[4]~input_o  & ((\Mux51~19_combout )))

	.dataa(\my_rf.rsel2[4]~input_o ),
	.datab(\Mux51~9_combout ),
	.datac(\Mux51~19_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux51~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~20 .lut_mask = 16'hD8D8;
defparam \Mux51~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X47_Y0_N8
cycloneive_io_ibuf \my_rf.wdat[13]~input (
	.i(\my_rf.wdat [13]),
	.ibar(gnd),
	.o(\my_rf.wdat[13]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[13]~input .bus_hold = "false";
defparam \my_rf.wdat[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X54_Y37_N15
dffeas \registerArray[4][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][13] .is_wysiwyg = "true";
defparam \registerArray[4][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N29
dffeas \registerArray[5][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][13] .is_wysiwyg = "true";
defparam \registerArray[5][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N28
cycloneive_lcell_comb \Mux50~10 (
// Equation(s):
// \Mux50~10_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & ((\registerArray[5][13]~q ))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][13]~q ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[4][13]~q ),
	.datac(\registerArray[5][13]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux50~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~10 .lut_mask = 16'hFA44;
defparam \Mux50~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N5
dffeas \registerArray[6][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][13] .is_wysiwyg = "true";
defparam \registerArray[6][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N4
cycloneive_lcell_comb \Mux50~11 (
// Equation(s):
// \Mux50~11_combout  = (\Mux50~10_combout  & ((\registerArray[7][13]~q ) # ((!\my_rf.rsel2[1]~input_o )))) # (!\Mux50~10_combout  & (((\registerArray[6][13]~q  & \my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[7][13]~q ),
	.datab(\Mux50~10_combout ),
	.datac(\registerArray[6][13]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux50~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~11 .lut_mask = 16'hB8CC;
defparam \Mux50~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y36_N9
dffeas \registerArray[13][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][13] .is_wysiwyg = "true";
defparam \registerArray[13][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y36_N27
dffeas \registerArray[12][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][13] .is_wysiwyg = "true";
defparam \registerArray[12][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y36_N8
cycloneive_lcell_comb \Mux50~17 (
// Equation(s):
// \Mux50~17_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[13][13]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[12][13]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[13][13]~q ),
	.datad(\registerArray[12][13]~q ),
	.cin(gnd),
	.combout(\Mux50~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~17 .lut_mask = 16'hB9A8;
defparam \Mux50~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N27
dffeas \registerArray[14][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][13] .is_wysiwyg = "true";
defparam \registerArray[14][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N29
dffeas \registerArray[15][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][13] .is_wysiwyg = "true";
defparam \registerArray[15][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N26
cycloneive_lcell_comb \Mux50~18 (
// Equation(s):
// \Mux50~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux50~17_combout  & ((\registerArray[15][13]~q ))) # (!\Mux50~17_combout  & (\registerArray[14][13]~q )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux50~17_combout ))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux50~17_combout ),
	.datac(\registerArray[14][13]~q ),
	.datad(\registerArray[15][13]~q ),
	.cin(gnd),
	.combout(\Mux50~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~18 .lut_mask = 16'hEC64;
defparam \Mux50~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N26
cycloneive_lcell_comb \Mux50~19 (
// Equation(s):
// \Mux50~19_combout  = (\Mux50~16_combout  & (((\Mux50~18_combout ) # (!\my_rf.rsel2[2]~input_o )))) # (!\Mux50~16_combout  & (\Mux50~11_combout  & (\my_rf.rsel2[2]~input_o )))

	.dataa(\Mux50~16_combout ),
	.datab(\Mux50~11_combout ),
	.datac(\my_rf.rsel2[2]~input_o ),
	.datad(\Mux50~18_combout ),
	.cin(gnd),
	.combout(\Mux50~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~19 .lut_mask = 16'hEA4A;
defparam \Mux50~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y33_N13
dffeas \registerArray[23][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][13] .is_wysiwyg = "true";
defparam \registerArray[23][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N17
dffeas \registerArray[27][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][13] .is_wysiwyg = "true";
defparam \registerArray[27][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N16
cycloneive_lcell_comb \Mux50~7 (
// Equation(s):
// \Mux50~7_combout  = (\my_rf.rsel2[3]~input_o  & (((\registerArray[27][13]~q ) # (\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[19][13]~q  & ((!\my_rf.rsel2[2]~input_o ))))

	.dataa(\registerArray[19][13]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][13]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux50~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~7 .lut_mask = 16'hCCE2;
defparam \Mux50~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N12
cycloneive_lcell_comb \Mux50~8 (
// Equation(s):
// \Mux50~8_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux50~7_combout  & (\registerArray[31][13]~q )) # (!\Mux50~7_combout  & ((\registerArray[23][13]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux50~7_combout ))))

	.dataa(\registerArray[31][13]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[23][13]~q ),
	.datad(\Mux50~7_combout ),
	.cin(gnd),
	.combout(\Mux50~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~8 .lut_mask = 16'hBBC0;
defparam \Mux50~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N11
dffeas \registerArray[26][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][13] .is_wysiwyg = "true";
defparam \registerArray[26][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y35_N27
dffeas \registerArray[30][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][13] .is_wysiwyg = "true";
defparam \registerArray[30][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N10
cycloneive_lcell_comb \Mux50~3 (
// Equation(s):
// \Mux50~3_combout  = (\Mux50~2_combout  & (((\registerArray[30][13]~q )) # (!\my_rf.rsel2[3]~input_o ))) # (!\Mux50~2_combout  & (\my_rf.rsel2[3]~input_o  & (\registerArray[26][13]~q )))

	.dataa(\Mux50~2_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[26][13]~q ),
	.datad(\registerArray[30][13]~q ),
	.cin(gnd),
	.combout(\Mux50~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~3 .lut_mask = 16'hEA62;
defparam \Mux50~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N22
cycloneive_lcell_comb \Mux50~6 (
// Equation(s):
// \Mux50~6_combout  = (\my_rf.rsel2[0]~input_o  & (((\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\Mux50~3_combout ))) # (!\my_rf.rsel2[1]~input_o  & (\Mux50~5_combout ))))

	.dataa(\Mux50~5_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\my_rf.rsel2[1]~input_o ),
	.datad(\Mux50~3_combout ),
	.cin(gnd),
	.combout(\Mux50~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~6 .lut_mask = 16'hF2C2;
defparam \Mux50~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N8
cycloneive_lcell_comb \Mux50~9 (
// Equation(s):
// \Mux50~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux50~6_combout  & ((\Mux50~8_combout ))) # (!\Mux50~6_combout  & (\Mux50~1_combout )))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux50~6_combout ))))

	.dataa(\Mux50~1_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux50~8_combout ),
	.datad(\Mux50~6_combout ),
	.cin(gnd),
	.combout(\Mux50~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~9 .lut_mask = 16'hF388;
defparam \Mux50~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N12
cycloneive_lcell_comb \Mux50~20 (
// Equation(s):
// \Mux50~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux50~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux50~19_combout ))

	.dataa(\Mux50~19_combout ),
	.datab(\Mux50~9_combout ),
	.datac(\my_rf.rsel2[4]~input_o ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux50~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~20 .lut_mask = 16'hCACA;
defparam \Mux50~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X0_Y32_N15
cycloneive_io_ibuf \my_rf.wdat[14]~input (
	.i(\my_rf.wdat [14]),
	.ibar(gnd),
	.o(\my_rf.wdat[14]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[14]~input .bus_hold = "false";
defparam \my_rf.wdat[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X42_Y35_N13
dffeas \registerArray[14][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][14] .is_wysiwyg = "true";
defparam \registerArray[14][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y36_N29
dffeas \registerArray[13][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][14] .is_wysiwyg = "true";
defparam \registerArray[13][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y36_N28
cycloneive_lcell_comb \Mux49~17 (
// Equation(s):
// \Mux49~17_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[13][14]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[12][14]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[12][14]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[13][14]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux49~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~17 .lut_mask = 16'hCCE2;
defparam \Mux49~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N12
cycloneive_lcell_comb \Mux49~18 (
// Equation(s):
// \Mux49~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux49~17_combout  & (\registerArray[15][14]~q )) # (!\Mux49~17_combout  & ((\registerArray[14][14]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux49~17_combout ))))

	.dataa(\registerArray[15][14]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][14]~q ),
	.datad(\Mux49~17_combout ),
	.cin(gnd),
	.combout(\Mux49~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~18 .lut_mask = 16'hBBC0;
defparam \Mux49~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y37_N17
dffeas \registerArray[9][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][14] .is_wysiwyg = "true";
defparam \registerArray[9][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y37_N19
dffeas \registerArray[11][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][14] .is_wysiwyg = "true";
defparam \registerArray[11][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y37_N16
cycloneive_lcell_comb \Mux49~11 (
// Equation(s):
// \Mux49~11_combout  = (\Mux49~10_combout  & (((\registerArray[11][14]~q )) # (!\my_rf.rsel2[0]~input_o ))) # (!\Mux49~10_combout  & (\my_rf.rsel2[0]~input_o  & (\registerArray[9][14]~q )))

	.dataa(\Mux49~10_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[9][14]~q ),
	.datad(\registerArray[11][14]~q ),
	.cin(gnd),
	.combout(\Mux49~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~11 .lut_mask = 16'hEA62;
defparam \Mux49~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N8
cycloneive_lcell_comb \Mux49~19 (
// Equation(s):
// \Mux49~19_combout  = (\Mux49~16_combout  & (((\Mux49~18_combout )) # (!\my_rf.rsel2[3]~input_o ))) # (!\Mux49~16_combout  & (\my_rf.rsel2[3]~input_o  & ((\Mux49~11_combout ))))

	.dataa(\Mux49~16_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux49~18_combout ),
	.datad(\Mux49~11_combout ),
	.cin(gnd),
	.combout(\Mux49~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~19 .lut_mask = 16'hE6A2;
defparam \Mux49~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N21
dffeas \registerArray[20][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][14] .is_wysiwyg = "true";
defparam \registerArray[20][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N25
dffeas \registerArray[24][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][14] .is_wysiwyg = "true";
defparam \registerArray[24][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N19
dffeas \registerArray[16][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][14] .is_wysiwyg = "true";
defparam \registerArray[16][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N24
cycloneive_lcell_comb \Mux49~4 (
// Equation(s):
// \Mux49~4_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[24][14]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][14]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][14]~q ),
	.datad(\registerArray[16][14]~q ),
	.cin(gnd),
	.combout(\Mux49~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~4 .lut_mask = 16'hD9C8;
defparam \Mux49~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N20
cycloneive_lcell_comb \Mux49~5 (
// Equation(s):
// \Mux49~5_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux49~4_combout  & (\registerArray[28][14]~q )) # (!\Mux49~4_combout  & ((\registerArray[20][14]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux49~4_combout ))))

	.dataa(\registerArray[28][14]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[20][14]~q ),
	.datad(\Mux49~4_combout ),
	.cin(gnd),
	.combout(\Mux49~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~5 .lut_mask = 16'hBBC0;
defparam \Mux49~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y36_N5
dffeas \registerArray[22][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][14] .is_wysiwyg = "true";
defparam \registerArray[22][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y36_N31
dffeas \registerArray[18][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][14] .is_wysiwyg = "true";
defparam \registerArray[18][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y38_N19
dffeas \registerArray[26][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][14] .is_wysiwyg = "true";
defparam \registerArray[26][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y38_N18
cycloneive_lcell_comb \Mux49~2 (
// Equation(s):
// \Mux49~2_combout  = (\my_rf.rsel2[3]~input_o  & (((\registerArray[26][14]~q ) # (\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[18][14]~q  & ((!\my_rf.rsel2[2]~input_o ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[18][14]~q ),
	.datac(\registerArray[26][14]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux49~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~2 .lut_mask = 16'hAAE4;
defparam \Mux49~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N4
cycloneive_lcell_comb \Mux49~3 (
// Equation(s):
// \Mux49~3_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux49~2_combout  & (\registerArray[30][14]~q )) # (!\Mux49~2_combout  & ((\registerArray[22][14]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux49~2_combout ))))

	.dataa(\registerArray[30][14]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][14]~q ),
	.datad(\Mux49~2_combout ),
	.cin(gnd),
	.combout(\Mux49~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~3 .lut_mask = 16'hBBC0;
defparam \Mux49~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N16
cycloneive_lcell_comb \Mux49~6 (
// Equation(s):
// \Mux49~6_combout  = (\my_rf.rsel2[0]~input_o  & (\my_rf.rsel2[1]~input_o )) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\Mux49~3_combout ))) # (!\my_rf.rsel2[1]~input_o  & (\Mux49~5_combout ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\Mux49~5_combout ),
	.datad(\Mux49~3_combout ),
	.cin(gnd),
	.combout(\Mux49~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~6 .lut_mask = 16'hDC98;
defparam \Mux49~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N21
dffeas \registerArray[27][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][14] .is_wysiwyg = "true";
defparam \registerArray[27][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N9
dffeas \registerArray[31][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][14] .is_wysiwyg = "true";
defparam \registerArray[31][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N20
cycloneive_lcell_comb \Mux49~8 (
// Equation(s):
// \Mux49~8_combout  = (\Mux49~7_combout  & (((\registerArray[31][14]~q )) # (!\my_rf.rsel2[3]~input_o ))) # (!\Mux49~7_combout  & (\my_rf.rsel2[3]~input_o  & (\registerArray[27][14]~q )))

	.dataa(\Mux49~7_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][14]~q ),
	.datad(\registerArray[31][14]~q ),
	.cin(gnd),
	.combout(\Mux49~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~8 .lut_mask = 16'hEA62;
defparam \Mux49~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N17
dffeas \registerArray[29][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][14] .is_wysiwyg = "true";
defparam \registerArray[29][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N13
dffeas \registerArray[21][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][14] .is_wysiwyg = "true";
defparam \registerArray[21][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N12
cycloneive_lcell_comb \Mux49~0 (
// Equation(s):
// \Mux49~0_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & ((\registerArray[21][14]~q ))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[17][14]~q ))))

	.dataa(\registerArray[17][14]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[21][14]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux49~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~0 .lut_mask = 16'hFC22;
defparam \Mux49~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X0_Y32_N17
dffeas \registerArray[25][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[14]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][14] .is_wysiwyg = "true";
defparam \registerArray[25][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N26
cycloneive_lcell_comb \Mux49~1 (
// Equation(s):
// \Mux49~1_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux49~0_combout  & (\registerArray[29][14]~q )) # (!\Mux49~0_combout  & ((\registerArray[25][14]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux49~0_combout ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[29][14]~q ),
	.datac(\Mux49~0_combout ),
	.datad(\registerArray[25][14]~q ),
	.cin(gnd),
	.combout(\Mux49~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~1 .lut_mask = 16'hDAD0;
defparam \Mux49~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N18
cycloneive_lcell_comb \Mux49~9 (
// Equation(s):
// \Mux49~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux49~6_combout  & (\Mux49~8_combout )) # (!\Mux49~6_combout  & ((\Mux49~1_combout ))))) # (!\my_rf.rsel2[0]~input_o  & (\Mux49~6_combout ))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\Mux49~6_combout ),
	.datac(\Mux49~8_combout ),
	.datad(\Mux49~1_combout ),
	.cin(gnd),
	.combout(\Mux49~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~9 .lut_mask = 16'hE6C4;
defparam \Mux49~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N2
cycloneive_lcell_comb \Mux49~20 (
// Equation(s):
// \Mux49~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux49~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux49~19_combout ))

	.dataa(\my_rf.rsel2[4]~input_o ),
	.datab(gnd),
	.datac(\Mux49~19_combout ),
	.datad(\Mux49~9_combout ),
	.cin(gnd),
	.combout(\Mux49~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~20 .lut_mask = 16'hFA50;
defparam \Mux49~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N15
cycloneive_io_ibuf \my_rf.wdat[15]~input (
	.i(\my_rf.wdat [15]),
	.ibar(gnd),
	.o(\my_rf.wdat[15]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[15]~input .bus_hold = "false";
defparam \my_rf.wdat[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X47_Y37_N5
dffeas \registerArray[7][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][15] .is_wysiwyg = "true";
defparam \registerArray[7][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y37_N3
dffeas \registerArray[6][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][15] .is_wysiwyg = "true";
defparam \registerArray[6][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N5
dffeas \registerArray[5][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][15] .is_wysiwyg = "true";
defparam \registerArray[5][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N4
cycloneive_lcell_comb \Mux48~10 (
// Equation(s):
// \Mux48~10_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & ((\registerArray[5][15]~q ))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][15]~q ))))

	.dataa(\registerArray[4][15]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[5][15]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux48~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~10 .lut_mask = 16'hFC22;
defparam \Mux48~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N2
cycloneive_lcell_comb \Mux48~11 (
// Equation(s):
// \Mux48~11_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux48~10_combout  & (\registerArray[7][15]~q )) # (!\Mux48~10_combout  & ((\registerArray[6][15]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux48~10_combout ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[7][15]~q ),
	.datac(\registerArray[6][15]~q ),
	.datad(\Mux48~10_combout ),
	.cin(gnd),
	.combout(\Mux48~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~11 .lut_mask = 16'hDDA0;
defparam \Mux48~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y36_N17
dffeas \registerArray[3][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][15] .is_wysiwyg = "true";
defparam \registerArray[3][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N3
dffeas \registerArray[1][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][15] .is_wysiwyg = "true";
defparam \registerArray[1][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N16
cycloneive_lcell_comb \Mux48~14 (
// Equation(s):
// \Mux48~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][15]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][15]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][15]~q ),
	.datad(\registerArray[1][15]~q ),
	.cin(gnd),
	.combout(\Mux48~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~14 .lut_mask = 16'hC480;
defparam \Mux48~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N11
dffeas \registerArray[2][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][15] .is_wysiwyg = "true";
defparam \registerArray[2][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N10
cycloneive_lcell_comb \Mux48~15 (
// Equation(s):
// \Mux48~15_combout  = (\Mux48~14_combout ) # ((!\my_rf.rsel2[0]~input_o  & (\registerArray[2][15]~q  & \my_rf.rsel2[1]~input_o )))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\Mux48~14_combout ),
	.datac(\registerArray[2][15]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux48~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~15 .lut_mask = 16'hDCCC;
defparam \Mux48~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N6
cycloneive_lcell_comb \Mux48~16 (
// Equation(s):
// \Mux48~16_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux48~13_combout ) # ((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (((!\my_rf.rsel2[2]~input_o  & \Mux48~15_combout ))))

	.dataa(\Mux48~13_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\my_rf.rsel2[2]~input_o ),
	.datad(\Mux48~15_combout ),
	.cin(gnd),
	.combout(\Mux48~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~16 .lut_mask = 16'hCBC8;
defparam \Mux48~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N24
cycloneive_lcell_comb \Mux48~19 (
// Equation(s):
// \Mux48~19_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux48~16_combout  & (\Mux48~18_combout )) # (!\Mux48~16_combout  & ((\Mux48~11_combout ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux48~16_combout ))))

	.dataa(\Mux48~18_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\Mux48~11_combout ),
	.datad(\Mux48~16_combout ),
	.cin(gnd),
	.combout(\Mux48~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~19 .lut_mask = 16'hBBC0;
defparam \Mux48~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y35_N23
dffeas \registerArray[20][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][15] .is_wysiwyg = "true";
defparam \registerArray[20][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N23
dffeas \registerArray[16][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][15] .is_wysiwyg = "true";
defparam \registerArray[16][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N22
cycloneive_lcell_comb \Mux48~4 (
// Equation(s):
// \Mux48~4_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[20][15]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][15]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[20][15]~q ),
	.datad(\registerArray[16][15]~q ),
	.cin(gnd),
	.combout(\Mux48~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~4 .lut_mask = 16'hB9A8;
defparam \Mux48~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N3
dffeas \registerArray[24][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][15] .is_wysiwyg = "true";
defparam \registerArray[24][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N2
cycloneive_lcell_comb \Mux48~5 (
// Equation(s):
// \Mux48~5_combout  = (\Mux48~4_combout  & ((\registerArray[28][15]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux48~4_combout  & (((\registerArray[24][15]~q  & \my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[28][15]~q ),
	.datab(\Mux48~4_combout ),
	.datac(\registerArray[24][15]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux48~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~5 .lut_mask = 16'hB8CC;
defparam \Mux48~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y35_N29
dffeas \registerArray[30][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][15] .is_wysiwyg = "true";
defparam \registerArray[30][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y34_N25
dffeas \registerArray[26][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][15] .is_wysiwyg = "true";
defparam \registerArray[26][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N24
cycloneive_lcell_comb \Mux48~3 (
// Equation(s):
// \Mux48~3_combout  = (\Mux48~2_combout  & ((\registerArray[30][15]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux48~2_combout  & (((\registerArray[26][15]~q  & \my_rf.rsel2[3]~input_o ))))

	.dataa(\Mux48~2_combout ),
	.datab(\registerArray[30][15]~q ),
	.datac(\registerArray[26][15]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux48~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~3 .lut_mask = 16'hD8AA;
defparam \Mux48~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N4
cycloneive_lcell_comb \Mux48~6 (
// Equation(s):
// \Mux48~6_combout  = (\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o ) # ((\Mux48~3_combout )))) # (!\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & (\Mux48~5_combout )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux48~5_combout ),
	.datad(\Mux48~3_combout ),
	.cin(gnd),
	.combout(\Mux48~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~6 .lut_mask = 16'hBA98;
defparam \Mux48~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N17
dffeas \registerArray[27][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][15] .is_wysiwyg = "true";
defparam \registerArray[27][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N19
dffeas \registerArray[19][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][15] .is_wysiwyg = "true";
defparam \registerArray[19][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N16
cycloneive_lcell_comb \Mux48~7 (
// Equation(s):
// \Mux48~7_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[27][15]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[19][15]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][15]~q ),
	.datad(\registerArray[19][15]~q ),
	.cin(gnd),
	.combout(\Mux48~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~7 .lut_mask = 16'hD9C8;
defparam \Mux48~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y33_N1
dffeas \registerArray[23][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][15] .is_wysiwyg = "true";
defparam \registerArray[23][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N0
cycloneive_lcell_comb \Mux48~8 (
// Equation(s):
// \Mux48~8_combout  = (\Mux48~7_combout  & ((\registerArray[31][15]~q ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux48~7_combout  & (((\registerArray[23][15]~q  & \my_rf.rsel2[2]~input_o ))))

	.dataa(\registerArray[31][15]~q ),
	.datab(\Mux48~7_combout ),
	.datac(\registerArray[23][15]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux48~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~8 .lut_mask = 16'hB8CC;
defparam \Mux48~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N17
dffeas \registerArray[29][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][15] .is_wysiwyg = "true";
defparam \registerArray[29][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N1
dffeas \registerArray[17][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][15] .is_wysiwyg = "true";
defparam \registerArray[17][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y34_N15
dffeas \registerArray[25][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][15] .is_wysiwyg = "true";
defparam \registerArray[25][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N14
cycloneive_lcell_comb \Mux48~0 (
// Equation(s):
// \Mux48~0_combout  = (\my_rf.rsel2[3]~input_o  & (((\registerArray[25][15]~q ) # (\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[17][15]~q  & ((!\my_rf.rsel2[2]~input_o ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[17][15]~q ),
	.datac(\registerArray[25][15]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux48~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~0 .lut_mask = 16'hAAE4;
defparam \Mux48~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y0_N17
dffeas \registerArray[21][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[15]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][15] .is_wysiwyg = "true";
defparam \registerArray[21][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N4
cycloneive_lcell_comb \Mux48~1 (
// Equation(s):
// \Mux48~1_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux48~0_combout  & (\registerArray[29][15]~q )) # (!\Mux48~0_combout  & ((\registerArray[21][15]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux48~0_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[29][15]~q ),
	.datac(\Mux48~0_combout ),
	.datad(\registerArray[21][15]~q ),
	.cin(gnd),
	.combout(\Mux48~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~1 .lut_mask = 16'hDAD0;
defparam \Mux48~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N8
cycloneive_lcell_comb \Mux48~9 (
// Equation(s):
// \Mux48~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux48~6_combout  & (\Mux48~8_combout )) # (!\Mux48~6_combout  & ((\Mux48~1_combout ))))) # (!\my_rf.rsel2[0]~input_o  & (\Mux48~6_combout ))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\Mux48~6_combout ),
	.datac(\Mux48~8_combout ),
	.datad(\Mux48~1_combout ),
	.cin(gnd),
	.combout(\Mux48~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~9 .lut_mask = 16'hE6C4;
defparam \Mux48~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N26
cycloneive_lcell_comb \Mux48~20 (
// Equation(s):
// \Mux48~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux48~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux48~19_combout ))

	.dataa(gnd),
	.datab(\Mux48~19_combout ),
	.datac(\Mux48~9_combout ),
	.datad(\my_rf.rsel2[4]~input_o ),
	.cin(gnd),
	.combout(\Mux48~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~20 .lut_mask = 16'hF0CC;
defparam \Mux48~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X0_Y35_N1
cycloneive_io_ibuf \my_rf.wdat[16]~input (
	.i(\my_rf.wdat [16]),
	.ibar(gnd),
	.o(\my_rf.wdat[16]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[16]~input .bus_hold = "false";
defparam \my_rf.wdat[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X43_Y39_N15
dffeas \registerArray[11][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][16] .is_wysiwyg = "true";
defparam \registerArray[11][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y39_N5
dffeas \registerArray[9][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][16] .is_wysiwyg = "true";
defparam \registerArray[9][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N4
cycloneive_lcell_comb \Mux47~11 (
// Equation(s):
// \Mux47~11_combout  = (\Mux47~10_combout  & ((\registerArray[11][16]~q ) # ((!\my_rf.rsel2[0]~input_o )))) # (!\Mux47~10_combout  & (((\registerArray[9][16]~q  & \my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux47~10_combout ),
	.datab(\registerArray[11][16]~q ),
	.datac(\registerArray[9][16]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux47~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~11 .lut_mask = 16'hD8AA;
defparam \Mux47~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y36_N9
dffeas \registerArray[14][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][16] .is_wysiwyg = "true";
defparam \registerArray[14][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y36_N3
dffeas \registerArray[15][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][16] .is_wysiwyg = "true";
defparam \registerArray[15][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N8
cycloneive_lcell_comb \Mux47~18 (
// Equation(s):
// \Mux47~18_combout  = (\Mux47~17_combout  & (((\registerArray[15][16]~q )) # (!\my_rf.rsel2[1]~input_o ))) # (!\Mux47~17_combout  & (\my_rf.rsel2[1]~input_o  & (\registerArray[14][16]~q )))

	.dataa(\Mux47~17_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][16]~q ),
	.datad(\registerArray[15][16]~q ),
	.cin(gnd),
	.combout(\Mux47~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~18 .lut_mask = 16'hEA62;
defparam \Mux47~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N20
cycloneive_lcell_comb \Mux47~19 (
// Equation(s):
// \Mux47~19_combout  = (\Mux47~16_combout  & (((\Mux47~18_combout ) # (!\my_rf.rsel2[3]~input_o )))) # (!\Mux47~16_combout  & (\Mux47~11_combout  & ((\my_rf.rsel2[3]~input_o ))))

	.dataa(\Mux47~16_combout ),
	.datab(\Mux47~11_combout ),
	.datac(\Mux47~18_combout ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux47~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~19 .lut_mask = 16'hE4AA;
defparam \Mux47~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X0_Y35_N3
dffeas \registerArray[25][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[16]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][16] .is_wysiwyg = "true";
defparam \registerArray[25][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N3
dffeas \registerArray[21][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][16] .is_wysiwyg = "true";
defparam \registerArray[21][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N29
dffeas \registerArray[17][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][16] .is_wysiwyg = "true";
defparam \registerArray[17][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N2
cycloneive_lcell_comb \Mux47~0 (
// Equation(s):
// \Mux47~0_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[21][16]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[17][16]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[21][16]~q ),
	.datad(\registerArray[17][16]~q ),
	.cin(gnd),
	.combout(\Mux47~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~0 .lut_mask = 16'hB9A8;
defparam \Mux47~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N0
cycloneive_lcell_comb \Mux47~1 (
// Equation(s):
// \Mux47~1_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux47~0_combout  & (\registerArray[29][16]~q )) # (!\Mux47~0_combout  & ((\registerArray[25][16]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux47~0_combout ))))

	.dataa(\registerArray[29][16]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[25][16]~q ),
	.datad(\Mux47~0_combout ),
	.cin(gnd),
	.combout(\Mux47~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~1 .lut_mask = 16'hBBC0;
defparam \Mux47~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y38_N31
dffeas \registerArray[22][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][16] .is_wysiwyg = "true";
defparam \registerArray[22][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y35_N31
dffeas \registerArray[30][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][16] .is_wysiwyg = "true";
defparam \registerArray[30][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N30
cycloneive_lcell_comb \Mux47~3 (
// Equation(s):
// \Mux47~3_combout  = (\Mux47~2_combout  & (((\registerArray[30][16]~q )) # (!\my_rf.rsel2[2]~input_o ))) # (!\Mux47~2_combout  & (\my_rf.rsel2[2]~input_o  & (\registerArray[22][16]~q )))

	.dataa(\Mux47~2_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[22][16]~q ),
	.datad(\registerArray[30][16]~q ),
	.cin(gnd),
	.combout(\Mux47~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~3 .lut_mask = 16'hEA62;
defparam \Mux47~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N18
cycloneive_lcell_comb \Mux47~6 (
// Equation(s):
// \Mux47~6_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o ) # (\Mux47~3_combout )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux47~5_combout  & (!\my_rf.rsel2[0]~input_o )))

	.dataa(\Mux47~5_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux47~3_combout ),
	.cin(gnd),
	.combout(\Mux47~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~6 .lut_mask = 16'hCEC2;
defparam \Mux47~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N4
cycloneive_lcell_comb \Mux47~9 (
// Equation(s):
// \Mux47~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux47~6_combout  & (\Mux47~8_combout )) # (!\Mux47~6_combout  & ((\Mux47~1_combout ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux47~6_combout ))))

	.dataa(\Mux47~8_combout ),
	.datab(\Mux47~1_combout ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux47~6_combout ),
	.cin(gnd),
	.combout(\Mux47~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~9 .lut_mask = 16'hAFC0;
defparam \Mux47~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N6
cycloneive_lcell_comb \Mux47~20 (
// Equation(s):
// \Mux47~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux47~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux47~19_combout ))

	.dataa(gnd),
	.datab(\Mux47~19_combout ),
	.datac(\Mux47~9_combout ),
	.datad(\my_rf.rsel2[4]~input_o ),
	.cin(gnd),
	.combout(\Mux47~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~20 .lut_mask = 16'hF0CC;
defparam \Mux47~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X45_Y0_N15
cycloneive_io_ibuf \my_rf.wdat[17]~input (
	.i(\my_rf.wdat [17]),
	.ibar(gnd),
	.o(\my_rf.wdat[17]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[17]~input .bus_hold = "false";
defparam \my_rf.wdat[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X47_Y37_N19
dffeas \registerArray[7][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][17] .is_wysiwyg = "true";
defparam \registerArray[7][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y37_N17
dffeas \registerArray[6][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][17] .is_wysiwyg = "true";
defparam \registerArray[6][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N16
cycloneive_lcell_comb \Mux46~11 (
// Equation(s):
// \Mux46~11_combout  = (\Mux46~10_combout  & ((\registerArray[7][17]~q ) # ((!\my_rf.rsel2[1]~input_o )))) # (!\Mux46~10_combout  & (((\registerArray[6][17]~q  & \my_rf.rsel2[1]~input_o ))))

	.dataa(\Mux46~10_combout ),
	.datab(\registerArray[7][17]~q ),
	.datac(\registerArray[6][17]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux46~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~11 .lut_mask = 16'hD8AA;
defparam \Mux46~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y36_N11
dffeas \registerArray[14][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][17] .is_wysiwyg = "true";
defparam \registerArray[14][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y36_N29
dffeas \registerArray[15][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][17] .is_wysiwyg = "true";
defparam \registerArray[15][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N10
cycloneive_lcell_comb \Mux46~18 (
// Equation(s):
// \Mux46~18_combout  = (\Mux46~17_combout  & (((\registerArray[15][17]~q )) # (!\my_rf.rsel2[1]~input_o ))) # (!\Mux46~17_combout  & (\my_rf.rsel2[1]~input_o  & (\registerArray[14][17]~q )))

	.dataa(\Mux46~17_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][17]~q ),
	.datad(\registerArray[15][17]~q ),
	.cin(gnd),
	.combout(\Mux46~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~18 .lut_mask = 16'hEA62;
defparam \Mux46~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N14
cycloneive_lcell_comb \Mux46~19 (
// Equation(s):
// \Mux46~19_combout  = (\Mux46~16_combout  & (((\Mux46~18_combout ) # (!\my_rf.rsel2[2]~input_o )))) # (!\Mux46~16_combout  & (\Mux46~11_combout  & ((\my_rf.rsel2[2]~input_o ))))

	.dataa(\Mux46~16_combout ),
	.datab(\Mux46~11_combout ),
	.datac(\Mux46~18_combout ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux46~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~19 .lut_mask = 16'hE4AA;
defparam \Mux46~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y0_N17
dffeas \registerArray[21][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[17]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][17] .is_wysiwyg = "true";
defparam \registerArray[21][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y32_N25
dffeas \registerArray[29][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][17] .is_wysiwyg = "true";
defparam \registerArray[29][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N10
cycloneive_lcell_comb \Mux46~1 (
// Equation(s):
// \Mux46~1_combout  = (\Mux46~0_combout  & (((\registerArray[29][17]~q ) # (!\my_rf.rsel2[2]~input_o )))) # (!\Mux46~0_combout  & (\registerArray[21][17]~q  & (\my_rf.rsel2[2]~input_o )))

	.dataa(\Mux46~0_combout ),
	.datab(\registerArray[21][17]~q ),
	.datac(\my_rf.rsel2[2]~input_o ),
	.datad(\registerArray[29][17]~q ),
	.cin(gnd),
	.combout(\Mux46~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~1 .lut_mask = 16'hEA4A;
defparam \Mux46~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y35_N25
dffeas \registerArray[26][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][17] .is_wysiwyg = "true";
defparam \registerArray[26][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y37_N3
dffeas \registerArray[18][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][17] .is_wysiwyg = "true";
defparam \registerArray[18][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y37_N17
dffeas \registerArray[22][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][17] .is_wysiwyg = "true";
defparam \registerArray[22][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N16
cycloneive_lcell_comb \Mux46~2 (
// Equation(s):
// \Mux46~2_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[22][17]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[18][17]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[18][17]~q ),
	.datac(\registerArray[22][17]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux46~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~2 .lut_mask = 16'hAAE4;
defparam \Mux46~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N24
cycloneive_lcell_comb \Mux46~3 (
// Equation(s):
// \Mux46~3_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux46~2_combout  & (\registerArray[30][17]~q )) # (!\Mux46~2_combout  & ((\registerArray[26][17]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux46~2_combout ))))

	.dataa(\registerArray[30][17]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[26][17]~q ),
	.datad(\Mux46~2_combout ),
	.cin(gnd),
	.combout(\Mux46~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~3 .lut_mask = 16'hBBC0;
defparam \Mux46~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N10
cycloneive_lcell_comb \Mux46~6 (
// Equation(s):
// \Mux46~6_combout  = (\my_rf.rsel2[0]~input_o  & (((\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\Mux46~3_combout ))) # (!\my_rf.rsel2[1]~input_o  & (\Mux46~5_combout ))))

	.dataa(\Mux46~5_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\my_rf.rsel2[1]~input_o ),
	.datad(\Mux46~3_combout ),
	.cin(gnd),
	.combout(\Mux46~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~6 .lut_mask = 16'hF2C2;
defparam \Mux46~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N20
cycloneive_lcell_comb \Mux46~9 (
// Equation(s):
// \Mux46~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux46~6_combout  & (\Mux46~8_combout )) # (!\Mux46~6_combout  & ((\Mux46~1_combout ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux46~6_combout ))))

	.dataa(\Mux46~8_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux46~1_combout ),
	.datad(\Mux46~6_combout ),
	.cin(gnd),
	.combout(\Mux46~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~9 .lut_mask = 16'hBBC0;
defparam \Mux46~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N24
cycloneive_lcell_comb \Mux46~20 (
// Equation(s):
// \Mux46~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux46~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux46~19_combout ))

	.dataa(gnd),
	.datab(\Mux46~19_combout ),
	.datac(\Mux46~9_combout ),
	.datad(\my_rf.rsel2[4]~input_o ),
	.cin(gnd),
	.combout(\Mux46~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~20 .lut_mask = 16'hF0CC;
defparam \Mux46~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X45_Y0_N22
cycloneive_io_ibuf \my_rf.wdat[18]~input (
	.i(\my_rf.wdat [18]),
	.ibar(gnd),
	.o(\my_rf.wdat[18]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[18]~input .bus_hold = "false";
defparam \my_rf.wdat[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X49_Y29_N21
dffeas \registerArray[6][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][18] .is_wysiwyg = "true";
defparam \registerArray[6][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y29_N29
dffeas \registerArray[5][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][18] .is_wysiwyg = "true";
defparam \registerArray[5][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N28
cycloneive_lcell_comb \Mux45~12 (
// Equation(s):
// \Mux45~12_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[5][18]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][18]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[4][18]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][18]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux45~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~12 .lut_mask = 16'hCCE2;
defparam \Mux45~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N20
cycloneive_lcell_comb \Mux45~13 (
// Equation(s):
// \Mux45~13_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux45~12_combout  & (\registerArray[7][18]~q )) # (!\Mux45~12_combout  & ((\registerArray[6][18]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux45~12_combout ))))

	.dataa(\registerArray[7][18]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[6][18]~q ),
	.datad(\Mux45~12_combout ),
	.cin(gnd),
	.combout(\Mux45~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~13 .lut_mask = 16'hBBC0;
defparam \Mux45~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N29
dffeas \registerArray[2][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][18] .is_wysiwyg = "true";
defparam \registerArray[2][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N17
dffeas \registerArray[3][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][18] .is_wysiwyg = "true";
defparam \registerArray[3][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N19
dffeas \registerArray[1][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][18] .is_wysiwyg = "true";
defparam \registerArray[1][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N16
cycloneive_lcell_comb \Mux45~14 (
// Equation(s):
// \Mux45~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][18]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][18]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][18]~q ),
	.datad(\registerArray[1][18]~q ),
	.cin(gnd),
	.combout(\Mux45~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~14 .lut_mask = 16'hC480;
defparam \Mux45~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N28
cycloneive_lcell_comb \Mux45~15 (
// Equation(s):
// \Mux45~15_combout  = (\Mux45~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][18]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][18]~q ),
	.datad(\Mux45~14_combout ),
	.cin(gnd),
	.combout(\Mux45~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~15 .lut_mask = 16'hFF20;
defparam \Mux45~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N0
cycloneive_lcell_comb \Mux45~16 (
// Equation(s):
// \Mux45~16_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\Mux45~13_combout )) # (!\my_rf.rsel2[2]~input_o  & ((\Mux45~15_combout )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux45~13_combout ),
	.datac(\my_rf.rsel2[2]~input_o ),
	.datad(\Mux45~15_combout ),
	.cin(gnd),
	.combout(\Mux45~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~16 .lut_mask = 16'hE5E0;
defparam \Mux45~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N17
dffeas \registerArray[13][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][18] .is_wysiwyg = "true";
defparam \registerArray[13][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y36_N19
dffeas \registerArray[12][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][18] .is_wysiwyg = "true";
defparam \registerArray[12][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N16
cycloneive_lcell_comb \Mux45~17 (
// Equation(s):
// \Mux45~17_combout  = (\my_rf.rsel2[1]~input_o  & (\my_rf.rsel2[0]~input_o )) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & (\registerArray[13][18]~q )) # (!\my_rf.rsel2[0]~input_o  & ((\registerArray[12][18]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[13][18]~q ),
	.datad(\registerArray[12][18]~q ),
	.cin(gnd),
	.combout(\Mux45~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~17 .lut_mask = 16'hD9C8;
defparam \Mux45~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N21
dffeas \registerArray[14][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][18] .is_wysiwyg = "true";
defparam \registerArray[14][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N7
dffeas \registerArray[15][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][18] .is_wysiwyg = "true";
defparam \registerArray[15][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N20
cycloneive_lcell_comb \Mux45~18 (
// Equation(s):
// \Mux45~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux45~17_combout  & ((\registerArray[15][18]~q ))) # (!\Mux45~17_combout  & (\registerArray[14][18]~q )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux45~17_combout ))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux45~17_combout ),
	.datac(\registerArray[14][18]~q ),
	.datad(\registerArray[15][18]~q ),
	.cin(gnd),
	.combout(\Mux45~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~18 .lut_mask = 16'hEC64;
defparam \Mux45~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y31_N9
dffeas \registerArray[9][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][18] .is_wysiwyg = "true";
defparam \registerArray[9][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y31_N19
dffeas \registerArray[11][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][18] .is_wysiwyg = "true";
defparam \registerArray[11][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N8
cycloneive_lcell_comb \Mux45~11 (
// Equation(s):
// \Mux45~11_combout  = (\Mux45~10_combout  & (((\registerArray[11][18]~q )) # (!\my_rf.rsel2[0]~input_o ))) # (!\Mux45~10_combout  & (\my_rf.rsel2[0]~input_o  & (\registerArray[9][18]~q )))

	.dataa(\Mux45~10_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[9][18]~q ),
	.datad(\registerArray[11][18]~q ),
	.cin(gnd),
	.combout(\Mux45~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~11 .lut_mask = 16'hEA62;
defparam \Mux45~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y30_N10
cycloneive_lcell_comb \Mux45~19 (
// Equation(s):
// \Mux45~19_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux45~16_combout  & (\Mux45~18_combout )) # (!\Mux45~16_combout  & ((\Mux45~11_combout ))))) # (!\my_rf.rsel2[3]~input_o  & (\Mux45~16_combout ))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux45~16_combout ),
	.datac(\Mux45~18_combout ),
	.datad(\Mux45~11_combout ),
	.cin(gnd),
	.combout(\Mux45~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~19 .lut_mask = 16'hE6C4;
defparam \Mux45~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N29
dffeas \registerArray[29][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][18] .is_wysiwyg = "true";
defparam \registerArray[29][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N7
dffeas \registerArray[21][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][18] .is_wysiwyg = "true";
defparam \registerArray[21][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N25
dffeas \registerArray[17][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][18] .is_wysiwyg = "true";
defparam \registerArray[17][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N6
cycloneive_lcell_comb \Mux45~0 (
// Equation(s):
// \Mux45~0_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[21][18]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[17][18]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[21][18]~q ),
	.datad(\registerArray[17][18]~q ),
	.cin(gnd),
	.combout(\Mux45~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~0 .lut_mask = 16'hB9A8;
defparam \Mux45~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y0_N24
dffeas \registerArray[25][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[18]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][18] .is_wysiwyg = "true";
defparam \registerArray[25][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N24
cycloneive_lcell_comb \Mux45~1 (
// Equation(s):
// \Mux45~1_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux45~0_combout  & (\registerArray[29][18]~q )) # (!\Mux45~0_combout  & ((\registerArray[25][18]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux45~0_combout ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[29][18]~q ),
	.datac(\Mux45~0_combout ),
	.datad(\registerArray[25][18]~q ),
	.cin(gnd),
	.combout(\Mux45~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~1 .lut_mask = 16'hDAD0;
defparam \Mux45~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y32_N19
dffeas \registerArray[20][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][18] .is_wysiwyg = "true";
defparam \registerArray[20][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y32_N21
dffeas \registerArray[28][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][18] .is_wysiwyg = "true";
defparam \registerArray[28][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N18
cycloneive_lcell_comb \Mux45~5 (
// Equation(s):
// \Mux45~5_combout  = (\Mux45~4_combout  & (((\registerArray[28][18]~q )) # (!\my_rf.rsel2[2]~input_o ))) # (!\Mux45~4_combout  & (\my_rf.rsel2[2]~input_o  & (\registerArray[20][18]~q )))

	.dataa(\Mux45~4_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[20][18]~q ),
	.datad(\registerArray[28][18]~q ),
	.cin(gnd),
	.combout(\Mux45~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~5 .lut_mask = 16'hEA62;
defparam \Mux45~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y38_N27
dffeas \registerArray[26][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][18] .is_wysiwyg = "true";
defparam \registerArray[26][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y38_N29
dffeas \registerArray[18][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][18] .is_wysiwyg = "true";
defparam \registerArray[18][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N26
cycloneive_lcell_comb \Mux45~2 (
// Equation(s):
// \Mux45~2_combout  = (\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o ) # ((\registerArray[26][18]~q )))) # (!\my_rf.rsel2[3]~input_o  & (!\my_rf.rsel2[2]~input_o  & ((\registerArray[18][18]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[26][18]~q ),
	.datad(\registerArray[18][18]~q ),
	.cin(gnd),
	.combout(\Mux45~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~2 .lut_mask = 16'hB9A8;
defparam \Mux45~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y37_N21
dffeas \registerArray[22][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][18] .is_wysiwyg = "true";
defparam \registerArray[22][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y37_N31
dffeas \registerArray[30][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][18] .is_wysiwyg = "true";
defparam \registerArray[30][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N20
cycloneive_lcell_comb \Mux45~3 (
// Equation(s):
// \Mux45~3_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux45~2_combout  & ((\registerArray[30][18]~q ))) # (!\Mux45~2_combout  & (\registerArray[22][18]~q )))) # (!\my_rf.rsel2[2]~input_o  & (\Mux45~2_combout ))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux45~2_combout ),
	.datac(\registerArray[22][18]~q ),
	.datad(\registerArray[30][18]~q ),
	.cin(gnd),
	.combout(\Mux45~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~3 .lut_mask = 16'hEC64;
defparam \Mux45~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N22
cycloneive_lcell_comb \Mux45~6 (
// Equation(s):
// \Mux45~6_combout  = (\my_rf.rsel2[1]~input_o  & (((\Mux45~3_combout ) # (\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux45~5_combout  & ((!\my_rf.rsel2[0]~input_o ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux45~5_combout ),
	.datac(\Mux45~3_combout ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux45~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~6 .lut_mask = 16'hAAE4;
defparam \Mux45~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y28_N9
dffeas \registerArray[19][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][18] .is_wysiwyg = "true";
defparam \registerArray[19][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N15
dffeas \registerArray[23][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][18] .is_wysiwyg = "true";
defparam \registerArray[23][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N14
cycloneive_lcell_comb \Mux45~7 (
// Equation(s):
// \Mux45~7_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & ((\registerArray[23][18]~q ))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[19][18]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\registerArray[19][18]~q ),
	.datac(\registerArray[23][18]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux45~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~7 .lut_mask = 16'hFA44;
defparam \Mux45~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y32_N13
dffeas \registerArray[27][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][18] .is_wysiwyg = "true";
defparam \registerArray[27][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N12
cycloneive_lcell_comb \Mux45~8 (
// Equation(s):
// \Mux45~8_combout  = (\Mux45~7_combout  & ((\registerArray[31][18]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux45~7_combout  & (((\registerArray[27][18]~q  & \my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[31][18]~q ),
	.datab(\Mux45~7_combout ),
	.datac(\registerArray[27][18]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux45~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~8 .lut_mask = 16'hB8CC;
defparam \Mux45~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N16
cycloneive_lcell_comb \Mux45~9 (
// Equation(s):
// \Mux45~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux45~6_combout  & ((\Mux45~8_combout ))) # (!\Mux45~6_combout  & (\Mux45~1_combout )))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux45~6_combout ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\Mux45~1_combout ),
	.datac(\Mux45~6_combout ),
	.datad(\Mux45~8_combout ),
	.cin(gnd),
	.combout(\Mux45~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~9 .lut_mask = 16'hF858;
defparam \Mux45~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N2
cycloneive_lcell_comb \Mux45~20 (
// Equation(s):
// \Mux45~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux45~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux45~19_combout ))

	.dataa(\my_rf.rsel2[4]~input_o ),
	.datab(gnd),
	.datac(\Mux45~19_combout ),
	.datad(\Mux45~9_combout ),
	.cin(gnd),
	.combout(\Mux45~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~20 .lut_mask = 16'hFA50;
defparam \Mux45~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N8
cycloneive_io_ibuf \my_rf.wdat[19]~input (
	.i(\my_rf.wdat [19]),
	.ibar(gnd),
	.o(\my_rf.wdat[19]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[19]~input .bus_hold = "false";
defparam \my_rf.wdat[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X52_Y34_N13
dffeas \registerArray[9][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][19] .is_wysiwyg = "true";
defparam \registerArray[9][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y31_N21
dffeas \registerArray[10][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][19] .is_wysiwyg = "true";
defparam \registerArray[10][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N20
cycloneive_lcell_comb \Mux44~12 (
// Equation(s):
// \Mux44~12_combout  = (\my_rf.rsel2[0]~input_o  & (((\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[10][19]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[8][19]~q ))))

	.dataa(\registerArray[8][19]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[10][19]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux44~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~12 .lut_mask = 16'hFC22;
defparam \Mux44~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N12
cycloneive_lcell_comb \Mux44~13 (
// Equation(s):
// \Mux44~13_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux44~12_combout  & (\registerArray[11][19]~q )) # (!\Mux44~12_combout  & ((\registerArray[9][19]~q ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux44~12_combout ))))

	.dataa(\registerArray[11][19]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[9][19]~q ),
	.datad(\Mux44~12_combout ),
	.cin(gnd),
	.combout(\Mux44~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~13 .lut_mask = 16'hBBC0;
defparam \Mux44~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N3
dffeas \registerArray[2][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][19] .is_wysiwyg = "true";
defparam \registerArray[2][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N21
dffeas \registerArray[3][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][19] .is_wysiwyg = "true";
defparam \registerArray[3][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N20
cycloneive_lcell_comb \Mux44~14 (
// Equation(s):
// \Mux44~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[3][19]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[1][19]~q ))))

	.dataa(\registerArray[1][19]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][19]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux44~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~14 .lut_mask = 16'hC088;
defparam \Mux44~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N2
cycloneive_lcell_comb \Mux44~15 (
// Equation(s):
// \Mux44~15_combout  = (\Mux44~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][19]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][19]~q ),
	.datad(\Mux44~14_combout ),
	.cin(gnd),
	.combout(\Mux44~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~15 .lut_mask = 16'hFF20;
defparam \Mux44~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N8
cycloneive_lcell_comb \Mux44~16 (
// Equation(s):
// \Mux44~16_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\Mux44~13_combout )) # (!\my_rf.rsel2[3]~input_o  & ((\Mux44~15_combout )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux44~13_combout ),
	.datac(\my_rf.rsel2[3]~input_o ),
	.datad(\Mux44~15_combout ),
	.cin(gnd),
	.combout(\Mux44~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~16 .lut_mask = 16'hE5E0;
defparam \Mux44~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N25
dffeas \registerArray[15][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][19] .is_wysiwyg = "true";
defparam \registerArray[15][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N23
dffeas \registerArray[14][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][19] .is_wysiwyg = "true";
defparam \registerArray[14][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N23
dffeas \registerArray[13][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][19] .is_wysiwyg = "true";
defparam \registerArray[13][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N17
dffeas \registerArray[12][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][19] .is_wysiwyg = "true";
defparam \registerArray[12][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N22
cycloneive_lcell_comb \Mux44~17 (
// Equation(s):
// \Mux44~17_combout  = (\my_rf.rsel2[1]~input_o  & (\my_rf.rsel2[0]~input_o )) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & (\registerArray[13][19]~q )) # (!\my_rf.rsel2[0]~input_o  & ((\registerArray[12][19]~q )))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[13][19]~q ),
	.datad(\registerArray[12][19]~q ),
	.cin(gnd),
	.combout(\Mux44~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~17 .lut_mask = 16'hD9C8;
defparam \Mux44~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N22
cycloneive_lcell_comb \Mux44~18 (
// Equation(s):
// \Mux44~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux44~17_combout  & (\registerArray[15][19]~q )) # (!\Mux44~17_combout  & ((\registerArray[14][19]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux44~17_combout ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[15][19]~q ),
	.datac(\registerArray[14][19]~q ),
	.datad(\Mux44~17_combout ),
	.cin(gnd),
	.combout(\Mux44~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~18 .lut_mask = 16'hDDA0;
defparam \Mux44~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N15
dffeas \registerArray[7][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][19] .is_wysiwyg = "true";
defparam \registerArray[7][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N21
dffeas \registerArray[6][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][19] .is_wysiwyg = "true";
defparam \registerArray[6][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N17
dffeas \registerArray[5][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][19] .is_wysiwyg = "true";
defparam \registerArray[5][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N16
cycloneive_lcell_comb \Mux44~10 (
// Equation(s):
// \Mux44~10_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[5][19]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][19]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[4][19]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[5][19]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux44~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~10 .lut_mask = 16'hCCE2;
defparam \Mux44~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N20
cycloneive_lcell_comb \Mux44~11 (
// Equation(s):
// \Mux44~11_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux44~10_combout  & (\registerArray[7][19]~q )) # (!\Mux44~10_combout  & ((\registerArray[6][19]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux44~10_combout ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[7][19]~q ),
	.datac(\registerArray[6][19]~q ),
	.datad(\Mux44~10_combout ),
	.cin(gnd),
	.combout(\Mux44~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~11 .lut_mask = 16'hDDA0;
defparam \Mux44~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N18
cycloneive_lcell_comb \Mux44~19 (
// Equation(s):
// \Mux44~19_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux44~16_combout  & (\Mux44~18_combout )) # (!\Mux44~16_combout  & ((\Mux44~11_combout ))))) # (!\my_rf.rsel2[2]~input_o  & (\Mux44~16_combout ))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux44~16_combout ),
	.datac(\Mux44~18_combout ),
	.datad(\Mux44~11_combout ),
	.cin(gnd),
	.combout(\Mux44~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~19 .lut_mask = 16'hE6C4;
defparam \Mux44~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y32_N17
dffeas \registerArray[31][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][19] .is_wysiwyg = "true";
defparam \registerArray[31][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y32_N13
dffeas \registerArray[23][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][19] .is_wysiwyg = "true";
defparam \registerArray[23][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N12
cycloneive_lcell_comb \Mux44~8 (
// Equation(s):
// \Mux44~8_combout  = (\Mux44~7_combout  & ((\registerArray[31][19]~q ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux44~7_combout  & (((\registerArray[23][19]~q  & \my_rf.rsel2[2]~input_o ))))

	.dataa(\Mux44~7_combout ),
	.datab(\registerArray[31][19]~q ),
	.datac(\registerArray[23][19]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux44~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~8 .lut_mask = 16'hD8AA;
defparam \Mux44~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y0_N10
dffeas \registerArray[21][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[19]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][19] .is_wysiwyg = "true";
defparam \registerArray[21][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N25
dffeas \registerArray[25][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][19] .is_wysiwyg = "true";
defparam \registerArray[25][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N19
dffeas \registerArray[17][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][19] .is_wysiwyg = "true";
defparam \registerArray[17][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N24
cycloneive_lcell_comb \Mux44~0 (
// Equation(s):
// \Mux44~0_combout  = (\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o ) # ((\registerArray[25][19]~q )))) # (!\my_rf.rsel2[3]~input_o  & (!\my_rf.rsel2[2]~input_o  & ((\registerArray[17][19]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[25][19]~q ),
	.datad(\registerArray[17][19]~q ),
	.cin(gnd),
	.combout(\Mux44~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~0 .lut_mask = 16'hB9A8;
defparam \Mux44~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N28
cycloneive_lcell_comb \Mux44~1 (
// Equation(s):
// \Mux44~1_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux44~0_combout  & (\registerArray[29][19]~q )) # (!\Mux44~0_combout  & ((\registerArray[21][19]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux44~0_combout ))))

	.dataa(\registerArray[29][19]~q ),
	.datab(\registerArray[21][19]~q ),
	.datac(\my_rf.rsel2[2]~input_o ),
	.datad(\Mux44~0_combout ),
	.cin(gnd),
	.combout(\Mux44~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~1 .lut_mask = 16'hAFC0;
defparam \Mux44~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N2
cycloneive_lcell_comb \Mux44~9 (
// Equation(s):
// \Mux44~9_combout  = (\Mux44~6_combout  & (((\Mux44~8_combout )) # (!\my_rf.rsel2[0]~input_o ))) # (!\Mux44~6_combout  & (\my_rf.rsel2[0]~input_o  & ((\Mux44~1_combout ))))

	.dataa(\Mux44~6_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux44~8_combout ),
	.datad(\Mux44~1_combout ),
	.cin(gnd),
	.combout(\Mux44~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~9 .lut_mask = 16'hE6A2;
defparam \Mux44~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N20
cycloneive_lcell_comb \Mux44~20 (
// Equation(s):
// \Mux44~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux44~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux44~19_combout ))

	.dataa(gnd),
	.datab(\Mux44~19_combout ),
	.datac(\my_rf.rsel2[4]~input_o ),
	.datad(\Mux44~9_combout ),
	.cin(gnd),
	.combout(\Mux44~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~20 .lut_mask = 16'hFC0C;
defparam \Mux44~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X47_Y73_N15
cycloneive_io_ibuf \my_rf.wdat[20]~input (
	.i(\my_rf.wdat [20]),
	.ibar(gnd),
	.o(\my_rf.wdat[20]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[20]~input .bus_hold = "false";
defparam \my_rf.wdat[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X43_Y39_N29
dffeas \registerArray[9][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][20] .is_wysiwyg = "true";
defparam \registerArray[9][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y39_N21
dffeas \registerArray[10][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][20] .is_wysiwyg = "true";
defparam \registerArray[10][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N20
cycloneive_lcell_comb \Mux43~10 (
// Equation(s):
// \Mux43~10_combout  = (\my_rf.rsel2[1]~input_o  & (((\registerArray[10][20]~q ) # (\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[8][20]~q  & ((!\my_rf.rsel2[0]~input_o ))))

	.dataa(\registerArray[8][20]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[10][20]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux43~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~10 .lut_mask = 16'hCCE2;
defparam \Mux43~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N28
cycloneive_lcell_comb \Mux43~11 (
// Equation(s):
// \Mux43~11_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux43~10_combout  & (\registerArray[11][20]~q )) # (!\Mux43~10_combout  & ((\registerArray[9][20]~q ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux43~10_combout ))))

	.dataa(\registerArray[11][20]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[9][20]~q ),
	.datad(\Mux43~10_combout ),
	.cin(gnd),
	.combout(\Mux43~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~11 .lut_mask = 16'hBBC0;
defparam \Mux43~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y31_N19
dffeas \registerArray[5][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][20] .is_wysiwyg = "true";
defparam \registerArray[5][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N29
dffeas \registerArray[4][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][20] .is_wysiwyg = "true";
defparam \registerArray[4][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N18
cycloneive_lcell_comb \Mux43~12 (
// Equation(s):
// \Mux43~12_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[5][20]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[4][20]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[5][20]~q ),
	.datad(\registerArray[4][20]~q ),
	.cin(gnd),
	.combout(\Mux43~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~12 .lut_mask = 16'hB9A8;
defparam \Mux43~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y37_N29
dffeas \registerArray[6][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][20] .is_wysiwyg = "true";
defparam \registerArray[6][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N28
cycloneive_lcell_comb \Mux43~13 (
// Equation(s):
// \Mux43~13_combout  = (\Mux43~12_combout  & ((\registerArray[7][20]~q ) # ((!\my_rf.rsel2[1]~input_o )))) # (!\Mux43~12_combout  & (((\registerArray[6][20]~q  & \my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[7][20]~q ),
	.datab(\Mux43~12_combout ),
	.datac(\registerArray[6][20]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux43~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~13 .lut_mask = 16'hB8CC;
defparam \Mux43~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N0
cycloneive_lcell_comb \Mux43~16 (
// Equation(s):
// \Mux43~16_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & ((\Mux43~13_combout ))) # (!\my_rf.rsel2[2]~input_o  & (\Mux43~15_combout ))))

	.dataa(\Mux43~15_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\my_rf.rsel2[2]~input_o ),
	.datad(\Mux43~13_combout ),
	.cin(gnd),
	.combout(\Mux43~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~16 .lut_mask = 16'hF2C2;
defparam \Mux43~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N10
cycloneive_lcell_comb \Mux43~19 (
// Equation(s):
// \Mux43~19_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux43~16_combout  & (\Mux43~18_combout )) # (!\Mux43~16_combout  & ((\Mux43~11_combout ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux43~16_combout ))))

	.dataa(\Mux43~18_combout ),
	.datab(\Mux43~11_combout ),
	.datac(\my_rf.rsel2[3]~input_o ),
	.datad(\Mux43~16_combout ),
	.cin(gnd),
	.combout(\Mux43~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~19 .lut_mask = 16'hAFC0;
defparam \Mux43~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y33_N13
dffeas \registerArray[23][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][20] .is_wysiwyg = "true";
defparam \registerArray[23][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y33_N13
dffeas \registerArray[19][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][20] .is_wysiwyg = "true";
defparam \registerArray[19][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N12
cycloneive_lcell_comb \Mux43~7 (
// Equation(s):
// \Mux43~7_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\registerArray[23][20]~q )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\registerArray[19][20]~q ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[23][20]~q ),
	.datad(\registerArray[19][20]~q ),
	.cin(gnd),
	.combout(\Mux43~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~7 .lut_mask = 16'hB9A8;
defparam \Mux43~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y33_N19
dffeas \registerArray[27][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][20] .is_wysiwyg = "true";
defparam \registerArray[27][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y33_N31
dffeas \registerArray[31][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][20] .is_wysiwyg = "true";
defparam \registerArray[31][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N18
cycloneive_lcell_comb \Mux43~8 (
// Equation(s):
// \Mux43~8_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux43~7_combout  & ((\registerArray[31][20]~q ))) # (!\Mux43~7_combout  & (\registerArray[27][20]~q )))) # (!\my_rf.rsel2[3]~input_o  & (\Mux43~7_combout ))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux43~7_combout ),
	.datac(\registerArray[27][20]~q ),
	.datad(\registerArray[31][20]~q ),
	.cin(gnd),
	.combout(\Mux43~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~8 .lut_mask = 16'hEC64;
defparam \Mux43~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N25
dffeas \registerArray[21][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][20] .is_wysiwyg = "true";
defparam \registerArray[21][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N24
cycloneive_lcell_comb \Mux43~0 (
// Equation(s):
// \Mux43~0_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[21][20]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[17][20]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[17][20]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[21][20]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux43~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~0 .lut_mask = 16'hCCE2;
defparam \Mux43~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y73_N17
dffeas \registerArray[25][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[20]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][20] .is_wysiwyg = "true";
defparam \registerArray[25][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y38_N25
dffeas \registerArray[29][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][20] .is_wysiwyg = "true";
defparam \registerArray[29][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N18
cycloneive_lcell_comb \Mux43~1 (
// Equation(s):
// \Mux43~1_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux43~0_combout  & ((\registerArray[29][20]~q ))) # (!\Mux43~0_combout  & (\registerArray[25][20]~q )))) # (!\my_rf.rsel2[3]~input_o  & (\Mux43~0_combout ))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux43~0_combout ),
	.datac(\registerArray[25][20]~q ),
	.datad(\registerArray[29][20]~q ),
	.cin(gnd),
	.combout(\Mux43~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~1 .lut_mask = 16'hEC64;
defparam \Mux43~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N16
cycloneive_lcell_comb \Mux43~9 (
// Equation(s):
// \Mux43~9_combout  = (\Mux43~6_combout  & (((\Mux43~8_combout )) # (!\my_rf.rsel2[0]~input_o ))) # (!\Mux43~6_combout  & (\my_rf.rsel2[0]~input_o  & ((\Mux43~1_combout ))))

	.dataa(\Mux43~6_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux43~8_combout ),
	.datad(\Mux43~1_combout ),
	.cin(gnd),
	.combout(\Mux43~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~9 .lut_mask = 16'hE6A2;
defparam \Mux43~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N12
cycloneive_lcell_comb \Mux43~20 (
// Equation(s):
// \Mux43~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux43~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux43~19_combout ))

	.dataa(\Mux43~19_combout ),
	.datab(\Mux43~9_combout ),
	.datac(gnd),
	.datad(\my_rf.rsel2[4]~input_o ),
	.cin(gnd),
	.combout(\Mux43~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~20 .lut_mask = 16'hCCAA;
defparam \Mux43~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X0_Y32_N22
cycloneive_io_ibuf \my_rf.wdat[21]~input (
	.i(\my_rf.wdat [21]),
	.ibar(gnd),
	.o(\my_rf.wdat[21]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[21]~input .bus_hold = "false";
defparam \my_rf.wdat[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X48_Y33_N19
dffeas \registerArray[31][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][21] .is_wysiwyg = "true";
defparam \registerArray[31][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y33_N17
dffeas \registerArray[23][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][21] .is_wysiwyg = "true";
defparam \registerArray[23][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N11
dffeas \registerArray[27][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][21] .is_wysiwyg = "true";
defparam \registerArray[27][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N29
dffeas \registerArray[19][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][21] .is_wysiwyg = "true";
defparam \registerArray[19][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N10
cycloneive_lcell_comb \Mux42~7 (
// Equation(s):
// \Mux42~7_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[27][21]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[19][21]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][21]~q ),
	.datad(\registerArray[19][21]~q ),
	.cin(gnd),
	.combout(\Mux42~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~7 .lut_mask = 16'hD9C8;
defparam \Mux42~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N16
cycloneive_lcell_comb \Mux42~8 (
// Equation(s):
// \Mux42~8_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux42~7_combout  & (\registerArray[31][21]~q )) # (!\Mux42~7_combout  & ((\registerArray[23][21]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux42~7_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[31][21]~q ),
	.datac(\registerArray[23][21]~q ),
	.datad(\Mux42~7_combout ),
	.cin(gnd),
	.combout(\Mux42~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~8 .lut_mask = 16'hDDA0;
defparam \Mux42~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y38_N13
dffeas \registerArray[18][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][21] .is_wysiwyg = "true";
defparam \registerArray[18][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y37_N23
dffeas \registerArray[22][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][21] .is_wysiwyg = "true";
defparam \registerArray[22][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N22
cycloneive_lcell_comb \Mux42~2 (
// Equation(s):
// \Mux42~2_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[22][21]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[18][21]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[18][21]~q ),
	.datac(\registerArray[22][21]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux42~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~2 .lut_mask = 16'hAAE4;
defparam \Mux42~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y38_N3
dffeas \registerArray[26][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][21] .is_wysiwyg = "true";
defparam \registerArray[26][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N2
cycloneive_lcell_comb \Mux42~3 (
// Equation(s):
// \Mux42~3_combout  = (\Mux42~2_combout  & ((\registerArray[30][21]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux42~2_combout  & (((\registerArray[26][21]~q  & \my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[30][21]~q ),
	.datab(\Mux42~2_combout ),
	.datac(\registerArray[26][21]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux42~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~3 .lut_mask = 16'hB8CC;
defparam \Mux42~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y32_N16
cycloneive_lcell_comb \Mux42~6 (
// Equation(s):
// \Mux42~6_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o ) # (\Mux42~3_combout )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux42~5_combout  & (!\my_rf.rsel2[0]~input_o )))

	.dataa(\Mux42~5_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux42~3_combout ),
	.cin(gnd),
	.combout(\Mux42~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~6 .lut_mask = 16'hCEC2;
defparam \Mux42~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y32_N2
cycloneive_lcell_comb \Mux42~9 (
// Equation(s):
// \Mux42~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux42~6_combout  & ((\Mux42~8_combout ))) # (!\Mux42~6_combout  & (\Mux42~1_combout )))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux42~6_combout ))))

	.dataa(\Mux42~1_combout ),
	.datab(\Mux42~8_combout ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux42~6_combout ),
	.cin(gnd),
	.combout(\Mux42~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~9 .lut_mask = 16'hCFA0;
defparam \Mux42~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N29
dffeas \registerArray[14][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][21] .is_wysiwyg = "true";
defparam \registerArray[14][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y35_N7
dffeas \registerArray[15][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][21] .is_wysiwyg = "true";
defparam \registerArray[15][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N28
cycloneive_lcell_comb \Mux42~18 (
// Equation(s):
// \Mux42~18_combout  = (\Mux42~17_combout  & (((\registerArray[15][21]~q )) # (!\my_rf.rsel2[1]~input_o ))) # (!\Mux42~17_combout  & (\my_rf.rsel2[1]~input_o  & (\registerArray[14][21]~q )))

	.dataa(\Mux42~17_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][21]~q ),
	.datad(\registerArray[15][21]~q ),
	.cin(gnd),
	.combout(\Mux42~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~18 .lut_mask = 16'hEA62;
defparam \Mux42~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y31_N9
dffeas \registerArray[6][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][21] .is_wysiwyg = "true";
defparam \registerArray[6][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N7
dffeas \registerArray[5][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][21] .is_wysiwyg = "true";
defparam \registerArray[5][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N9
dffeas \registerArray[4][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][21] .is_wysiwyg = "true";
defparam \registerArray[4][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N6
cycloneive_lcell_comb \Mux42~10 (
// Equation(s):
// \Mux42~10_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[5][21]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[4][21]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[5][21]~q ),
	.datad(\registerArray[4][21]~q ),
	.cin(gnd),
	.combout(\Mux42~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~10 .lut_mask = 16'hB9A8;
defparam \Mux42~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y31_N8
cycloneive_lcell_comb \Mux42~11 (
// Equation(s):
// \Mux42~11_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux42~10_combout  & (\registerArray[7][21]~q )) # (!\Mux42~10_combout  & ((\registerArray[6][21]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux42~10_combout ))))

	.dataa(\registerArray[7][21]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[6][21]~q ),
	.datad(\Mux42~10_combout ),
	.cin(gnd),
	.combout(\Mux42~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~11 .lut_mask = 16'hBBC0;
defparam \Mux42~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N17
dffeas \registerArray[9][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][21] .is_wysiwyg = "true";
defparam \registerArray[9][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y39_N11
dffeas \registerArray[11][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][21] .is_wysiwyg = "true";
defparam \registerArray[11][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N16
cycloneive_lcell_comb \Mux42~13 (
// Equation(s):
// \Mux42~13_combout  = (\Mux42~12_combout  & (((\registerArray[11][21]~q )) # (!\my_rf.rsel2[0]~input_o ))) # (!\Mux42~12_combout  & (\my_rf.rsel2[0]~input_o  & (\registerArray[9][21]~q )))

	.dataa(\Mux42~12_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[9][21]~q ),
	.datad(\registerArray[11][21]~q ),
	.cin(gnd),
	.combout(\Mux42~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~13 .lut_mask = 16'hEA62;
defparam \Mux42~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y32_N13
dffeas \registerArray[2][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][21] .is_wysiwyg = "true";
defparam \registerArray[2][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y32_N12
cycloneive_lcell_comb \Mux42~15 (
// Equation(s):
// \Mux42~15_combout  = (\Mux42~14_combout ) # ((!\my_rf.rsel2[0]~input_o  & (\registerArray[2][21]~q  & \my_rf.rsel2[1]~input_o )))

	.dataa(\Mux42~14_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][21]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux42~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~15 .lut_mask = 16'hBAAA;
defparam \Mux42~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y32_N6
cycloneive_lcell_comb \Mux42~16 (
// Equation(s):
// \Mux42~16_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\Mux42~13_combout )) # (!\my_rf.rsel2[3]~input_o  & ((\Mux42~15_combout )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux42~13_combout ),
	.datad(\Mux42~15_combout ),
	.cin(gnd),
	.combout(\Mux42~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~16 .lut_mask = 16'hD9C8;
defparam \Mux42~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y32_N0
cycloneive_lcell_comb \Mux42~19 (
// Equation(s):
// \Mux42~19_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux42~16_combout  & (\Mux42~18_combout )) # (!\Mux42~16_combout  & ((\Mux42~11_combout ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux42~16_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux42~18_combout ),
	.datac(\Mux42~11_combout ),
	.datad(\Mux42~16_combout ),
	.cin(gnd),
	.combout(\Mux42~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~19 .lut_mask = 16'hDDA0;
defparam \Mux42~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y32_N10
cycloneive_lcell_comb \Mux42~20 (
// Equation(s):
// \Mux42~20_combout  = (\my_rf.rsel2[4]~input_o  & (\Mux42~9_combout )) # (!\my_rf.rsel2[4]~input_o  & ((\Mux42~19_combout )))

	.dataa(\my_rf.rsel2[4]~input_o ),
	.datab(\Mux42~9_combout ),
	.datac(gnd),
	.datad(\Mux42~19_combout ),
	.cin(gnd),
	.combout(\Mux42~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~20 .lut_mask = 16'hDD88;
defparam \Mux42~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X45_Y73_N8
cycloneive_io_ibuf \my_rf.wdat[22]~input (
	.i(\my_rf.wdat [22]),
	.ibar(gnd),
	.o(\my_rf.wdat[22]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[22]~input .bus_hold = "false";
defparam \my_rf.wdat[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X47_Y33_N23
dffeas \registerArray[27][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][22] .is_wysiwyg = "true";
defparam \registerArray[27][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y31_N17
dffeas \registerArray[23][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][22] .is_wysiwyg = "true";
defparam \registerArray[23][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N16
cycloneive_lcell_comb \Mux41~7 (
// Equation(s):
// \Mux41~7_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[23][22]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[19][22]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[19][22]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[23][22]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux41~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~7 .lut_mask = 16'hCCE2;
defparam \Mux41~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N22
cycloneive_lcell_comb \Mux41~8 (
// Equation(s):
// \Mux41~8_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux41~7_combout  & (\registerArray[31][22]~q )) # (!\Mux41~7_combout  & ((\registerArray[27][22]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux41~7_combout ))))

	.dataa(\registerArray[31][22]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][22]~q ),
	.datad(\Mux41~7_combout ),
	.cin(gnd),
	.combout(\Mux41~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~8 .lut_mask = 16'hBBC0;
defparam \Mux41~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y73_N10
dffeas \registerArray[25][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[22]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][22] .is_wysiwyg = "true";
defparam \registerArray[25][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N5
dffeas \registerArray[21][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][22] .is_wysiwyg = "true";
defparam \registerArray[21][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N4
cycloneive_lcell_comb \Mux41~0 (
// Equation(s):
// \Mux41~0_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[21][22]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[17][22]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[17][22]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[21][22]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux41~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~0 .lut_mask = 16'hCCE2;
defparam \Mux41~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y31_N20
cycloneive_lcell_comb \Mux41~1 (
// Equation(s):
// \Mux41~1_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux41~0_combout  & (\registerArray[29][22]~q )) # (!\Mux41~0_combout  & ((\registerArray[25][22]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux41~0_combout ))))

	.dataa(\registerArray[29][22]~q ),
	.datab(\registerArray[25][22]~q ),
	.datac(\my_rf.rsel2[3]~input_o ),
	.datad(\Mux41~0_combout ),
	.cin(gnd),
	.combout(\Mux41~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~1 .lut_mask = 16'hAFC0;
defparam \Mux41~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y31_N16
cycloneive_lcell_comb \Mux41~9 (
// Equation(s):
// \Mux41~9_combout  = (\Mux41~6_combout  & (((\Mux41~8_combout )) # (!\my_rf.rsel2[0]~input_o ))) # (!\Mux41~6_combout  & (\my_rf.rsel2[0]~input_o  & ((\Mux41~1_combout ))))

	.dataa(\Mux41~6_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux41~8_combout ),
	.datad(\Mux41~1_combout ),
	.cin(gnd),
	.combout(\Mux41~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~9 .lut_mask = 16'hE6A2;
defparam \Mux41~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y39_N13
dffeas \registerArray[10][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][22] .is_wysiwyg = "true";
defparam \registerArray[10][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y39_N31
dffeas \registerArray[8][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][22] .is_wysiwyg = "true";
defparam \registerArray[8][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N12
cycloneive_lcell_comb \Mux41~10 (
// Equation(s):
// \Mux41~10_combout  = (\my_rf.rsel2[0]~input_o  & (\my_rf.rsel2[1]~input_o )) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[10][22]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[8][22]~q )))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[10][22]~q ),
	.datad(\registerArray[8][22]~q ),
	.cin(gnd),
	.combout(\Mux41~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~10 .lut_mask = 16'hD9C8;
defparam \Mux41~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N13
dffeas \registerArray[9][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][22] .is_wysiwyg = "true";
defparam \registerArray[9][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N12
cycloneive_lcell_comb \Mux41~11 (
// Equation(s):
// \Mux41~11_combout  = (\Mux41~10_combout  & ((\registerArray[11][22]~q ) # ((!\my_rf.rsel2[0]~input_o )))) # (!\Mux41~10_combout  & (((\registerArray[9][22]~q  & \my_rf.rsel2[0]~input_o ))))

	.dataa(\registerArray[11][22]~q ),
	.datab(\Mux41~10_combout ),
	.datac(\registerArray[9][22]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux41~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~11 .lut_mask = 16'hB8CC;
defparam \Mux41~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N9
dffeas \registerArray[2][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][22] .is_wysiwyg = "true";
defparam \registerArray[2][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N8
cycloneive_lcell_comb \Mux41~15 (
// Equation(s):
// \Mux41~15_combout  = (\Mux41~14_combout ) # ((!\my_rf.rsel2[0]~input_o  & (\registerArray[2][22]~q  & \my_rf.rsel2[1]~input_o )))

	.dataa(\Mux41~14_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][22]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux41~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~15 .lut_mask = 16'hBAAA;
defparam \Mux41~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y31_N5
dffeas \registerArray[7][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][22] .is_wysiwyg = "true";
defparam \registerArray[7][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y31_N27
dffeas \registerArray[6][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][22] .is_wysiwyg = "true";
defparam \registerArray[6][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N5
dffeas \registerArray[4][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][22] .is_wysiwyg = "true";
defparam \registerArray[4][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N3
dffeas \registerArray[5][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][22] .is_wysiwyg = "true";
defparam \registerArray[5][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N2
cycloneive_lcell_comb \Mux41~12 (
// Equation(s):
// \Mux41~12_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[5][22]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][22]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\registerArray[4][22]~q ),
	.datac(\registerArray[5][22]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux41~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~12 .lut_mask = 16'hAAE4;
defparam \Mux41~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y31_N26
cycloneive_lcell_comb \Mux41~13 (
// Equation(s):
// \Mux41~13_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux41~12_combout  & (\registerArray[7][22]~q )) # (!\Mux41~12_combout  & ((\registerArray[6][22]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux41~12_combout ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[7][22]~q ),
	.datac(\registerArray[6][22]~q ),
	.datad(\Mux41~12_combout ),
	.cin(gnd),
	.combout(\Mux41~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~13 .lut_mask = 16'hDDA0;
defparam \Mux41~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y31_N30
cycloneive_lcell_comb \Mux41~16 (
// Equation(s):
// \Mux41~16_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & ((\Mux41~13_combout ))) # (!\my_rf.rsel2[2]~input_o  & (\Mux41~15_combout ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux41~15_combout ),
	.datac(\Mux41~13_combout ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux41~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~16 .lut_mask = 16'hFA44;
defparam \Mux41~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N25
dffeas \registerArray[14][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][22] .is_wysiwyg = "true";
defparam \registerArray[14][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y35_N11
dffeas \registerArray[15][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][22] .is_wysiwyg = "true";
defparam \registerArray[15][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N24
cycloneive_lcell_comb \Mux41~18 (
// Equation(s):
// \Mux41~18_combout  = (\Mux41~17_combout  & (((\registerArray[15][22]~q )) # (!\my_rf.rsel2[1]~input_o ))) # (!\Mux41~17_combout  & (\my_rf.rsel2[1]~input_o  & (\registerArray[14][22]~q )))

	.dataa(\Mux41~17_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][22]~q ),
	.datad(\registerArray[15][22]~q ),
	.cin(gnd),
	.combout(\Mux41~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~18 .lut_mask = 16'hEA62;
defparam \Mux41~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y31_N0
cycloneive_lcell_comb \Mux41~19 (
// Equation(s):
// \Mux41~19_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux41~16_combout  & ((\Mux41~18_combout ))) # (!\Mux41~16_combout  & (\Mux41~11_combout )))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux41~16_combout ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux41~11_combout ),
	.datac(\Mux41~16_combout ),
	.datad(\Mux41~18_combout ),
	.cin(gnd),
	.combout(\Mux41~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~19 .lut_mask = 16'hF858;
defparam \Mux41~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y31_N18
cycloneive_lcell_comb \Mux41~20 (
// Equation(s):
// \Mux41~20_combout  = (\my_rf.rsel2[4]~input_o  & (\Mux41~9_combout )) # (!\my_rf.rsel2[4]~input_o  & ((\Mux41~19_combout )))

	.dataa(\my_rf.rsel2[4]~input_o ),
	.datab(\Mux41~9_combout ),
	.datac(gnd),
	.datad(\Mux41~19_combout ),
	.cin(gnd),
	.combout(\Mux41~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~20 .lut_mask = 16'hDD88;
defparam \Mux41~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X0_Y34_N15
cycloneive_io_ibuf \my_rf.wdat[23]~input (
	.i(\my_rf.wdat [23]),
	.ibar(gnd),
	.o(\my_rf.wdat[23]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[23]~input .bus_hold = "false";
defparam \my_rf.wdat[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X48_Y33_N9
dffeas \registerArray[31][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][23] .is_wysiwyg = "true";
defparam \registerArray[31][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y33_N23
dffeas \registerArray[23][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][23] .is_wysiwyg = "true";
defparam \registerArray[23][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N9
dffeas \registerArray[27][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][23] .is_wysiwyg = "true";
defparam \registerArray[27][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N3
dffeas \registerArray[19][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][23] .is_wysiwyg = "true";
defparam \registerArray[19][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N8
cycloneive_lcell_comb \Mux40~7 (
// Equation(s):
// \Mux40~7_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[27][23]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[19][23]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][23]~q ),
	.datad(\registerArray[19][23]~q ),
	.cin(gnd),
	.combout(\Mux40~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~7 .lut_mask = 16'hD9C8;
defparam \Mux40~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N22
cycloneive_lcell_comb \Mux40~8 (
// Equation(s):
// \Mux40~8_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux40~7_combout  & (\registerArray[31][23]~q )) # (!\Mux40~7_combout  & ((\registerArray[23][23]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux40~7_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[31][23]~q ),
	.datac(\registerArray[23][23]~q ),
	.datad(\Mux40~7_combout ),
	.cin(gnd),
	.combout(\Mux40~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~8 .lut_mask = 16'hDDA0;
defparam \Mux40~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N21
dffeas \registerArray[29][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][23] .is_wysiwyg = "true";
defparam \registerArray[29][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X0_Y34_N17
dffeas \registerArray[21][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[23]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][23] .is_wysiwyg = "true";
defparam \registerArray[21][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N6
cycloneive_lcell_comb \Mux40~1 (
// Equation(s):
// \Mux40~1_combout  = (\Mux40~0_combout  & ((\registerArray[29][23]~q ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux40~0_combout  & (((\registerArray[21][23]~q  & \my_rf.rsel2[2]~input_o ))))

	.dataa(\Mux40~0_combout ),
	.datab(\registerArray[29][23]~q ),
	.datac(\registerArray[21][23]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux40~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~1 .lut_mask = 16'hD8AA;
defparam \Mux40~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N30
cycloneive_lcell_comb \Mux40~9 (
// Equation(s):
// \Mux40~9_combout  = (\Mux40~6_combout  & ((\Mux40~8_combout ) # ((!\my_rf.rsel2[0]~input_o )))) # (!\Mux40~6_combout  & (((\Mux40~1_combout  & \my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux40~6_combout ),
	.datab(\Mux40~8_combout ),
	.datac(\Mux40~1_combout ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux40~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~9 .lut_mask = 16'hD8AA;
defparam \Mux40~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y34_N15
dffeas \registerArray[12][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][23] .is_wysiwyg = "true";
defparam \registerArray[12][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y34_N21
dffeas \registerArray[13][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][23] .is_wysiwyg = "true";
defparam \registerArray[13][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N20
cycloneive_lcell_comb \Mux40~17 (
// Equation(s):
// \Mux40~17_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[13][23]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[12][23]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\registerArray[12][23]~q ),
	.datac(\registerArray[13][23]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux40~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~17 .lut_mask = 16'hAAE4;
defparam \Mux40~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N25
dffeas \registerArray[14][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][23] .is_wysiwyg = "true";
defparam \registerArray[14][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N11
dffeas \registerArray[15][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][23] .is_wysiwyg = "true";
defparam \registerArray[15][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N24
cycloneive_lcell_comb \Mux40~18 (
// Equation(s):
// \Mux40~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux40~17_combout  & ((\registerArray[15][23]~q ))) # (!\Mux40~17_combout  & (\registerArray[14][23]~q )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux40~17_combout ))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux40~17_combout ),
	.datac(\registerArray[14][23]~q ),
	.datad(\registerArray[15][23]~q ),
	.cin(gnd),
	.combout(\Mux40~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~18 .lut_mask = 16'hEC64;
defparam \Mux40~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y31_N15
dffeas \registerArray[7][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][23] .is_wysiwyg = "true";
defparam \registerArray[7][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y31_N13
dffeas \registerArray[6][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][23] .is_wysiwyg = "true";
defparam \registerArray[6][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N23
dffeas \registerArray[5][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][23] .is_wysiwyg = "true";
defparam \registerArray[5][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N25
dffeas \registerArray[4][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][23] .is_wysiwyg = "true";
defparam \registerArray[4][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N22
cycloneive_lcell_comb \Mux40~10 (
// Equation(s):
// \Mux40~10_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[5][23]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[4][23]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[5][23]~q ),
	.datad(\registerArray[4][23]~q ),
	.cin(gnd),
	.combout(\Mux40~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~10 .lut_mask = 16'hB9A8;
defparam \Mux40~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y31_N12
cycloneive_lcell_comb \Mux40~11 (
// Equation(s):
// \Mux40~11_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux40~10_combout  & (\registerArray[7][23]~q )) # (!\Mux40~10_combout  & ((\registerArray[6][23]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux40~10_combout ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[7][23]~q ),
	.datac(\registerArray[6][23]~q ),
	.datad(\Mux40~10_combout ),
	.cin(gnd),
	.combout(\Mux40~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~11 .lut_mask = 16'hDDA0;
defparam \Mux40~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N24
cycloneive_lcell_comb \Mux40~19 (
// Equation(s):
// \Mux40~19_combout  = (\Mux40~16_combout  & ((\Mux40~18_combout ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux40~16_combout  & (((\my_rf.rsel2[2]~input_o  & \Mux40~11_combout ))))

	.dataa(\Mux40~16_combout ),
	.datab(\Mux40~18_combout ),
	.datac(\my_rf.rsel2[2]~input_o ),
	.datad(\Mux40~11_combout ),
	.cin(gnd),
	.combout(\Mux40~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~19 .lut_mask = 16'hDA8A;
defparam \Mux40~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N18
cycloneive_lcell_comb \Mux40~20 (
// Equation(s):
// \Mux40~20_combout  = (\my_rf.rsel2[4]~input_o  & (\Mux40~9_combout )) # (!\my_rf.rsel2[4]~input_o  & ((\Mux40~19_combout )))

	.dataa(\my_rf.rsel2[4]~input_o ),
	.datab(gnd),
	.datac(\Mux40~9_combout ),
	.datad(\Mux40~19_combout ),
	.cin(gnd),
	.combout(\Mux40~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~20 .lut_mask = 16'hF5A0;
defparam \Mux40~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X42_Y0_N22
cycloneive_io_ibuf \my_rf.wdat[24]~input (
	.i(\my_rf.wdat [24]),
	.ibar(gnd),
	.o(\my_rf.wdat[24]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[24]~input .bus_hold = "false";
defparam \my_rf.wdat[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X47_Y34_N1
dffeas \registerArray[6][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][24] .is_wysiwyg = "true";
defparam \registerArray[6][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N11
dffeas \registerArray[5][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][24] .is_wysiwyg = "true";
defparam \registerArray[5][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N21
dffeas \registerArray[4][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][24] .is_wysiwyg = "true";
defparam \registerArray[4][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N10
cycloneive_lcell_comb \Mux39~12 (
// Equation(s):
// \Mux39~12_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[5][24]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[4][24]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[5][24]~q ),
	.datad(\registerArray[4][24]~q ),
	.cin(gnd),
	.combout(\Mux39~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~12 .lut_mask = 16'hB9A8;
defparam \Mux39~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N0
cycloneive_lcell_comb \Mux39~13 (
// Equation(s):
// \Mux39~13_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux39~12_combout  & (\registerArray[7][24]~q )) # (!\Mux39~12_combout  & ((\registerArray[6][24]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux39~12_combout ))))

	.dataa(\registerArray[7][24]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[6][24]~q ),
	.datad(\Mux39~12_combout ),
	.cin(gnd),
	.combout(\Mux39~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~13 .lut_mask = 16'hBBC0;
defparam \Mux39~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N28
cycloneive_lcell_comb \Mux39~16 (
// Equation(s):
// \Mux39~16_combout  = (\my_rf.rsel2[3]~input_o  & (((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & ((\Mux39~13_combout ))) # (!\my_rf.rsel2[2]~input_o  & (\Mux39~15_combout ))))

	.dataa(\Mux39~15_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux39~13_combout ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux39~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~16 .lut_mask = 16'hFC22;
defparam \Mux39~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N25
dffeas \registerArray[10][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][24] .is_wysiwyg = "true";
defparam \registerArray[10][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N24
cycloneive_lcell_comb \Mux39~10 (
// Equation(s):
// \Mux39~10_combout  = (\my_rf.rsel2[1]~input_o  & (((\registerArray[10][24]~q ) # (\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[8][24]~q  & ((!\my_rf.rsel2[0]~input_o ))))

	.dataa(\registerArray[8][24]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[10][24]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux39~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~10 .lut_mask = 16'hCCE2;
defparam \Mux39~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y33_N25
dffeas \registerArray[9][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][24] .is_wysiwyg = "true";
defparam \registerArray[9][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y33_N3
dffeas \registerArray[11][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][24] .is_wysiwyg = "true";
defparam \registerArray[11][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N24
cycloneive_lcell_comb \Mux39~11 (
// Equation(s):
// \Mux39~11_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux39~10_combout  & ((\registerArray[11][24]~q ))) # (!\Mux39~10_combout  & (\registerArray[9][24]~q )))) # (!\my_rf.rsel2[0]~input_o  & (\Mux39~10_combout ))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\Mux39~10_combout ),
	.datac(\registerArray[9][24]~q ),
	.datad(\registerArray[11][24]~q ),
	.cin(gnd),
	.combout(\Mux39~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~11 .lut_mask = 16'hEC64;
defparam \Mux39~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N30
cycloneive_lcell_comb \Mux39~19 (
// Equation(s):
// \Mux39~19_combout  = (\Mux39~16_combout  & ((\Mux39~18_combout ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux39~16_combout  & (((\my_rf.rsel2[3]~input_o  & \Mux39~11_combout ))))

	.dataa(\Mux39~18_combout ),
	.datab(\Mux39~16_combout ),
	.datac(\my_rf.rsel2[3]~input_o ),
	.datad(\Mux39~11_combout ),
	.cin(gnd),
	.combout(\Mux39~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~19 .lut_mask = 16'hBC8C;
defparam \Mux39~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N1
dffeas \registerArray[29][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][24] .is_wysiwyg = "true";
defparam \registerArray[29][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y0_N24
dffeas \registerArray[25][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[24]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][24] .is_wysiwyg = "true";
defparam \registerArray[25][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N10
cycloneive_lcell_comb \Mux39~1 (
// Equation(s):
// \Mux39~1_combout  = (\Mux39~0_combout  & ((\registerArray[29][24]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux39~0_combout  & (((\registerArray[25][24]~q  & \my_rf.rsel2[3]~input_o ))))

	.dataa(\Mux39~0_combout ),
	.datab(\registerArray[29][24]~q ),
	.datac(\registerArray[25][24]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux39~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~1 .lut_mask = 16'hD8AA;
defparam \Mux39~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N27
dffeas \registerArray[24][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][24] .is_wysiwyg = "true";
defparam \registerArray[24][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N29
dffeas \registerArray[16][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][24] .is_wysiwyg = "true";
defparam \registerArray[16][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N26
cycloneive_lcell_comb \Mux39~4 (
// Equation(s):
// \Mux39~4_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[24][24]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][24]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][24]~q ),
	.datad(\registerArray[16][24]~q ),
	.cin(gnd),
	.combout(\Mux39~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~4 .lut_mask = 16'hD9C8;
defparam \Mux39~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y35_N25
dffeas \registerArray[20][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][24] .is_wysiwyg = "true";
defparam \registerArray[20][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N24
cycloneive_lcell_comb \Mux39~5 (
// Equation(s):
// \Mux39~5_combout  = (\Mux39~4_combout  & ((\registerArray[28][24]~q ) # ((!\my_rf.rsel2[2]~input_o )))) # (!\Mux39~4_combout  & (((\registerArray[20][24]~q  & \my_rf.rsel2[2]~input_o ))))

	.dataa(\registerArray[28][24]~q ),
	.datab(\Mux39~4_combout ),
	.datac(\registerArray[20][24]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux39~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~5 .lut_mask = 16'hB8CC;
defparam \Mux39~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N8
cycloneive_lcell_comb \Mux39~6 (
// Equation(s):
// \Mux39~6_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux39~3_combout ) # ((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux39~5_combout  & !\my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux39~3_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\Mux39~5_combout ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux39~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~6 .lut_mask = 16'hCCB8;
defparam \Mux39~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N10
cycloneive_lcell_comb \Mux39~9 (
// Equation(s):
// \Mux39~9_combout  = (\Mux39~6_combout  & ((\Mux39~8_combout ) # ((!\my_rf.rsel2[0]~input_o )))) # (!\Mux39~6_combout  & (((\Mux39~1_combout  & \my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux39~8_combout ),
	.datab(\Mux39~1_combout ),
	.datac(\Mux39~6_combout ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux39~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~9 .lut_mask = 16'hACF0;
defparam \Mux39~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N24
cycloneive_lcell_comb \Mux39~20 (
// Equation(s):
// \Mux39~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux39~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux39~19_combout ))

	.dataa(gnd),
	.datab(\my_rf.rsel2[4]~input_o ),
	.datac(\Mux39~19_combout ),
	.datad(\Mux39~9_combout ),
	.cin(gnd),
	.combout(\Mux39~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~20 .lut_mask = 16'hFC30;
defparam \Mux39~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X0_Y33_N22
cycloneive_io_ibuf \my_rf.wdat[25]~input (
	.i(\my_rf.wdat [25]),
	.ibar(gnd),
	.o(\my_rf.wdat[25]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[25]~input .bus_hold = "false";
defparam \my_rf.wdat[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X40_Y34_N13
dffeas \registerArray[13][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][25] .is_wysiwyg = "true";
defparam \registerArray[13][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y34_N7
dffeas \registerArray[12][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][25] .is_wysiwyg = "true";
defparam \registerArray[12][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N12
cycloneive_lcell_comb \Mux38~17 (
// Equation(s):
// \Mux38~17_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[13][25]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[12][25]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[13][25]~q ),
	.datad(\registerArray[12][25]~q ),
	.cin(gnd),
	.combout(\Mux38~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~17 .lut_mask = 16'hB9A8;
defparam \Mux38~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N9
dffeas \registerArray[14][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][25] .is_wysiwyg = "true";
defparam \registerArray[14][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N3
dffeas \registerArray[15][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][25] .is_wysiwyg = "true";
defparam \registerArray[15][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N8
cycloneive_lcell_comb \Mux38~18 (
// Equation(s):
// \Mux38~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux38~17_combout  & ((\registerArray[15][25]~q ))) # (!\Mux38~17_combout  & (\registerArray[14][25]~q )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux38~17_combout ))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux38~17_combout ),
	.datac(\registerArray[14][25]~q ),
	.datad(\registerArray[15][25]~q ),
	.cin(gnd),
	.combout(\Mux38~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~18 .lut_mask = 16'hEC64;
defparam \Mux38~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y34_N15
dffeas \registerArray[1][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][25] .is_wysiwyg = "true";
defparam \registerArray[1][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y34_N21
dffeas \registerArray[3][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][25] .is_wysiwyg = "true";
defparam \registerArray[3][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N20
cycloneive_lcell_comb \Mux38~14 (
// Equation(s):
// \Mux38~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[3][25]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[1][25]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\registerArray[1][25]~q ),
	.datac(\registerArray[3][25]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux38~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~14 .lut_mask = 16'hA088;
defparam \Mux38~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N15
dffeas \registerArray[2][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][25] .is_wysiwyg = "true";
defparam \registerArray[2][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N14
cycloneive_lcell_comb \Mux38~15 (
// Equation(s):
// \Mux38~15_combout  = (\Mux38~14_combout ) # ((!\my_rf.rsel2[0]~input_o  & (\registerArray[2][25]~q  & \my_rf.rsel2[1]~input_o )))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\Mux38~14_combout ),
	.datac(\registerArray[2][25]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux38~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~15 .lut_mask = 16'hDCCC;
defparam \Mux38~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N7
dffeas \registerArray[8][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][25] .is_wysiwyg = "true";
defparam \registerArray[8][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y33_N29
dffeas \registerArray[10][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][25] .is_wysiwyg = "true";
defparam \registerArray[10][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N28
cycloneive_lcell_comb \Mux38~12 (
// Equation(s):
// \Mux38~12_combout  = (\my_rf.rsel2[1]~input_o  & (((\registerArray[10][25]~q ) # (\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[8][25]~q  & ((!\my_rf.rsel2[0]~input_o ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[8][25]~q ),
	.datac(\registerArray[10][25]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux38~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~12 .lut_mask = 16'hAAE4;
defparam \Mux38~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y33_N13
dffeas \registerArray[9][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][25] .is_wysiwyg = "true";
defparam \registerArray[9][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N12
cycloneive_lcell_comb \Mux38~13 (
// Equation(s):
// \Mux38~13_combout  = (\Mux38~12_combout  & ((\registerArray[11][25]~q ) # ((!\my_rf.rsel2[0]~input_o )))) # (!\Mux38~12_combout  & (((\registerArray[9][25]~q  & \my_rf.rsel2[0]~input_o ))))

	.dataa(\registerArray[11][25]~q ),
	.datab(\Mux38~12_combout ),
	.datac(\registerArray[9][25]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux38~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~13 .lut_mask = 16'hB8CC;
defparam \Mux38~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N8
cycloneive_lcell_comb \Mux38~16 (
// Equation(s):
// \Mux38~16_combout  = (\my_rf.rsel2[3]~input_o  & (((\Mux38~13_combout ) # (\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (\Mux38~15_combout  & ((!\my_rf.rsel2[2]~input_o ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux38~15_combout ),
	.datac(\Mux38~13_combout ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux38~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~16 .lut_mask = 16'hAAE4;
defparam \Mux38~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N29
dffeas \registerArray[5][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][25] .is_wysiwyg = "true";
defparam \registerArray[5][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N28
cycloneive_lcell_comb \Mux38~10 (
// Equation(s):
// \Mux38~10_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & ((\registerArray[5][25]~q ))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][25]~q ))))

	.dataa(\registerArray[4][25]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[5][25]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux38~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~10 .lut_mask = 16'hFC22;
defparam \Mux38~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N21
dffeas \registerArray[6][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][25] .is_wysiwyg = "true";
defparam \registerArray[6][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N20
cycloneive_lcell_comb \Mux38~11 (
// Equation(s):
// \Mux38~11_combout  = (\Mux38~10_combout  & ((\registerArray[7][25]~q ) # ((!\my_rf.rsel2[1]~input_o )))) # (!\Mux38~10_combout  & (((\registerArray[6][25]~q  & \my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[7][25]~q ),
	.datab(\Mux38~10_combout ),
	.datac(\registerArray[6][25]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux38~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~11 .lut_mask = 16'hB8CC;
defparam \Mux38~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N18
cycloneive_lcell_comb \Mux38~19 (
// Equation(s):
// \Mux38~19_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux38~16_combout  & (\Mux38~18_combout )) # (!\Mux38~16_combout  & ((\Mux38~11_combout ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux38~16_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux38~18_combout ),
	.datac(\Mux38~16_combout ),
	.datad(\Mux38~11_combout ),
	.cin(gnd),
	.combout(\Mux38~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~19 .lut_mask = 16'hDAD0;
defparam \Mux38~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N13
dffeas \registerArray[25][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][25] .is_wysiwyg = "true";
defparam \registerArray[25][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N21
dffeas \registerArray[17][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][25] .is_wysiwyg = "true";
defparam \registerArray[17][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N12
cycloneive_lcell_comb \Mux38~0 (
// Equation(s):
// \Mux38~0_combout  = (\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o ) # ((\registerArray[25][25]~q )))) # (!\my_rf.rsel2[3]~input_o  & (!\my_rf.rsel2[2]~input_o  & ((\registerArray[17][25]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[25][25]~q ),
	.datad(\registerArray[17][25]~q ),
	.cin(gnd),
	.combout(\Mux38~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~0 .lut_mask = 16'hB9A8;
defparam \Mux38~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N23
dffeas \registerArray[29][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][25] .is_wysiwyg = "true";
defparam \registerArray[29][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N16
cycloneive_lcell_comb \Mux38~1 (
// Equation(s):
// \Mux38~1_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux38~0_combout  & ((\registerArray[29][25]~q ))) # (!\Mux38~0_combout  & (\registerArray[21][25]~q )))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux38~0_combout ))))

	.dataa(\registerArray[21][25]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\Mux38~0_combout ),
	.datad(\registerArray[29][25]~q ),
	.cin(gnd),
	.combout(\Mux38~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~1 .lut_mask = 16'hF838;
defparam \Mux38~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y38_N9
dffeas \registerArray[26][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][25] .is_wysiwyg = "true";
defparam \registerArray[26][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y37_N27
dffeas \registerArray[18][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][25] .is_wysiwyg = "true";
defparam \registerArray[18][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y37_N1
dffeas \registerArray[22][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][25] .is_wysiwyg = "true";
defparam \registerArray[22][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N0
cycloneive_lcell_comb \Mux38~2 (
// Equation(s):
// \Mux38~2_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[22][25]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[18][25]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[18][25]~q ),
	.datac(\registerArray[22][25]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux38~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~2 .lut_mask = 16'hAAE4;
defparam \Mux38~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y38_N8
cycloneive_lcell_comb \Mux38~3 (
// Equation(s):
// \Mux38~3_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux38~2_combout  & (\registerArray[30][25]~q )) # (!\Mux38~2_combout  & ((\registerArray[26][25]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux38~2_combout ))))

	.dataa(\registerArray[30][25]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[26][25]~q ),
	.datad(\Mux38~2_combout ),
	.cin(gnd),
	.combout(\Mux38~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~3 .lut_mask = 16'hBBC0;
defparam \Mux38~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y38_N28
cycloneive_lcell_comb \Mux38~6 (
// Equation(s):
// \Mux38~6_combout  = (\my_rf.rsel2[0]~input_o  & (((\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\Mux38~3_combout ))) # (!\my_rf.rsel2[1]~input_o  & (\Mux38~5_combout ))))

	.dataa(\Mux38~5_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\my_rf.rsel2[1]~input_o ),
	.datad(\Mux38~3_combout ),
	.cin(gnd),
	.combout(\Mux38~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~6 .lut_mask = 16'hF2C2;
defparam \Mux38~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y38_N6
cycloneive_lcell_comb \Mux38~9 (
// Equation(s):
// \Mux38~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux38~6_combout  & (\Mux38~8_combout )) # (!\Mux38~6_combout  & ((\Mux38~1_combout ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux38~6_combout ))))

	.dataa(\Mux38~8_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux38~1_combout ),
	.datad(\Mux38~6_combout ),
	.cin(gnd),
	.combout(\Mux38~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~9 .lut_mask = 16'hBBC0;
defparam \Mux38~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y38_N24
cycloneive_lcell_comb \Mux38~20 (
// Equation(s):
// \Mux38~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux38~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux38~19_combout ))

	.dataa(gnd),
	.datab(\Mux38~19_combout ),
	.datac(\my_rf.rsel2[4]~input_o ),
	.datad(\Mux38~9_combout ),
	.cin(gnd),
	.combout(\Mux38~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~20 .lut_mask = 16'hFC0C;
defparam \Mux38~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X0_Y34_N22
cycloneive_io_ibuf \my_rf.wdat[26]~input (
	.i(\my_rf.wdat [26]),
	.ibar(gnd),
	.o(\my_rf.wdat[26]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[26]~input .bus_hold = "false";
defparam \my_rf.wdat[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X39_Y34_N25
dffeas \registerArray[14][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][26] .is_wysiwyg = "true";
defparam \registerArray[14][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y34_N17
dffeas \registerArray[13][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][26] .is_wysiwyg = "true";
defparam \registerArray[13][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N16
cycloneive_lcell_comb \Mux37~17 (
// Equation(s):
// \Mux37~17_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[13][26]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[12][26]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[12][26]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[13][26]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux37~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~17 .lut_mask = 16'hCCE2;
defparam \Mux37~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y34_N24
cycloneive_lcell_comb \Mux37~18 (
// Equation(s):
// \Mux37~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux37~17_combout  & (\registerArray[15][26]~q )) # (!\Mux37~17_combout  & ((\registerArray[14][26]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux37~17_combout ))))

	.dataa(\registerArray[15][26]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][26]~q ),
	.datad(\Mux37~17_combout ),
	.cin(gnd),
	.combout(\Mux37~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~18 .lut_mask = 16'hBBC0;
defparam \Mux37~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N17
dffeas \registerArray[5][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][26] .is_wysiwyg = "true";
defparam \registerArray[5][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N16
cycloneive_lcell_comb \Mux37~12 (
// Equation(s):
// \Mux37~12_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & ((\registerArray[5][26]~q ))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][26]~q ))))

	.dataa(\registerArray[4][26]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[5][26]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux37~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~12 .lut_mask = 16'hFC22;
defparam \Mux37~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N5
dffeas \registerArray[6][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][26] .is_wysiwyg = "true";
defparam \registerArray[6][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N4
cycloneive_lcell_comb \Mux37~13 (
// Equation(s):
// \Mux37~13_combout  = (\Mux37~12_combout  & ((\registerArray[7][26]~q ) # ((!\my_rf.rsel2[1]~input_o )))) # (!\Mux37~12_combout  & (((\registerArray[6][26]~q  & \my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[7][26]~q ),
	.datab(\Mux37~12_combout ),
	.datac(\registerArray[6][26]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux37~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~13 .lut_mask = 16'hB8CC;
defparam \Mux37~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N21
dffeas \registerArray[2][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][26] .is_wysiwyg = "true";
defparam \registerArray[2][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y34_N7
dffeas \registerArray[3][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][26] .is_wysiwyg = "true";
defparam \registerArray[3][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y34_N17
dffeas \registerArray[1][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][26] .is_wysiwyg = "true";
defparam \registerArray[1][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N6
cycloneive_lcell_comb \Mux37~14 (
// Equation(s):
// \Mux37~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][26]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][26]~q )))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[3][26]~q ),
	.datad(\registerArray[1][26]~q ),
	.cin(gnd),
	.combout(\Mux37~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~14 .lut_mask = 16'hA280;
defparam \Mux37~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N20
cycloneive_lcell_comb \Mux37~15 (
// Equation(s):
// \Mux37~15_combout  = (\Mux37~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][26]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][26]~q ),
	.datad(\Mux37~14_combout ),
	.cin(gnd),
	.combout(\Mux37~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~15 .lut_mask = 16'hFF20;
defparam \Mux37~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N28
cycloneive_lcell_comb \Mux37~16 (
// Equation(s):
// \Mux37~16_combout  = (\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o ) # ((\Mux37~13_combout )))) # (!\my_rf.rsel2[2]~input_o  & (!\my_rf.rsel2[3]~input_o  & ((\Mux37~15_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux37~13_combout ),
	.datad(\Mux37~15_combout ),
	.cin(gnd),
	.combout(\Mux37~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~16 .lut_mask = 16'hB9A8;
defparam \Mux37~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N6
cycloneive_lcell_comb \Mux37~19 (
// Equation(s):
// \Mux37~19_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux37~16_combout  & ((\Mux37~18_combout ))) # (!\Mux37~16_combout  & (\Mux37~11_combout )))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux37~16_combout ))))

	.dataa(\Mux37~11_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux37~18_combout ),
	.datad(\Mux37~16_combout ),
	.cin(gnd),
	.combout(\Mux37~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~19 .lut_mask = 16'hF388;
defparam \Mux37~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y34_N27
dffeas \registerArray[29][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][26] .is_wysiwyg = "true";
defparam \registerArray[29][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N7
dffeas \registerArray[21][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][26] .is_wysiwyg = "true";
defparam \registerArray[21][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N17
dffeas \registerArray[17][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][26] .is_wysiwyg = "true";
defparam \registerArray[17][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N6
cycloneive_lcell_comb \Mux37~0 (
// Equation(s):
// \Mux37~0_combout  = (\my_rf.rsel2[3]~input_o  & (\my_rf.rsel2[2]~input_o )) # (!\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o  & (\registerArray[21][26]~q )) # (!\my_rf.rsel2[2]~input_o  & ((\registerArray[17][26]~q )))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[21][26]~q ),
	.datad(\registerArray[17][26]~q ),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~0 .lut_mask = 16'hD9C8;
defparam \Mux37~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N24
cycloneive_lcell_comb \Mux37~1 (
// Equation(s):
// \Mux37~1_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux37~0_combout  & ((\registerArray[29][26]~q ))) # (!\Mux37~0_combout  & (\registerArray[25][26]~q )))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux37~0_combout ))))

	.dataa(\registerArray[25][26]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[29][26]~q ),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\Mux37~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~1 .lut_mask = 16'hF388;
defparam \Mux37~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y33_N19
dffeas \registerArray[27][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][26] .is_wysiwyg = "true";
defparam \registerArray[27][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y33_N13
dffeas \registerArray[31][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][26] .is_wysiwyg = "true";
defparam \registerArray[31][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N18
cycloneive_lcell_comb \Mux37~8 (
// Equation(s):
// \Mux37~8_combout  = (\Mux37~7_combout  & (((\registerArray[31][26]~q )) # (!\my_rf.rsel2[3]~input_o ))) # (!\Mux37~7_combout  & (\my_rf.rsel2[3]~input_o  & (\registerArray[27][26]~q )))

	.dataa(\Mux37~7_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][26]~q ),
	.datad(\registerArray[31][26]~q ),
	.cin(gnd),
	.combout(\Mux37~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~8 .lut_mask = 16'hEA62;
defparam \Mux37~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N4
cycloneive_lcell_comb \Mux37~9 (
// Equation(s):
// \Mux37~9_combout  = (\Mux37~6_combout  & (((\Mux37~8_combout ) # (!\my_rf.rsel2[0]~input_o )))) # (!\Mux37~6_combout  & (\Mux37~1_combout  & (\my_rf.rsel2[0]~input_o )))

	.dataa(\Mux37~6_combout ),
	.datab(\Mux37~1_combout ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux37~8_combout ),
	.cin(gnd),
	.combout(\Mux37~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~9 .lut_mask = 16'hEA4A;
defparam \Mux37~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N2
cycloneive_lcell_comb \Mux37~20 (
// Equation(s):
// \Mux37~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux37~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux37~19_combout ))

	.dataa(gnd),
	.datab(\my_rf.rsel2[4]~input_o ),
	.datac(\Mux37~19_combout ),
	.datad(\Mux37~9_combout ),
	.cin(gnd),
	.combout(\Mux37~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~20 .lut_mask = 16'hFC30;
defparam \Mux37~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X38_Y0_N8
cycloneive_io_ibuf \my_rf.wdat[27]~input (
	.i(\my_rf.wdat [27]),
	.ibar(gnd),
	.o(\my_rf.wdat[27]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[27]~input .bus_hold = "false";
defparam \my_rf.wdat[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X48_Y37_N21
dffeas \registerArray[5][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][27] .is_wysiwyg = "true";
defparam \registerArray[5][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N20
cycloneive_lcell_comb \Mux36~10 (
// Equation(s):
// \Mux36~10_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & ((\registerArray[5][27]~q ))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][27]~q ))))

	.dataa(\registerArray[4][27]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[5][27]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux36~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~10 .lut_mask = 16'hFC22;
defparam \Mux36~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N25
dffeas \registerArray[6][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][27] .is_wysiwyg = "true";
defparam \registerArray[6][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y34_N3
dffeas \registerArray[7][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][27] .is_wysiwyg = "true";
defparam \registerArray[7][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N24
cycloneive_lcell_comb \Mux36~11 (
// Equation(s):
// \Mux36~11_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux36~10_combout  & ((\registerArray[7][27]~q ))) # (!\Mux36~10_combout  & (\registerArray[6][27]~q )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux36~10_combout ))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\Mux36~10_combout ),
	.datac(\registerArray[6][27]~q ),
	.datad(\registerArray[7][27]~q ),
	.cin(gnd),
	.combout(\Mux36~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~11 .lut_mask = 16'hEC64;
defparam \Mux36~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N21
dffeas \registerArray[10][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][27] .is_wysiwyg = "true";
defparam \registerArray[10][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N20
cycloneive_lcell_comb \Mux36~12 (
// Equation(s):
// \Mux36~12_combout  = (\my_rf.rsel2[1]~input_o  & (((\registerArray[10][27]~q ) # (\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[8][27]~q  & ((!\my_rf.rsel2[0]~input_o ))))

	.dataa(\registerArray[8][27]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[10][27]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux36~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~12 .lut_mask = 16'hCCE2;
defparam \Mux36~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y33_N17
dffeas \registerArray[9][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][27] .is_wysiwyg = "true";
defparam \registerArray[9][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N16
cycloneive_lcell_comb \Mux36~13 (
// Equation(s):
// \Mux36~13_combout  = (\Mux36~12_combout  & ((\registerArray[11][27]~q ) # ((!\my_rf.rsel2[0]~input_o )))) # (!\Mux36~12_combout  & (((\registerArray[9][27]~q  & \my_rf.rsel2[0]~input_o ))))

	.dataa(\registerArray[11][27]~q ),
	.datab(\Mux36~12_combout ),
	.datac(\registerArray[9][27]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux36~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~13 .lut_mask = 16'hB8CC;
defparam \Mux36~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N17
dffeas \registerArray[2][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][27] .is_wysiwyg = "true";
defparam \registerArray[2][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y34_N23
dffeas \registerArray[1][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][27] .is_wysiwyg = "true";
defparam \registerArray[1][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y34_N13
dffeas \registerArray[3][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][27] .is_wysiwyg = "true";
defparam \registerArray[3][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N12
cycloneive_lcell_comb \Mux36~14 (
// Equation(s):
// \Mux36~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[3][27]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[1][27]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\registerArray[1][27]~q ),
	.datac(\registerArray[3][27]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux36~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~14 .lut_mask = 16'hA088;
defparam \Mux36~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N16
cycloneive_lcell_comb \Mux36~15 (
// Equation(s):
// \Mux36~15_combout  = (\Mux36~14_combout ) # ((!\my_rf.rsel2[0]~input_o  & (\my_rf.rsel2[1]~input_o  & \registerArray[2][27]~q )))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[2][27]~q ),
	.datad(\Mux36~14_combout ),
	.cin(gnd),
	.combout(\Mux36~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~15 .lut_mask = 16'hFF40;
defparam \Mux36~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N4
cycloneive_lcell_comb \Mux36~16 (
// Equation(s):
// \Mux36~16_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\Mux36~13_combout )) # (!\my_rf.rsel2[3]~input_o  & ((\Mux36~15_combout )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux36~13_combout ),
	.datad(\Mux36~15_combout ),
	.cin(gnd),
	.combout(\Mux36~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~16 .lut_mask = 16'hD9C8;
defparam \Mux36~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y34_N15
dffeas \registerArray[15][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][27] .is_wysiwyg = "true";
defparam \registerArray[15][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X39_Y34_N13
dffeas \registerArray[14][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][27] .is_wysiwyg = "true";
defparam \registerArray[14][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y34_N12
cycloneive_lcell_comb \Mux36~18 (
// Equation(s):
// \Mux36~18_combout  = (\Mux36~17_combout  & ((\registerArray[15][27]~q ) # ((!\my_rf.rsel2[1]~input_o )))) # (!\Mux36~17_combout  & (((\registerArray[14][27]~q  & \my_rf.rsel2[1]~input_o ))))

	.dataa(\Mux36~17_combout ),
	.datab(\registerArray[15][27]~q ),
	.datac(\registerArray[14][27]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux36~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~18 .lut_mask = 16'hD8AA;
defparam \Mux36~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N30
cycloneive_lcell_comb \Mux36~19 (
// Equation(s):
// \Mux36~19_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux36~16_combout  & ((\Mux36~18_combout ))) # (!\Mux36~16_combout  & (\Mux36~11_combout )))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux36~16_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux36~11_combout ),
	.datac(\Mux36~16_combout ),
	.datad(\Mux36~18_combout ),
	.cin(gnd),
	.combout(\Mux36~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~19 .lut_mask = 16'hF858;
defparam \Mux36~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N31
dffeas \registerArray[29][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][27] .is_wysiwyg = "true";
defparam \registerArray[29][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y32_N23
dffeas \registerArray[25][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][27] .is_wysiwyg = "true";
defparam \registerArray[25][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N22
cycloneive_lcell_comb \Mux36~0 (
// Equation(s):
// \Mux36~0_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & ((\registerArray[25][27]~q ))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[17][27]~q ))))

	.dataa(\registerArray[17][27]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[25][27]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux36~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~0 .lut_mask = 16'hFC22;
defparam \Mux36~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N8
cycloneive_lcell_comb \Mux36~1 (
// Equation(s):
// \Mux36~1_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux36~0_combout  & ((\registerArray[29][27]~q ))) # (!\Mux36~0_combout  & (\registerArray[21][27]~q )))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux36~0_combout ))))

	.dataa(\registerArray[21][27]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[29][27]~q ),
	.datad(\Mux36~0_combout ),
	.cin(gnd),
	.combout(\Mux36~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~1 .lut_mask = 16'hF388;
defparam \Mux36~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y34_N1
dffeas \registerArray[24][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][27] .is_wysiwyg = "true";
defparam \registerArray[24][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N17
dffeas \registerArray[16][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][27] .is_wysiwyg = "true";
defparam \registerArray[16][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N7
dffeas \registerArray[20][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][27] .is_wysiwyg = "true";
defparam \registerArray[20][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N6
cycloneive_lcell_comb \Mux36~4 (
// Equation(s):
// \Mux36~4_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[20][27]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[16][27]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[16][27]~q ),
	.datac(\registerArray[20][27]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux36~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~4 .lut_mask = 16'hAAE4;
defparam \Mux36~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N0
cycloneive_lcell_comb \Mux36~5 (
// Equation(s):
// \Mux36~5_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux36~4_combout  & (\registerArray[28][27]~q )) # (!\Mux36~4_combout  & ((\registerArray[24][27]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux36~4_combout ))))

	.dataa(\registerArray[28][27]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][27]~q ),
	.datad(\Mux36~4_combout ),
	.cin(gnd),
	.combout(\Mux36~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~5 .lut_mask = 16'hBBC0;
defparam \Mux36~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N18
cycloneive_lcell_comb \Mux36~6 (
// Equation(s):
// \Mux36~6_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux36~3_combout ) # ((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux36~5_combout  & !\my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux36~3_combout ),
	.datab(\Mux36~5_combout ),
	.datac(\my_rf.rsel2[1]~input_o ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux36~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~6 .lut_mask = 16'hF0AC;
defparam \Mux36~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N28
cycloneive_lcell_comb \Mux36~9 (
// Equation(s):
// \Mux36~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux36~6_combout  & (\Mux36~8_combout )) # (!\Mux36~6_combout  & ((\Mux36~1_combout ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux36~6_combout ))))

	.dataa(\Mux36~8_combout ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\Mux36~1_combout ),
	.datad(\Mux36~6_combout ),
	.cin(gnd),
	.combout(\Mux36~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~9 .lut_mask = 16'hBBC0;
defparam \Mux36~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N30
cycloneive_lcell_comb \Mux36~20 (
// Equation(s):
// \Mux36~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux36~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux36~19_combout ))

	.dataa(\Mux36~19_combout ),
	.datab(gnd),
	.datac(\my_rf.rsel2[4]~input_o ),
	.datad(\Mux36~9_combout ),
	.cin(gnd),
	.combout(\Mux36~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~20 .lut_mask = 16'hFA0A;
defparam \Mux36~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X0_Y35_N15
cycloneive_io_ibuf \my_rf.wdat[28]~input (
	.i(\my_rf.wdat [28]),
	.ibar(gnd),
	.o(\my_rf.wdat[28]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[28]~input .bus_hold = "false";
defparam \my_rf.wdat[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X0_Y35_N17
dffeas \registerArray[25][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[28]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][28] .is_wysiwyg = "true";
defparam \registerArray[25][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y33_N21
dffeas \registerArray[29][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][28] .is_wysiwyg = "true";
defparam \registerArray[29][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N0
cycloneive_lcell_comb \Mux35~1 (
// Equation(s):
// \Mux35~1_combout  = (\Mux35~0_combout  & (((\registerArray[29][28]~q )) # (!\my_rf.rsel2[3]~input_o ))) # (!\Mux35~0_combout  & (\my_rf.rsel2[3]~input_o  & (\registerArray[25][28]~q )))

	.dataa(\Mux35~0_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[25][28]~q ),
	.datad(\registerArray[29][28]~q ),
	.cin(gnd),
	.combout(\Mux35~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~1 .lut_mask = 16'hEA62;
defparam \Mux35~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y35_N17
dffeas \registerArray[28][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][28] .is_wysiwyg = "true";
defparam \registerArray[28][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N11
dffeas \registerArray[20][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][28] .is_wysiwyg = "true";
defparam \registerArray[20][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N31
dffeas \registerArray[24][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][28] .is_wysiwyg = "true";
defparam \registerArray[24][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N13
dffeas \registerArray[16][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][28] .is_wysiwyg = "true";
defparam \registerArray[16][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N30
cycloneive_lcell_comb \Mux35~4 (
// Equation(s):
// \Mux35~4_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[24][28]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[16][28]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[24][28]~q ),
	.datad(\registerArray[16][28]~q ),
	.cin(gnd),
	.combout(\Mux35~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~4 .lut_mask = 16'hD9C8;
defparam \Mux35~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N10
cycloneive_lcell_comb \Mux35~5 (
// Equation(s):
// \Mux35~5_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux35~4_combout  & (\registerArray[28][28]~q )) # (!\Mux35~4_combout  & ((\registerArray[20][28]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux35~4_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[28][28]~q ),
	.datac(\registerArray[20][28]~q ),
	.datad(\Mux35~4_combout ),
	.cin(gnd),
	.combout(\Mux35~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~5 .lut_mask = 16'hDDA0;
defparam \Mux35~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N8
cycloneive_lcell_comb \Mux35~6 (
// Equation(s):
// \Mux35~6_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux35~3_combout ) # ((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux35~5_combout  & !\my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux35~3_combout ),
	.datab(\Mux35~5_combout ),
	.datac(\my_rf.rsel2[1]~input_o ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux35~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~6 .lut_mask = 16'hF0AC;
defparam \Mux35~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N26
cycloneive_lcell_comb \Mux35~9 (
// Equation(s):
// \Mux35~9_combout  = (\Mux35~6_combout  & ((\Mux35~8_combout ) # ((!\my_rf.rsel2[0]~input_o )))) # (!\Mux35~6_combout  & (((\Mux35~1_combout  & \my_rf.rsel2[0]~input_o ))))

	.dataa(\Mux35~8_combout ),
	.datab(\Mux35~1_combout ),
	.datac(\Mux35~6_combout ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux35~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~9 .lut_mask = 16'hACF0;
defparam \Mux35~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y34_N17
dffeas \registerArray[14][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][28] .is_wysiwyg = "true";
defparam \registerArray[14][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X39_Y34_N19
dffeas \registerArray[15][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][28] .is_wysiwyg = "true";
defparam \registerArray[15][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y34_N16
cycloneive_lcell_comb \Mux35~18 (
// Equation(s):
// \Mux35~18_combout  = (\Mux35~17_combout  & (((\registerArray[15][28]~q )) # (!\my_rf.rsel2[1]~input_o ))) # (!\Mux35~17_combout  & (\my_rf.rsel2[1]~input_o  & (\registerArray[14][28]~q )))

	.dataa(\Mux35~17_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][28]~q ),
	.datad(\registerArray[15][28]~q ),
	.cin(gnd),
	.combout(\Mux35~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~18 .lut_mask = 16'hEA62;
defparam \Mux35~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y31_N21
dffeas \registerArray[9][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][28] .is_wysiwyg = "true";
defparam \registerArray[9][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y33_N3
dffeas \registerArray[8][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][28] .is_wysiwyg = "true";
defparam \registerArray[8][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y33_N1
dffeas \registerArray[10][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][28] .is_wysiwyg = "true";
defparam \registerArray[10][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N0
cycloneive_lcell_comb \Mux35~10 (
// Equation(s):
// \Mux35~10_combout  = (\my_rf.rsel2[1]~input_o  & (((\registerArray[10][28]~q ) # (\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[8][28]~q  & ((!\my_rf.rsel2[0]~input_o ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[8][28]~q ),
	.datac(\registerArray[10][28]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux35~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~10 .lut_mask = 16'hAAE4;
defparam \Mux35~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N20
cycloneive_lcell_comb \Mux35~11 (
// Equation(s):
// \Mux35~11_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux35~10_combout  & (\registerArray[11][28]~q )) # (!\Mux35~10_combout  & ((\registerArray[9][28]~q ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux35~10_combout ))))

	.dataa(\registerArray[11][28]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[9][28]~q ),
	.datad(\Mux35~10_combout ),
	.cin(gnd),
	.combout(\Mux35~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~11 .lut_mask = 16'hBBC0;
defparam \Mux35~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N15
dffeas \registerArray[7][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][28] .is_wysiwyg = "true";
defparam \registerArray[7][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y34_N29
dffeas \registerArray[6][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][28] .is_wysiwyg = "true";
defparam \registerArray[6][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N31
dffeas \registerArray[5][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][28] .is_wysiwyg = "true";
defparam \registerArray[5][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y31_N1
dffeas \registerArray[4][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][28] .is_wysiwyg = "true";
defparam \registerArray[4][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N30
cycloneive_lcell_comb \Mux35~12 (
// Equation(s):
// \Mux35~12_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[5][28]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[4][28]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[5][28]~q ),
	.datad(\registerArray[4][28]~q ),
	.cin(gnd),
	.combout(\Mux35~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~12 .lut_mask = 16'hB9A8;
defparam \Mux35~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N28
cycloneive_lcell_comb \Mux35~13 (
// Equation(s):
// \Mux35~13_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux35~12_combout  & (\registerArray[7][28]~q )) # (!\Mux35~12_combout  & ((\registerArray[6][28]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux35~12_combout ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[7][28]~q ),
	.datac(\registerArray[6][28]~q ),
	.datad(\Mux35~12_combout ),
	.cin(gnd),
	.combout(\Mux35~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~13 .lut_mask = 16'hDDA0;
defparam \Mux35~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N15
dffeas \registerArray[2][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][28] .is_wysiwyg = "true";
defparam \registerArray[2][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y34_N9
dffeas \registerArray[3][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][28] .is_wysiwyg = "true";
defparam \registerArray[3][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y34_N19
dffeas \registerArray[1][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][28] .is_wysiwyg = "true";
defparam \registerArray[1][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N8
cycloneive_lcell_comb \Mux35~14 (
// Equation(s):
// \Mux35~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & (\registerArray[3][28]~q )) # (!\my_rf.rsel2[1]~input_o  & ((\registerArray[1][28]~q )))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[3][28]~q ),
	.datad(\registerArray[1][28]~q ),
	.cin(gnd),
	.combout(\Mux35~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~14 .lut_mask = 16'hA280;
defparam \Mux35~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N14
cycloneive_lcell_comb \Mux35~15 (
// Equation(s):
// \Mux35~15_combout  = (\Mux35~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][28]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][28]~q ),
	.datad(\Mux35~14_combout ),
	.cin(gnd),
	.combout(\Mux35~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~15 .lut_mask = 16'hFF20;
defparam \Mux35~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N16
cycloneive_lcell_comb \Mux35~16 (
// Equation(s):
// \Mux35~16_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux35~13_combout ) # ((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux35~15_combout  & !\my_rf.rsel2[3]~input_o ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux35~13_combout ),
	.datac(\Mux35~15_combout ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux35~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~16 .lut_mask = 16'hAAD8;
defparam \Mux35~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N26
cycloneive_lcell_comb \Mux35~19 (
// Equation(s):
// \Mux35~19_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux35~16_combout  & (\Mux35~18_combout )) # (!\Mux35~16_combout  & ((\Mux35~11_combout ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux35~16_combout ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\Mux35~18_combout ),
	.datac(\Mux35~11_combout ),
	.datad(\Mux35~16_combout ),
	.cin(gnd),
	.combout(\Mux35~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~19 .lut_mask = 16'hDDA0;
defparam \Mux35~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N20
cycloneive_lcell_comb \Mux35~20 (
// Equation(s):
// \Mux35~20_combout  = (\my_rf.rsel2[4]~input_o  & (\Mux35~9_combout )) # (!\my_rf.rsel2[4]~input_o  & ((\Mux35~19_combout )))

	.dataa(\Mux35~9_combout ),
	.datab(gnd),
	.datac(\my_rf.rsel2[4]~input_o ),
	.datad(\Mux35~19_combout ),
	.cin(gnd),
	.combout(\Mux35~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~20 .lut_mask = 16'hAFA0;
defparam \Mux35~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X0_Y33_N15
cycloneive_io_ibuf \my_rf.wdat[29]~input (
	.i(\my_rf.wdat [29]),
	.ibar(gnd),
	.o(\my_rf.wdat[29]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[29]~input .bus_hold = "false";
defparam \my_rf.wdat[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X43_Y34_N31
dffeas \registerArray[2][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][29] .is_wysiwyg = "true";
defparam \registerArray[2][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y34_N31
dffeas \registerArray[1][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][29] .is_wysiwyg = "true";
defparam \registerArray[1][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y34_N29
dffeas \registerArray[3][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][29] .is_wysiwyg = "true";
defparam \registerArray[3][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N28
cycloneive_lcell_comb \Mux34~14 (
// Equation(s):
// \Mux34~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[3][29]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[1][29]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\registerArray[1][29]~q ),
	.datac(\registerArray[3][29]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux34~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~14 .lut_mask = 16'hA088;
defparam \Mux34~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N30
cycloneive_lcell_comb \Mux34~15 (
// Equation(s):
// \Mux34~15_combout  = (\Mux34~14_combout ) # ((!\my_rf.rsel2[0]~input_o  & (\my_rf.rsel2[1]~input_o  & \registerArray[2][29]~q )))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[2][29]~q ),
	.datad(\Mux34~14_combout ),
	.cin(gnd),
	.combout(\Mux34~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~15 .lut_mask = 16'hFF40;
defparam \Mux34~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y33_N21
dffeas \registerArray[11][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][29] .is_wysiwyg = "true";
defparam \registerArray[11][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y33_N19
dffeas \registerArray[9][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][29] .is_wysiwyg = "true";
defparam \registerArray[9][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y33_N15
dffeas \registerArray[8][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][29] .is_wysiwyg = "true";
defparam \registerArray[8][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y33_N13
dffeas \registerArray[10][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][29] .is_wysiwyg = "true";
defparam \registerArray[10][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N12
cycloneive_lcell_comb \Mux34~12 (
// Equation(s):
// \Mux34~12_combout  = (\my_rf.rsel2[1]~input_o  & (((\registerArray[10][29]~q ) # (\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[8][29]~q  & ((!\my_rf.rsel2[0]~input_o ))))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\registerArray[8][29]~q ),
	.datac(\registerArray[10][29]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux34~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~12 .lut_mask = 16'hAAE4;
defparam \Mux34~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N18
cycloneive_lcell_comb \Mux34~13 (
// Equation(s):
// \Mux34~13_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux34~12_combout  & (\registerArray[11][29]~q )) # (!\Mux34~12_combout  & ((\registerArray[9][29]~q ))))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux34~12_combout ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\registerArray[11][29]~q ),
	.datac(\registerArray[9][29]~q ),
	.datad(\Mux34~12_combout ),
	.cin(gnd),
	.combout(\Mux34~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~13 .lut_mask = 16'hDDA0;
defparam \Mux34~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N24
cycloneive_lcell_comb \Mux34~16 (
// Equation(s):
// \Mux34~16_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & ((\Mux34~13_combout ))) # (!\my_rf.rsel2[3]~input_o  & (\Mux34~15_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux34~15_combout ),
	.datad(\Mux34~13_combout ),
	.cin(gnd),
	.combout(\Mux34~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~16 .lut_mask = 16'hDC98;
defparam \Mux34~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N1
dffeas \registerArray[5][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][29] .is_wysiwyg = "true";
defparam \registerArray[5][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N0
cycloneive_lcell_comb \Mux34~10 (
// Equation(s):
// \Mux34~10_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o )))) # (!\my_rf.rsel2[1]~input_o  & ((\my_rf.rsel2[0]~input_o  & ((\registerArray[5][29]~q ))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[4][29]~q ))))

	.dataa(\registerArray[4][29]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[5][29]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux34~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~10 .lut_mask = 16'hFC22;
defparam \Mux34~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N13
dffeas \registerArray[6][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][29] .is_wysiwyg = "true";
defparam \registerArray[6][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N12
cycloneive_lcell_comb \Mux34~11 (
// Equation(s):
// \Mux34~11_combout  = (\Mux34~10_combout  & ((\registerArray[7][29]~q ) # ((!\my_rf.rsel2[1]~input_o )))) # (!\Mux34~10_combout  & (((\registerArray[6][29]~q  & \my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[7][29]~q ),
	.datab(\Mux34~10_combout ),
	.datac(\registerArray[6][29]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux34~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~11 .lut_mask = 16'hB8CC;
defparam \Mux34~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N5
dffeas \registerArray[14][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][29] .is_wysiwyg = "true";
defparam \registerArray[14][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y34_N29
dffeas \registerArray[13][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][29] .is_wysiwyg = "true";
defparam \registerArray[13][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N28
cycloneive_lcell_comb \Mux34~17 (
// Equation(s):
// \Mux34~17_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[13][29]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[12][29]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\registerArray[12][29]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[13][29]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux34~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~17 .lut_mask = 16'hCCE2;
defparam \Mux34~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N4
cycloneive_lcell_comb \Mux34~18 (
// Equation(s):
// \Mux34~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux34~17_combout  & (\registerArray[15][29]~q )) # (!\Mux34~17_combout  & ((\registerArray[14][29]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux34~17_combout ))))

	.dataa(\registerArray[15][29]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][29]~q ),
	.datad(\Mux34~17_combout ),
	.cin(gnd),
	.combout(\Mux34~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~18 .lut_mask = 16'hBBC0;
defparam \Mux34~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N26
cycloneive_lcell_comb \Mux34~19 (
// Equation(s):
// \Mux34~19_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux34~16_combout  & ((\Mux34~18_combout ))) # (!\Mux34~16_combout  & (\Mux34~11_combout )))) # (!\my_rf.rsel2[2]~input_o  & (\Mux34~16_combout ))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux34~16_combout ),
	.datac(\Mux34~11_combout ),
	.datad(\Mux34~18_combout ),
	.cin(gnd),
	.combout(\Mux34~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~19 .lut_mask = 16'hEC64;
defparam \Mux34~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y33_N5
dffeas \registerArray[31][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][29] .is_wysiwyg = "true";
defparam \registerArray[31][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y33_N3
dffeas \registerArray[23][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][29] .is_wysiwyg = "true";
defparam \registerArray[23][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N21
dffeas \registerArray[27][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][29] .is_wysiwyg = "true";
defparam \registerArray[27][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y31_N3
dffeas \registerArray[19][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][29] .is_wysiwyg = "true";
defparam \registerArray[19][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N20
cycloneive_lcell_comb \Mux34~7 (
// Equation(s):
// \Mux34~7_combout  = (\my_rf.rsel2[2]~input_o  & (\my_rf.rsel2[3]~input_o )) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & (\registerArray[27][29]~q )) # (!\my_rf.rsel2[3]~input_o  & ((\registerArray[19][29]~q )))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][29]~q ),
	.datad(\registerArray[19][29]~q ),
	.cin(gnd),
	.combout(\Mux34~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~7 .lut_mask = 16'hD9C8;
defparam \Mux34~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N2
cycloneive_lcell_comb \Mux34~8 (
// Equation(s):
// \Mux34~8_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux34~7_combout  & (\registerArray[31][29]~q )) # (!\Mux34~7_combout  & ((\registerArray[23][29]~q ))))) # (!\my_rf.rsel2[2]~input_o  & (((\Mux34~7_combout ))))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\registerArray[31][29]~q ),
	.datac(\registerArray[23][29]~q ),
	.datad(\Mux34~7_combout ),
	.cin(gnd),
	.combout(\Mux34~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~8 .lut_mask = 16'hDDA0;
defparam \Mux34~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y36_N5
dffeas \registerArray[30][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][29] .is_wysiwyg = "true";
defparam \registerArray[30][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y36_N3
dffeas \registerArray[26][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][29] .is_wysiwyg = "true";
defparam \registerArray[26][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N2
cycloneive_lcell_comb \Mux34~3 (
// Equation(s):
// \Mux34~3_combout  = (\Mux34~2_combout  & ((\registerArray[30][29]~q ) # ((!\my_rf.rsel2[3]~input_o )))) # (!\Mux34~2_combout  & (((\registerArray[26][29]~q  & \my_rf.rsel2[3]~input_o ))))

	.dataa(\Mux34~2_combout ),
	.datab(\registerArray[30][29]~q ),
	.datac(\registerArray[26][29]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux34~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~3 .lut_mask = 16'hD8AA;
defparam \Mux34~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N18
cycloneive_lcell_comb \Mux34~6 (
// Equation(s):
// \Mux34~6_combout  = (\my_rf.rsel2[1]~input_o  & (((\my_rf.rsel2[0]~input_o ) # (\Mux34~3_combout )))) # (!\my_rf.rsel2[1]~input_o  & (\Mux34~5_combout  & (!\my_rf.rsel2[0]~input_o )))

	.dataa(\Mux34~5_combout ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux34~3_combout ),
	.cin(gnd),
	.combout(\Mux34~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~6 .lut_mask = 16'hCEC2;
defparam \Mux34~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N12
cycloneive_lcell_comb \Mux34~9 (
// Equation(s):
// \Mux34~9_combout  = (\my_rf.rsel2[0]~input_o  & ((\Mux34~6_combout  & ((\Mux34~8_combout ))) # (!\Mux34~6_combout  & (\Mux34~1_combout )))) # (!\my_rf.rsel2[0]~input_o  & (((\Mux34~6_combout ))))

	.dataa(\Mux34~1_combout ),
	.datab(\Mux34~8_combout ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux34~6_combout ),
	.cin(gnd),
	.combout(\Mux34~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~9 .lut_mask = 16'hCFA0;
defparam \Mux34~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N28
cycloneive_lcell_comb \Mux34~20 (
// Equation(s):
// \Mux34~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux34~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux34~19_combout ))

	.dataa(gnd),
	.datab(\my_rf.rsel2[4]~input_o ),
	.datac(\Mux34~19_combout ),
	.datad(\Mux34~9_combout ),
	.cin(gnd),
	.combout(\Mux34~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~20 .lut_mask = 16'hFC30;
defparam \Mux34~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X42_Y0_N15
cycloneive_io_ibuf \my_rf.wdat[30]~input (
	.i(\my_rf.wdat [30]),
	.ibar(gnd),
	.o(\my_rf.wdat[30]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[30]~input .bus_hold = "false";
defparam \my_rf.wdat[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X42_Y35_N21
dffeas \registerArray[14][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][30] .is_wysiwyg = "true";
defparam \registerArray[14][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y35_N15
dffeas \registerArray[12][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][30] .is_wysiwyg = "true";
defparam \registerArray[12][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y35_N13
dffeas \registerArray[13][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][30] .is_wysiwyg = "true";
defparam \registerArray[13][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N12
cycloneive_lcell_comb \Mux33~17 (
// Equation(s):
// \Mux33~17_combout  = (\my_rf.rsel2[0]~input_o  & (((\registerArray[13][30]~q ) # (\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & (\registerArray[12][30]~q  & ((!\my_rf.rsel2[1]~input_o ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\registerArray[12][30]~q ),
	.datac(\registerArray[13][30]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux33~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~17 .lut_mask = 16'hAAE4;
defparam \Mux33~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N20
cycloneive_lcell_comb \Mux33~18 (
// Equation(s):
// \Mux33~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux33~17_combout  & (\registerArray[15][30]~q )) # (!\Mux33~17_combout  & ((\registerArray[14][30]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux33~17_combout ))))

	.dataa(\registerArray[15][30]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][30]~q ),
	.datad(\Mux33~17_combout ),
	.cin(gnd),
	.combout(\Mux33~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~18 .lut_mask = 16'hBBC0;
defparam \Mux33~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y39_N15
dffeas \registerArray[8][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][30] .is_wysiwyg = "true";
defparam \registerArray[8][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y39_N5
dffeas \registerArray[10][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][30] .is_wysiwyg = "true";
defparam \registerArray[10][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N4
cycloneive_lcell_comb \Mux33~10 (
// Equation(s):
// \Mux33~10_combout  = (\my_rf.rsel2[0]~input_o  & (((\my_rf.rsel2[1]~input_o )))) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[10][30]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[8][30]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\registerArray[8][30]~q ),
	.datac(\registerArray[10][30]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux33~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~10 .lut_mask = 16'hFA44;
defparam \Mux33~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N21
dffeas \registerArray[9][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][30] .is_wysiwyg = "true";
defparam \registerArray[9][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N20
cycloneive_lcell_comb \Mux33~11 (
// Equation(s):
// \Mux33~11_combout  = (\Mux33~10_combout  & ((\registerArray[11][30]~q ) # ((!\my_rf.rsel2[0]~input_o )))) # (!\Mux33~10_combout  & (((\registerArray[9][30]~q  & \my_rf.rsel2[0]~input_o ))))

	.dataa(\registerArray[11][30]~q ),
	.datab(\Mux33~10_combout ),
	.datac(\registerArray[9][30]~q ),
	.datad(\my_rf.rsel2[0]~input_o ),
	.cin(gnd),
	.combout(\Mux33~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~11 .lut_mask = 16'hB8CC;
defparam \Mux33~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N10
cycloneive_lcell_comb \Mux33~19 (
// Equation(s):
// \Mux33~19_combout  = (\Mux33~16_combout  & (((\Mux33~18_combout )) # (!\my_rf.rsel2[3]~input_o ))) # (!\Mux33~16_combout  & (\my_rf.rsel2[3]~input_o  & ((\Mux33~11_combout ))))

	.dataa(\Mux33~16_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux33~18_combout ),
	.datad(\Mux33~11_combout ),
	.cin(gnd),
	.combout(\Mux33~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~19 .lut_mask = 16'hE6A2;
defparam \Mux33~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N17
dffeas \registerArray[20][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][30] .is_wysiwyg = "true";
defparam \registerArray[20][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y37_N11
dffeas \registerArray[28][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][30] .is_wysiwyg = "true";
defparam \registerArray[28][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N16
cycloneive_lcell_comb \Mux33~5 (
// Equation(s):
// \Mux33~5_combout  = (\Mux33~4_combout  & (((\registerArray[28][30]~q )) # (!\my_rf.rsel2[2]~input_o ))) # (!\Mux33~4_combout  & (\my_rf.rsel2[2]~input_o  & (\registerArray[20][30]~q )))

	.dataa(\Mux33~4_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[20][30]~q ),
	.datad(\registerArray[28][30]~q ),
	.cin(gnd),
	.combout(\Mux33~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~5 .lut_mask = 16'hEA62;
defparam \Mux33~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y38_N21
dffeas \registerArray[26][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][30] .is_wysiwyg = "true";
defparam \registerArray[26][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N20
cycloneive_lcell_comb \Mux33~2 (
// Equation(s):
// \Mux33~2_combout  = (\my_rf.rsel2[2]~input_o  & (((\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & ((\my_rf.rsel2[3]~input_o  & ((\registerArray[26][30]~q ))) # (!\my_rf.rsel2[3]~input_o  & (\registerArray[18][30]~q ))))

	.dataa(\registerArray[18][30]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[26][30]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux33~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~2 .lut_mask = 16'hFC22;
defparam \Mux33~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y38_N31
dffeas \registerArray[22][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][30] .is_wysiwyg = "true";
defparam \registerArray[22][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y38_N25
dffeas \registerArray[30][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][30] .is_wysiwyg = "true";
defparam \registerArray[30][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N30
cycloneive_lcell_comb \Mux33~3 (
// Equation(s):
// \Mux33~3_combout  = (\my_rf.rsel2[2]~input_o  & ((\Mux33~2_combout  & ((\registerArray[30][30]~q ))) # (!\Mux33~2_combout  & (\registerArray[22][30]~q )))) # (!\my_rf.rsel2[2]~input_o  & (\Mux33~2_combout ))

	.dataa(\my_rf.rsel2[2]~input_o ),
	.datab(\Mux33~2_combout ),
	.datac(\registerArray[22][30]~q ),
	.datad(\registerArray[30][30]~q ),
	.cin(gnd),
	.combout(\Mux33~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~3 .lut_mask = 16'hEC64;
defparam \Mux33~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N28
cycloneive_lcell_comb \Mux33~6 (
// Equation(s):
// \Mux33~6_combout  = (\my_rf.rsel2[0]~input_o  & (\my_rf.rsel2[1]~input_o )) # (!\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\Mux33~3_combout ))) # (!\my_rf.rsel2[1]~input_o  & (\Mux33~5_combout ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\Mux33~5_combout ),
	.datad(\Mux33~3_combout ),
	.cin(gnd),
	.combout(\Mux33~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~6 .lut_mask = 16'hDC98;
defparam \Mux33~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N23
dffeas \registerArray[27][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][30] .is_wysiwyg = "true";
defparam \registerArray[27][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y31_N21
dffeas \registerArray[23][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][30] .is_wysiwyg = "true";
defparam \registerArray[23][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N20
cycloneive_lcell_comb \Mux33~7 (
// Equation(s):
// \Mux33~7_combout  = (\my_rf.rsel2[2]~input_o  & (((\registerArray[23][30]~q ) # (\my_rf.rsel2[3]~input_o )))) # (!\my_rf.rsel2[2]~input_o  & (\registerArray[19][30]~q  & ((!\my_rf.rsel2[3]~input_o ))))

	.dataa(\registerArray[19][30]~q ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[23][30]~q ),
	.datad(\my_rf.rsel2[3]~input_o ),
	.cin(gnd),
	.combout(\Mux33~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~7 .lut_mask = 16'hCCE2;
defparam \Mux33~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N22
cycloneive_lcell_comb \Mux33~8 (
// Equation(s):
// \Mux33~8_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux33~7_combout  & (\registerArray[31][30]~q )) # (!\Mux33~7_combout  & ((\registerArray[27][30]~q ))))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux33~7_combout ))))

	.dataa(\registerArray[31][30]~q ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\registerArray[27][30]~q ),
	.datad(\Mux33~7_combout ),
	.cin(gnd),
	.combout(\Mux33~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~8 .lut_mask = 16'hBBC0;
defparam \Mux33~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N0
cycloneive_lcell_comb \Mux33~9 (
// Equation(s):
// \Mux33~9_combout  = (\Mux33~6_combout  & (((\Mux33~8_combout ) # (!\my_rf.rsel2[0]~input_o )))) # (!\Mux33~6_combout  & (\Mux33~1_combout  & (\my_rf.rsel2[0]~input_o )))

	.dataa(\Mux33~1_combout ),
	.datab(\Mux33~6_combout ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux33~8_combout ),
	.cin(gnd),
	.combout(\Mux33~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~9 .lut_mask = 16'hEC2C;
defparam \Mux33~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N20
cycloneive_lcell_comb \Mux33~20 (
// Equation(s):
// \Mux33~20_combout  = (\my_rf.rsel2[4]~input_o  & ((\Mux33~9_combout ))) # (!\my_rf.rsel2[4]~input_o  & (\Mux33~19_combout ))

	.dataa(\Mux33~19_combout ),
	.datab(\my_rf.rsel2[4]~input_o ),
	.datac(gnd),
	.datad(\Mux33~9_combout ),
	.cin(gnd),
	.combout(\Mux33~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~20 .lut_mask = 16'hEE22;
defparam \Mux33~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N8
cycloneive_io_ibuf \my_rf.wdat[31]~input (
	.i(\my_rf.wdat [31]),
	.ibar(gnd),
	.o(\my_rf.wdat[31]~input_o ));
// synopsys translate_off
defparam \my_rf.wdat[31]~input .bus_hold = "false";
defparam \my_rf.wdat[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X45_Y32_N19
dffeas \registerArray[25][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][31] .is_wysiwyg = "true";
defparam \registerArray[25][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y38_N9
dffeas \registerArray[17][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][31] .is_wysiwyg = "true";
defparam \registerArray[17][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N18
cycloneive_lcell_comb \Mux32~0 (
// Equation(s):
// \Mux32~0_combout  = (\my_rf.rsel2[3]~input_o  & ((\my_rf.rsel2[2]~input_o ) # ((\registerArray[25][31]~q )))) # (!\my_rf.rsel2[3]~input_o  & (!\my_rf.rsel2[2]~input_o  & ((\registerArray[17][31]~q ))))

	.dataa(\my_rf.rsel2[3]~input_o ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[25][31]~q ),
	.datad(\registerArray[17][31]~q ),
	.cin(gnd),
	.combout(\Mux32~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~0 .lut_mask = 16'hB9A8;
defparam \Mux32~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y38_N27
dffeas \registerArray[29][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][31] .is_wysiwyg = "true";
defparam \registerArray[29][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N28
cycloneive_lcell_comb \Mux32~1 (
// Equation(s):
// \Mux32~1_combout  = (\Mux32~0_combout  & (((\registerArray[29][31]~q ) # (!\my_rf.rsel2[2]~input_o )))) # (!\Mux32~0_combout  & (\registerArray[21][31]~q  & ((\my_rf.rsel2[2]~input_o ))))

	.dataa(\registerArray[21][31]~q ),
	.datab(\Mux32~0_combout ),
	.datac(\registerArray[29][31]~q ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux32~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~1 .lut_mask = 16'hE2CC;
defparam \Mux32~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y33_N3
dffeas \registerArray[23][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][31] .is_wysiwyg = "true";
defparam \registerArray[23][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N21
dffeas \registerArray[31][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][31] .is_wysiwyg = "true";
defparam \registerArray[31][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N2
cycloneive_lcell_comb \Mux32~8 (
// Equation(s):
// \Mux32~8_combout  = (\Mux32~7_combout  & (((\registerArray[31][31]~q )) # (!\my_rf.rsel2[2]~input_o ))) # (!\Mux32~7_combout  & (\my_rf.rsel2[2]~input_o  & (\registerArray[23][31]~q )))

	.dataa(\Mux32~7_combout ),
	.datab(\my_rf.rsel2[2]~input_o ),
	.datac(\registerArray[23][31]~q ),
	.datad(\registerArray[31][31]~q ),
	.cin(gnd),
	.combout(\Mux32~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~8 .lut_mask = 16'hEA62;
defparam \Mux32~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N16
cycloneive_lcell_comb \Mux32~9 (
// Equation(s):
// \Mux32~9_combout  = (\Mux32~6_combout  & (((\Mux32~8_combout ) # (!\my_rf.rsel2[0]~input_o )))) # (!\Mux32~6_combout  & (\Mux32~1_combout  & (\my_rf.rsel2[0]~input_o )))

	.dataa(\Mux32~6_combout ),
	.datab(\Mux32~1_combout ),
	.datac(\my_rf.rsel2[0]~input_o ),
	.datad(\Mux32~8_combout ),
	.cin(gnd),
	.combout(\Mux32~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~9 .lut_mask = 16'hEA4A;
defparam \Mux32~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N25
dffeas \registerArray[2][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][31] .is_wysiwyg = "true";
defparam \registerArray[2][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N29
dffeas \registerArray[3][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][31] .is_wysiwyg = "true";
defparam \registerArray[3][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N28
cycloneive_lcell_comb \Mux32~14 (
// Equation(s):
// \Mux32~14_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o  & ((\registerArray[3][31]~q ))) # (!\my_rf.rsel2[1]~input_o  & (\registerArray[1][31]~q ))))

	.dataa(\registerArray[1][31]~q ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[3][31]~q ),
	.datad(\my_rf.rsel2[1]~input_o ),
	.cin(gnd),
	.combout(\Mux32~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~14 .lut_mask = 16'hC088;
defparam \Mux32~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N24
cycloneive_lcell_comb \Mux32~15 (
// Equation(s):
// \Mux32~15_combout  = (\Mux32~14_combout ) # ((\my_rf.rsel2[1]~input_o  & (!\my_rf.rsel2[0]~input_o  & \registerArray[2][31]~q )))

	.dataa(\my_rf.rsel2[1]~input_o ),
	.datab(\my_rf.rsel2[0]~input_o ),
	.datac(\registerArray[2][31]~q ),
	.datad(\Mux32~14_combout ),
	.cin(gnd),
	.combout(\Mux32~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~15 .lut_mask = 16'hFF20;
defparam \Mux32~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N18
cycloneive_lcell_comb \Mux32~16 (
// Equation(s):
// \Mux32~16_combout  = (\my_rf.rsel2[3]~input_o  & ((\Mux32~13_combout ) # ((\my_rf.rsel2[2]~input_o )))) # (!\my_rf.rsel2[3]~input_o  & (((\Mux32~15_combout  & !\my_rf.rsel2[2]~input_o ))))

	.dataa(\Mux32~13_combout ),
	.datab(\my_rf.rsel2[3]~input_o ),
	.datac(\Mux32~15_combout ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux32~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~16 .lut_mask = 16'hCCB8;
defparam \Mux32~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y36_N27
dffeas \registerArray[14][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][31] .is_wysiwyg = "true";
defparam \registerArray[14][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y36_N25
dffeas \registerArray[13][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][31] .is_wysiwyg = "true";
defparam \registerArray[13][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y36_N3
dffeas \registerArray[12][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][31] .is_wysiwyg = "true";
defparam \registerArray[12][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y36_N24
cycloneive_lcell_comb \Mux32~17 (
// Equation(s):
// \Mux32~17_combout  = (\my_rf.rsel2[0]~input_o  & ((\my_rf.rsel2[1]~input_o ) # ((\registerArray[13][31]~q )))) # (!\my_rf.rsel2[0]~input_o  & (!\my_rf.rsel2[1]~input_o  & ((\registerArray[12][31]~q ))))

	.dataa(\my_rf.rsel2[0]~input_o ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[13][31]~q ),
	.datad(\registerArray[12][31]~q ),
	.cin(gnd),
	.combout(\Mux32~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~17 .lut_mask = 16'hB9A8;
defparam \Mux32~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N26
cycloneive_lcell_comb \Mux32~18 (
// Equation(s):
// \Mux32~18_combout  = (\my_rf.rsel2[1]~input_o  & ((\Mux32~17_combout  & (\registerArray[15][31]~q )) # (!\Mux32~17_combout  & ((\registerArray[14][31]~q ))))) # (!\my_rf.rsel2[1]~input_o  & (((\Mux32~17_combout ))))

	.dataa(\registerArray[15][31]~q ),
	.datab(\my_rf.rsel2[1]~input_o ),
	.datac(\registerArray[14][31]~q ),
	.datad(\Mux32~17_combout ),
	.cin(gnd),
	.combout(\Mux32~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~18 .lut_mask = 16'hBBC0;
defparam \Mux32~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N20
cycloneive_lcell_comb \Mux32~19 (
// Equation(s):
// \Mux32~19_combout  = (\Mux32~16_combout  & (((\Mux32~18_combout ) # (!\my_rf.rsel2[2]~input_o )))) # (!\Mux32~16_combout  & (\Mux32~11_combout  & ((\my_rf.rsel2[2]~input_o ))))

	.dataa(\Mux32~11_combout ),
	.datab(\Mux32~16_combout ),
	.datac(\Mux32~18_combout ),
	.datad(\my_rf.rsel2[2]~input_o ),
	.cin(gnd),
	.combout(\Mux32~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~19 .lut_mask = 16'hE2CC;
defparam \Mux32~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N22
cycloneive_lcell_comb \Mux32~20 (
// Equation(s):
// \Mux32~20_combout  = (\my_rf.rsel2[4]~input_o  & (\Mux32~9_combout )) # (!\my_rf.rsel2[4]~input_o  & ((\Mux32~19_combout )))

	.dataa(\my_rf.rsel2[4]~input_o ),
	.datab(\Mux32~9_combout ),
	.datac(gnd),
	.datad(\Mux32~19_combout ),
	.cin(gnd),
	.combout(\Mux32~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~20 .lut_mask = 16'hDD88;
defparam \Mux32~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X38_Y0_N1
cycloneive_io_ibuf \my_rf.rsel1[4]~input (
	.i(\my_rf.rsel1 [4]),
	.ibar(gnd),
	.o(\my_rf.rsel1[4]~input_o ));
// synopsys translate_off
defparam \my_rf.rsel1[4]~input .bus_hold = "false";
defparam \my_rf.rsel1[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X53_Y33_N27
dffeas \registerArray[15][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][0] .is_wysiwyg = "true";
defparam \registerArray[15][0] .power_up = "low";
// synopsys translate_on

// Location: IOIBUF_X40_Y0_N15
cycloneive_io_ibuf \my_rf.rsel1[1]~input (
	.i(\my_rf.rsel1 [1]),
	.ibar(gnd),
	.o(\my_rf.rsel1[1]~input_o ));
// synopsys translate_off
defparam \my_rf.rsel1[1]~input .bus_hold = "false";
defparam \my_rf.rsel1[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N26
cycloneive_lcell_comb \Mux31~18 (
// Equation(s):
// \Mux31~18_combout  = (\Mux31~17_combout  & (((\registerArray[15][0]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux31~17_combout  & (\registerArray[14][0]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux31~17_combout ),
	.datab(\registerArray[14][0]~q ),
	.datac(\registerArray[15][0]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux31~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~18 .lut_mask = 16'hE4AA;
defparam \Mux31~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N1
cycloneive_io_ibuf \my_rf.rsel1[3]~input (
	.i(\my_rf.rsel1 [3]),
	.ibar(gnd),
	.o(\my_rf.rsel1[3]~input_o ));
// synopsys translate_off
defparam \my_rf.rsel1[3]~input .bus_hold = "false";
defparam \my_rf.rsel1[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y0_N22
cycloneive_io_ibuf \my_rf.rsel1[0]~input (
	.i(\my_rf.rsel1 [0]),
	.ibar(gnd),
	.o(\my_rf.rsel1[0]~input_o ));
// synopsys translate_off
defparam \my_rf.rsel1[0]~input .bus_hold = "false";
defparam \my_rf.rsel1[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: FF_X52_Y31_N3
dffeas \registerArray[11][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][0] .is_wysiwyg = "true";
defparam \registerArray[11][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N2
cycloneive_lcell_comb \Mux31~11 (
// Equation(s):
// \Mux31~11_combout  = (\Mux31~10_combout  & (((\registerArray[11][0]~q )) # (!\my_rf.rsel1[0]~input_o ))) # (!\Mux31~10_combout  & (\my_rf.rsel1[0]~input_o  & ((\registerArray[9][0]~q ))))

	.dataa(\Mux31~10_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[11][0]~q ),
	.datad(\registerArray[9][0]~q ),
	.cin(gnd),
	.combout(\Mux31~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~11 .lut_mask = 16'hE6A2;
defparam \Mux31~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N8
cycloneive_lcell_comb \Mux31~19 (
// Equation(s):
// \Mux31~19_combout  = (\Mux31~16_combout  & ((\Mux31~18_combout ) # ((!\my_rf.rsel1[3]~input_o )))) # (!\Mux31~16_combout  & (((\my_rf.rsel1[3]~input_o  & \Mux31~11_combout ))))

	.dataa(\Mux31~16_combout ),
	.datab(\Mux31~18_combout ),
	.datac(\my_rf.rsel1[3]~input_o ),
	.datad(\Mux31~11_combout ),
	.cin(gnd),
	.combout(\Mux31~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~19 .lut_mask = 16'hDA8A;
defparam \Mux31~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y28_N27
dffeas \registerArray[31][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][0] .is_wysiwyg = "true";
defparam \registerArray[31][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y28_N17
dffeas \registerArray[27][0] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[0]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][0] .is_wysiwyg = "true";
defparam \registerArray[27][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N26
cycloneive_lcell_comb \Mux31~8 (
// Equation(s):
// \Mux31~8_combout  = (\Mux31~7_combout  & (((\registerArray[31][0]~q )) # (!\my_rf.rsel1[3]~input_o ))) # (!\Mux31~7_combout  & (\my_rf.rsel1[3]~input_o  & ((\registerArray[27][0]~q ))))

	.dataa(\Mux31~7_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[31][0]~q ),
	.datad(\registerArray[27][0]~q ),
	.cin(gnd),
	.combout(\Mux31~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~8 .lut_mask = 16'hE6A2;
defparam \Mux31~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X0_Y29_N22
cycloneive_io_ibuf \my_rf.rsel1[2]~input (
	.i(\my_rf.rsel1 [2]),
	.ibar(gnd),
	.o(\my_rf.rsel1[2]~input_o ));
// synopsys translate_off
defparam \my_rf.rsel1[2]~input .bus_hold = "false";
defparam \my_rf.rsel1[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N8
cycloneive_lcell_comb \Mux31~5 (
// Equation(s):
// \Mux31~5_combout  = (\Mux31~4_combout  & (((\registerArray[28][0]~q ) # (!\my_rf.rsel1[2]~input_o )))) # (!\Mux31~4_combout  & (\registerArray[20][0]~q  & ((\my_rf.rsel1[2]~input_o ))))

	.dataa(\Mux31~4_combout ),
	.datab(\registerArray[20][0]~q ),
	.datac(\registerArray[28][0]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux31~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~5 .lut_mask = 16'hE4AA;
defparam \Mux31~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N16
cycloneive_lcell_comb \Mux31~6 (
// Equation(s):
// \Mux31~6_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\Mux31~3_combout )) # (!\my_rf.rsel1[1]~input_o  & ((\Mux31~5_combout )))))

	.dataa(\Mux31~3_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\Mux31~5_combout ),
	.cin(gnd),
	.combout(\Mux31~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~6 .lut_mask = 16'hE3E0;
defparam \Mux31~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N18
cycloneive_lcell_comb \Mux31~9 (
// Equation(s):
// \Mux31~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux31~6_combout  & ((\Mux31~8_combout ))) # (!\Mux31~6_combout  & (\Mux31~1_combout )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux31~6_combout ))))

	.dataa(\Mux31~1_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux31~8_combout ),
	.datad(\Mux31~6_combout ),
	.cin(gnd),
	.combout(\Mux31~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~9 .lut_mask = 16'hF388;
defparam \Mux31~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N10
cycloneive_lcell_comb \Mux31~20 (
// Equation(s):
// \Mux31~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux31~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux31~19_combout ))

	.dataa(gnd),
	.datab(\my_rf.rsel1[4]~input_o ),
	.datac(\Mux31~19_combout ),
	.datad(\Mux31~9_combout ),
	.cin(gnd),
	.combout(\Mux31~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~20 .lut_mask = 16'hFC30;
defparam \Mux31~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N30
cycloneive_lcell_comb \Mux30~8 (
// Equation(s):
// \Mux30~8_combout  = (\Mux30~7_combout  & (((\registerArray[31][1]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux30~7_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[23][1]~q ))))

	.dataa(\Mux30~7_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[31][1]~q ),
	.datad(\registerArray[23][1]~q ),
	.cin(gnd),
	.combout(\Mux30~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~8 .lut_mask = 16'hE6A2;
defparam \Mux30~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y32_N27
dffeas \registerArray[30][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][1] .is_wysiwyg = "true";
defparam \registerArray[30][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N26
cycloneive_lcell_comb \Mux30~3 (
// Equation(s):
// \Mux30~3_combout  = (\Mux30~2_combout  & (((\registerArray[30][1]~q )) # (!\my_rf.rsel1[3]~input_o ))) # (!\Mux30~2_combout  & (\my_rf.rsel1[3]~input_o  & ((\registerArray[26][1]~q ))))

	.dataa(\Mux30~2_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[30][1]~q ),
	.datad(\registerArray[26][1]~q ),
	.cin(gnd),
	.combout(\Mux30~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~3 .lut_mask = 16'hE6A2;
defparam \Mux30~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N28
cycloneive_lcell_comb \Mux30~6 (
// Equation(s):
// \Mux30~6_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\Mux30~3_combout ))) # (!\my_rf.rsel1[1]~input_o  & (\Mux30~5_combout ))))

	.dataa(\Mux30~5_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\Mux30~3_combout ),
	.cin(gnd),
	.combout(\Mux30~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~6 .lut_mask = 16'hF2C2;
defparam \Mux30~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N6
cycloneive_lcell_comb \Mux30~9 (
// Equation(s):
// \Mux30~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux30~6_combout  & ((\Mux30~8_combout ))) # (!\Mux30~6_combout  & (\Mux30~1_combout )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux30~6_combout ))))

	.dataa(\Mux30~1_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux30~8_combout ),
	.datad(\Mux30~6_combout ),
	.cin(gnd),
	.combout(\Mux30~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~9 .lut_mask = 16'hF388;
defparam \Mux30~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y29_N7
dffeas \registerArray[7][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][1] .is_wysiwyg = "true";
defparam \registerArray[7][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y29_N23
dffeas \registerArray[4][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][1] .is_wysiwyg = "true";
defparam \registerArray[4][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N22
cycloneive_lcell_comb \Mux30~10 (
// Equation(s):
// \Mux30~10_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o ) # ((\registerArray[5][1]~q )))) # (!\my_rf.rsel1[0]~input_o  & (!\my_rf.rsel1[1]~input_o  & (\registerArray[4][1]~q )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[4][1]~q ),
	.datad(\registerArray[5][1]~q ),
	.cin(gnd),
	.combout(\Mux30~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~10 .lut_mask = 16'hBA98;
defparam \Mux30~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N6
cycloneive_lcell_comb \Mux30~11 (
// Equation(s):
// \Mux30~11_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux30~10_combout  & ((\registerArray[7][1]~q ))) # (!\Mux30~10_combout  & (\registerArray[6][1]~q )))) # (!\my_rf.rsel1[1]~input_o  & (((\Mux30~10_combout ))))

	.dataa(\registerArray[6][1]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[7][1]~q ),
	.datad(\Mux30~10_combout ),
	.cin(gnd),
	.combout(\Mux30~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~11 .lut_mask = 16'hF388;
defparam \Mux30~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N7
dffeas \registerArray[15][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][1] .is_wysiwyg = "true";
defparam \registerArray[15][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N7
dffeas \registerArray[12][1] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[1]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][1] .is_wysiwyg = "true";
defparam \registerArray[12][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N6
cycloneive_lcell_comb \Mux30~17 (
// Equation(s):
// \Mux30~17_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[13][1]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[12][1]~q )))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[13][1]~q ),
	.datac(\registerArray[12][1]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux30~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~17 .lut_mask = 16'hEE50;
defparam \Mux30~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N6
cycloneive_lcell_comb \Mux30~18 (
// Equation(s):
// \Mux30~18_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux30~17_combout  & ((\registerArray[15][1]~q ))) # (!\Mux30~17_combout  & (\registerArray[14][1]~q )))) # (!\my_rf.rsel1[1]~input_o  & (((\Mux30~17_combout ))))

	.dataa(\registerArray[14][1]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][1]~q ),
	.datad(\Mux30~17_combout ),
	.cin(gnd),
	.combout(\Mux30~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~18 .lut_mask = 16'hF388;
defparam \Mux30~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N4
cycloneive_lcell_comb \Mux30~19 (
// Equation(s):
// \Mux30~19_combout  = (\Mux30~16_combout  & (((\Mux30~18_combout ) # (!\my_rf.rsel1[2]~input_o )))) # (!\Mux30~16_combout  & (\Mux30~11_combout  & (\my_rf.rsel1[2]~input_o )))

	.dataa(\Mux30~16_combout ),
	.datab(\Mux30~11_combout ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux30~18_combout ),
	.cin(gnd),
	.combout(\Mux30~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~19 .lut_mask = 16'hEA4A;
defparam \Mux30~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N14
cycloneive_lcell_comb \Mux30~20 (
// Equation(s):
// \Mux30~20_combout  = (\my_rf.rsel1[4]~input_o  & (\Mux30~9_combout )) # (!\my_rf.rsel1[4]~input_o  & ((\Mux30~19_combout )))

	.dataa(\Mux30~9_combout ),
	.datab(\Mux30~19_combout ),
	.datac(gnd),
	.datad(\my_rf.rsel1[4]~input_o ),
	.cin(gnd),
	.combout(\Mux30~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~20 .lut_mask = 16'hAACC;
defparam \Mux30~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y31_N3
dffeas \registerArray[11][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][2] .is_wysiwyg = "true";
defparam \registerArray[11][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y31_N25
dffeas \registerArray[9][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][2] .is_wysiwyg = "true";
defparam \registerArray[9][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N2
cycloneive_lcell_comb \Mux29~11 (
// Equation(s):
// \Mux29~11_combout  = (\Mux29~10_combout  & (((\registerArray[11][2]~q )) # (!\my_rf.rsel1[0]~input_o ))) # (!\Mux29~10_combout  & (\my_rf.rsel1[0]~input_o  & ((\registerArray[9][2]~q ))))

	.dataa(\Mux29~10_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[11][2]~q ),
	.datad(\registerArray[9][2]~q ),
	.cin(gnd),
	.combout(\Mux29~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~11 .lut_mask = 16'hE6A2;
defparam \Mux29~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N18
cycloneive_lcell_comb \Mux29~18 (
// Equation(s):
// \Mux29~18_combout  = (\Mux29~17_combout  & (((\registerArray[15][2]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux29~17_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[14][2]~q ))))

	.dataa(\Mux29~17_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][2]~q ),
	.datad(\registerArray[14][2]~q ),
	.cin(gnd),
	.combout(\Mux29~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~18 .lut_mask = 16'hE6A2;
defparam \Mux29~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N24
cycloneive_lcell_comb \Mux29~19 (
// Equation(s):
// \Mux29~19_combout  = (\Mux29~16_combout  & (((\Mux29~18_combout )) # (!\my_rf.rsel1[3]~input_o ))) # (!\Mux29~16_combout  & (\my_rf.rsel1[3]~input_o  & (\Mux29~11_combout )))

	.dataa(\Mux29~16_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\Mux29~11_combout ),
	.datad(\Mux29~18_combout ),
	.cin(gnd),
	.combout(\Mux29~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~19 .lut_mask = 16'hEA62;
defparam \Mux29~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y0_N24
dffeas \registerArray[25][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[2]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][2] .is_wysiwyg = "true";
defparam \registerArray[25][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y38_N26
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// \Mux29~1_combout  = (\Mux29~0_combout  & (((\registerArray[29][2]~q ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux29~0_combout  & (\registerArray[25][2]~q  & ((\my_rf.rsel1[3]~input_o ))))

	.dataa(\Mux29~0_combout ),
	.datab(\registerArray[25][2]~q ),
	.datac(\registerArray[29][2]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'hE4AA;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y31_N5
dffeas \registerArray[24][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][2] .is_wysiwyg = "true";
defparam \registerArray[24][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y31_N23
dffeas \registerArray[16][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][2] .is_wysiwyg = "true";
defparam \registerArray[16][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N22
cycloneive_lcell_comb \Mux29~4 (
// Equation(s):
// \Mux29~4_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[24][2]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[16][2]~q )))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[24][2]~q ),
	.datac(\registerArray[16][2]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux29~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~4 .lut_mask = 16'hEE50;
defparam \Mux29~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N29
dffeas \registerArray[28][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][2] .is_wysiwyg = "true";
defparam \registerArray[28][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y35_N3
dffeas \registerArray[20][2] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[2]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][2] .is_wysiwyg = "true";
defparam \registerArray[20][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N28
cycloneive_lcell_comb \Mux29~5 (
// Equation(s):
// \Mux29~5_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux29~4_combout  & (\registerArray[28][2]~q )) # (!\Mux29~4_combout  & ((\registerArray[20][2]~q ))))) # (!\my_rf.rsel1[2]~input_o  & (\Mux29~4_combout ))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux29~4_combout ),
	.datac(\registerArray[28][2]~q ),
	.datad(\registerArray[20][2]~q ),
	.cin(gnd),
	.combout(\Mux29~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~5 .lut_mask = 16'hE6C4;
defparam \Mux29~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N0
cycloneive_lcell_comb \Mux29~6 (
// Equation(s):
// \Mux29~6_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\Mux29~3_combout )) # (!\my_rf.rsel1[1]~input_o  & ((\Mux29~5_combout )))))

	.dataa(\Mux29~3_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\Mux29~5_combout ),
	.cin(gnd),
	.combout(\Mux29~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~6 .lut_mask = 16'hE3E0;
defparam \Mux29~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N2
cycloneive_lcell_comb \Mux29~9 (
// Equation(s):
// \Mux29~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux29~6_combout  & (\Mux29~8_combout )) # (!\Mux29~6_combout  & ((\Mux29~1_combout ))))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux29~6_combout ))))

	.dataa(\Mux29~8_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux29~1_combout ),
	.datad(\Mux29~6_combout ),
	.cin(gnd),
	.combout(\Mux29~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~9 .lut_mask = 16'hBBC0;
defparam \Mux29~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N10
cycloneive_lcell_comb \Mux29~20 (
// Equation(s):
// \Mux29~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux29~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux29~19_combout ))

	.dataa(\my_rf.rsel1[4]~input_o ),
	.datab(\Mux29~19_combout ),
	.datac(gnd),
	.datad(\Mux29~9_combout ),
	.cin(gnd),
	.combout(\Mux29~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~20 .lut_mask = 16'hEE44;
defparam \Mux29~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y28_N15
dffeas \registerArray[31][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][3] .is_wysiwyg = "true";
defparam \registerArray[31][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y28_N14
cycloneive_lcell_comb \Mux28~8 (
// Equation(s):
// \Mux28~8_combout  = (\Mux28~7_combout  & (((\registerArray[31][3]~q ) # (!\my_rf.rsel1[2]~input_o )))) # (!\Mux28~7_combout  & (\registerArray[23][3]~q  & ((\my_rf.rsel1[2]~input_o ))))

	.dataa(\Mux28~7_combout ),
	.datab(\registerArray[23][3]~q ),
	.datac(\registerArray[31][3]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux28~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~8 .lut_mask = 16'hE4AA;
defparam \Mux28~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y32_N23
dffeas \registerArray[30][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][3] .is_wysiwyg = "true";
defparam \registerArray[30][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y32_N13
dffeas \registerArray[26][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][3] .is_wysiwyg = "true";
defparam \registerArray[26][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N22
cycloneive_lcell_comb \Mux28~3 (
// Equation(s):
// \Mux28~3_combout  = (\Mux28~2_combout  & (((\registerArray[30][3]~q )) # (!\my_rf.rsel1[3]~input_o ))) # (!\Mux28~2_combout  & (\my_rf.rsel1[3]~input_o  & ((\registerArray[26][3]~q ))))

	.dataa(\Mux28~2_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[30][3]~q ),
	.datad(\registerArray[26][3]~q ),
	.cin(gnd),
	.combout(\Mux28~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~3 .lut_mask = 16'hE6A2;
defparam \Mux28~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N31
dffeas \registerArray[24][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][3] .is_wysiwyg = "true";
defparam \registerArray[24][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N9
dffeas \registerArray[28][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][3] .is_wysiwyg = "true";
defparam \registerArray[28][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N8
cycloneive_lcell_comb \Mux28~5 (
// Equation(s):
// \Mux28~5_combout  = (\Mux28~4_combout  & (((\registerArray[28][3]~q ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux28~4_combout  & (\registerArray[24][3]~q  & ((\my_rf.rsel1[3]~input_o ))))

	.dataa(\Mux28~4_combout ),
	.datab(\registerArray[24][3]~q ),
	.datac(\registerArray[28][3]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux28~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~5 .lut_mask = 16'hE4AA;
defparam \Mux28~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N28
cycloneive_lcell_comb \Mux28~6 (
// Equation(s):
// \Mux28~6_combout  = (\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o )) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\Mux28~3_combout )) # (!\my_rf.rsel1[1]~input_o  & ((\Mux28~5_combout )))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\Mux28~3_combout ),
	.datad(\Mux28~5_combout ),
	.cin(gnd),
	.combout(\Mux28~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~6 .lut_mask = 16'hD9C8;
defparam \Mux28~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N30
cycloneive_lcell_comb \Mux28~9 (
// Equation(s):
// \Mux28~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux28~6_combout  & ((\Mux28~8_combout ))) # (!\Mux28~6_combout  & (\Mux28~1_combout )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux28~6_combout ))))

	.dataa(\Mux28~1_combout ),
	.datab(\Mux28~8_combout ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\Mux28~6_combout ),
	.cin(gnd),
	.combout(\Mux28~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~9 .lut_mask = 16'hCFA0;
defparam \Mux28~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N24
cycloneive_lcell_comb \Mux28~15 (
// Equation(s):
// \Mux28~15_combout  = (\Mux28~14_combout ) # ((\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & \registerArray[2][3]~q )))

	.dataa(\Mux28~14_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\registerArray[2][3]~q ),
	.cin(gnd),
	.combout(\Mux28~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~15 .lut_mask = 16'hAEAA;
defparam \Mux28~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N18
cycloneive_lcell_comb \Mux28~16 (
// Equation(s):
// \Mux28~16_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux28~13_combout ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((!\my_rf.rsel1[2]~input_o  & \Mux28~15_combout ))))

	.dataa(\Mux28~13_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux28~15_combout ),
	.cin(gnd),
	.combout(\Mux28~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~16 .lut_mask = 16'hCBC8;
defparam \Mux28~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N31
dffeas \registerArray[15][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][3] .is_wysiwyg = "true";
defparam \registerArray[15][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N30
cycloneive_lcell_comb \Mux28~18 (
// Equation(s):
// \Mux28~18_combout  = (\Mux28~17_combout  & (((\registerArray[15][3]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux28~17_combout  & (\registerArray[14][3]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux28~17_combout ),
	.datab(\registerArray[14][3]~q ),
	.datac(\registerArray[15][3]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux28~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~18 .lut_mask = 16'hE4AA;
defparam \Mux28~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y29_N31
dffeas \registerArray[4][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][3] .is_wysiwyg = "true";
defparam \registerArray[4][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y29_N13
dffeas \registerArray[5][3] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[3]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][3] .is_wysiwyg = "true";
defparam \registerArray[5][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y29_N30
cycloneive_lcell_comb \Mux28~10 (
// Equation(s):
// \Mux28~10_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o ) # ((\registerArray[5][3]~q )))) # (!\my_rf.rsel1[0]~input_o  & (!\my_rf.rsel1[1]~input_o  & (\registerArray[4][3]~q )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[4][3]~q ),
	.datad(\registerArray[5][3]~q ),
	.cin(gnd),
	.combout(\Mux28~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~10 .lut_mask = 16'hBA98;
defparam \Mux28~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N14
cycloneive_lcell_comb \Mux28~11 (
// Equation(s):
// \Mux28~11_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux28~10_combout  & (\registerArray[7][3]~q )) # (!\Mux28~10_combout  & ((\registerArray[6][3]~q ))))) # (!\my_rf.rsel1[1]~input_o  & (\Mux28~10_combout ))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\Mux28~10_combout ),
	.datac(\registerArray[7][3]~q ),
	.datad(\registerArray[6][3]~q ),
	.cin(gnd),
	.combout(\Mux28~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~11 .lut_mask = 16'hE6C4;
defparam \Mux28~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N20
cycloneive_lcell_comb \Mux28~19 (
// Equation(s):
// \Mux28~19_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux28~16_combout  & (\Mux28~18_combout )) # (!\Mux28~16_combout  & ((\Mux28~11_combout ))))) # (!\my_rf.rsel1[2]~input_o  & (\Mux28~16_combout ))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux28~16_combout ),
	.datac(\Mux28~18_combout ),
	.datad(\Mux28~11_combout ),
	.cin(gnd),
	.combout(\Mux28~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~19 .lut_mask = 16'hE6C4;
defparam \Mux28~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N14
cycloneive_lcell_comb \Mux28~20 (
// Equation(s):
// \Mux28~20_combout  = (\my_rf.rsel1[4]~input_o  & (\Mux28~9_combout )) # (!\my_rf.rsel1[4]~input_o  & ((\Mux28~19_combout )))

	.dataa(\Mux28~9_combout ),
	.datab(\Mux28~19_combout ),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux28~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~20 .lut_mask = 16'hACAC;
defparam \Mux28~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y31_N27
dffeas \registerArray[8][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][4] .is_wysiwyg = "true";
defparam \registerArray[8][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N26
cycloneive_lcell_comb \Mux27~10 (
// Equation(s):
// \Mux27~10_combout  = (\my_rf.rsel1[1]~input_o  & ((\registerArray[10][4]~q ) # ((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & (((\registerArray[8][4]~q  & !\my_rf.rsel1[0]~input_o ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[10][4]~q ),
	.datac(\registerArray[8][4]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux27~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~10 .lut_mask = 16'hAAD8;
defparam \Mux27~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y31_N11
dffeas \registerArray[11][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][4] .is_wysiwyg = "true";
defparam \registerArray[11][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N10
cycloneive_lcell_comb \Mux27~11 (
// Equation(s):
// \Mux27~11_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux27~10_combout  & (\registerArray[11][4]~q )) # (!\Mux27~10_combout  & ((\registerArray[9][4]~q ))))) # (!\my_rf.rsel1[0]~input_o  & (\Mux27~10_combout ))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux27~10_combout ),
	.datac(\registerArray[11][4]~q ),
	.datad(\registerArray[9][4]~q ),
	.cin(gnd),
	.combout(\Mux27~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~11 .lut_mask = 16'hE6C4;
defparam \Mux27~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y31_N9
dffeas \registerArray[3][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][4] .is_wysiwyg = "true";
defparam \registerArray[3][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N11
dffeas \registerArray[1][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][4] .is_wysiwyg = "true";
defparam \registerArray[1][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N10
cycloneive_lcell_comb \Mux27~14 (
// Equation(s):
// \Mux27~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\registerArray[3][4]~q )) # (!\my_rf.rsel1[1]~input_o  & ((\registerArray[1][4]~q )))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\registerArray[3][4]~q ),
	.datac(\registerArray[1][4]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux27~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~14 .lut_mask = 16'h88A0;
defparam \Mux27~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N23
dffeas \registerArray[2][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][4] .is_wysiwyg = "true";
defparam \registerArray[2][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N10
cycloneive_lcell_comb \Mux27~15 (
// Equation(s):
// \Mux27~15_combout  = (\Mux27~14_combout ) # ((!\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o  & \registerArray[2][4]~q )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux27~14_combout ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\registerArray[2][4]~q ),
	.cin(gnd),
	.combout(\Mux27~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~15 .lut_mask = 16'hDCCC;
defparam \Mux27~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N4
cycloneive_lcell_comb \Mux27~16 (
// Equation(s):
// \Mux27~16_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & (\Mux27~13_combout )) # (!\my_rf.rsel1[2]~input_o  & ((\Mux27~15_combout )))))

	.dataa(\Mux27~13_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux27~15_combout ),
	.cin(gnd),
	.combout(\Mux27~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~16 .lut_mask = 16'hE3E0;
defparam \Mux27~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N22
cycloneive_lcell_comb \Mux27~19 (
// Equation(s):
// \Mux27~19_combout  = (\Mux27~16_combout  & ((\Mux27~18_combout ) # ((!\my_rf.rsel1[3]~input_o )))) # (!\Mux27~16_combout  & (((\Mux27~11_combout  & \my_rf.rsel1[3]~input_o ))))

	.dataa(\Mux27~18_combout ),
	.datab(\Mux27~11_combout ),
	.datac(\Mux27~16_combout ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux27~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~19 .lut_mask = 16'hACF0;
defparam \Mux27~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N19
dffeas \registerArray[29][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][4] .is_wysiwyg = "true";
defparam \registerArray[29][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N10
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o ) # ((\registerArray[21][4]~q )))) # (!\my_rf.rsel1[2]~input_o  & (!\my_rf.rsel1[3]~input_o  & (\registerArray[17][4]~q )))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[17][4]~q ),
	.datad(\registerArray[21][4]~q ),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'hBA98;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N18
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// \Mux27~1_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux27~0_combout  & ((\registerArray[29][4]~q ))) # (!\Mux27~0_combout  & (\registerArray[25][4]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux27~0_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[25][4]~q ),
	.datac(\registerArray[29][4]~q ),
	.datad(\Mux27~0_combout ),
	.cin(gnd),
	.combout(\Mux27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hF588;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y31_N28
cycloneive_lcell_comb \Mux27~4 (
// Equation(s):
// \Mux27~4_combout  = (\my_rf.rsel1[2]~input_o  & (\my_rf.rsel1[3]~input_o )) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & ((\registerArray[24][4]~q ))) # (!\my_rf.rsel1[3]~input_o  & (\registerArray[16][4]~q ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[16][4]~q ),
	.datad(\registerArray[24][4]~q ),
	.cin(gnd),
	.combout(\Mux27~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~4 .lut_mask = 16'hDC98;
defparam \Mux27~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N26
cycloneive_lcell_comb \Mux27~5 (
// Equation(s):
// \Mux27~5_combout  = (\Mux27~4_combout  & (((\registerArray[28][4]~q ) # (!\my_rf.rsel1[2]~input_o )))) # (!\Mux27~4_combout  & (\registerArray[20][4]~q  & ((\my_rf.rsel1[2]~input_o ))))

	.dataa(\registerArray[20][4]~q ),
	.datab(\Mux27~4_combout ),
	.datac(\registerArray[28][4]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux27~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~5 .lut_mask = 16'hE2CC;
defparam \Mux27~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N8
cycloneive_lcell_comb \Mux27~6 (
// Equation(s):
// \Mux27~6_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux27~3_combout ) # ((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & (((!\my_rf.rsel1[0]~input_o  & \Mux27~5_combout ))))

	.dataa(\Mux27~3_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\Mux27~5_combout ),
	.cin(gnd),
	.combout(\Mux27~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~6 .lut_mask = 16'hCBC8;
defparam \Mux27~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y28_N27
dffeas \registerArray[19][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][4] .is_wysiwyg = "true";
defparam \registerArray[19][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N17
dffeas \registerArray[23][4] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[4]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][4] .is_wysiwyg = "true";
defparam \registerArray[23][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N26
cycloneive_lcell_comb \Mux27~7 (
// Equation(s):
// \Mux27~7_combout  = (\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o ) # ((\registerArray[23][4]~q )))) # (!\my_rf.rsel1[2]~input_o  & (!\my_rf.rsel1[3]~input_o  & (\registerArray[19][4]~q )))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[19][4]~q ),
	.datad(\registerArray[23][4]~q ),
	.cin(gnd),
	.combout(\Mux27~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~7 .lut_mask = 16'hBA98;
defparam \Mux27~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N18
cycloneive_lcell_comb \Mux27~8 (
// Equation(s):
// \Mux27~8_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux27~7_combout  & (\registerArray[31][4]~q )) # (!\Mux27~7_combout  & ((\registerArray[27][4]~q ))))) # (!\my_rf.rsel1[3]~input_o  & (\Mux27~7_combout ))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux27~7_combout ),
	.datac(\registerArray[31][4]~q ),
	.datad(\registerArray[27][4]~q ),
	.cin(gnd),
	.combout(\Mux27~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~8 .lut_mask = 16'hE6C4;
defparam \Mux27~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N2
cycloneive_lcell_comb \Mux27~9 (
// Equation(s):
// \Mux27~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux27~6_combout  & ((\Mux27~8_combout ))) # (!\Mux27~6_combout  & (\Mux27~1_combout )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux27~6_combout ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux27~1_combout ),
	.datac(\Mux27~6_combout ),
	.datad(\Mux27~8_combout ),
	.cin(gnd),
	.combout(\Mux27~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~9 .lut_mask = 16'hF858;
defparam \Mux27~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y32_N4
cycloneive_lcell_comb \Mux27~20 (
// Equation(s):
// \Mux27~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux27~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux27~19_combout ))

	.dataa(gnd),
	.datab(\Mux27~19_combout ),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux27~9_combout ),
	.cin(gnd),
	.combout(\Mux27~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~20 .lut_mask = 16'hFC0C;
defparam \Mux27~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y29_N5
dffeas \registerArray[6][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][5] .is_wysiwyg = "true";
defparam \registerArray[6][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y29_N23
dffeas \registerArray[7][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][5] .is_wysiwyg = "true";
defparam \registerArray[7][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N22
cycloneive_lcell_comb \Mux26~11 (
// Equation(s):
// \Mux26~11_combout  = (\Mux26~10_combout  & (((\registerArray[7][5]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux26~10_combout  & (\registerArray[6][5]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux26~10_combout ),
	.datab(\registerArray[6][5]~q ),
	.datac(\registerArray[7][5]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux26~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~11 .lut_mask = 16'hE4AA;
defparam \Mux26~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y31_N15
dffeas \registerArray[8][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][5] .is_wysiwyg = "true";
defparam \registerArray[8][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y31_N29
dffeas \registerArray[10][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][5] .is_wysiwyg = "true";
defparam \registerArray[10][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N14
cycloneive_lcell_comb \Mux26~12 (
// Equation(s):
// \Mux26~12_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\registerArray[10][5]~q )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & (\registerArray[8][5]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[8][5]~q ),
	.datad(\registerArray[10][5]~q ),
	.cin(gnd),
	.combout(\Mux26~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~12 .lut_mask = 16'hBA98;
defparam \Mux26~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y31_N7
dffeas \registerArray[11][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][5] .is_wysiwyg = "true";
defparam \registerArray[11][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N6
cycloneive_lcell_comb \Mux26~13 (
// Equation(s):
// \Mux26~13_combout  = (\Mux26~12_combout  & (((\registerArray[11][5]~q ) # (!\my_rf.rsel1[0]~input_o )))) # (!\Mux26~12_combout  & (\registerArray[9][5]~q  & ((\my_rf.rsel1[0]~input_o ))))

	.dataa(\registerArray[9][5]~q ),
	.datab(\Mux26~12_combout ),
	.datac(\registerArray[11][5]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux26~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~13 .lut_mask = 16'hE2CC;
defparam \Mux26~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y31_N5
dffeas \registerArray[3][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][5] .is_wysiwyg = "true";
defparam \registerArray[3][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N15
dffeas \registerArray[1][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][5] .is_wysiwyg = "true";
defparam \registerArray[1][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N14
cycloneive_lcell_comb \Mux26~14 (
// Equation(s):
// \Mux26~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\registerArray[3][5]~q )) # (!\my_rf.rsel1[1]~input_o  & ((\registerArray[1][5]~q )))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\registerArray[3][5]~q ),
	.datac(\registerArray[1][5]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux26~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~14 .lut_mask = 16'h88A0;
defparam \Mux26~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N28
cycloneive_lcell_comb \Mux26~15 (
// Equation(s):
// \Mux26~15_combout  = (\Mux26~14_combout ) # ((!\my_rf.rsel1[0]~input_o  & (\registerArray[2][5]~q  & \my_rf.rsel1[1]~input_o )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux26~14_combout ),
	.datac(\registerArray[2][5]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux26~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~15 .lut_mask = 16'hDCCC;
defparam \Mux26~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N22
cycloneive_lcell_comb \Mux26~16 (
// Equation(s):
// \Mux26~16_combout  = (\my_rf.rsel1[2]~input_o  & (\my_rf.rsel1[3]~input_o )) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\Mux26~13_combout )) # (!\my_rf.rsel1[3]~input_o  & ((\Mux26~15_combout )))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\Mux26~13_combout ),
	.datad(\Mux26~15_combout ),
	.cin(gnd),
	.combout(\Mux26~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~16 .lut_mask = 16'hD9C8;
defparam \Mux26~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N0
cycloneive_lcell_comb \Mux26~17 (
// Equation(s):
// \Mux26~17_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[13][5]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[12][5]~q )))))

	.dataa(\registerArray[13][5]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[12][5]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux26~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~17 .lut_mask = 16'hEE30;
defparam \Mux26~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N23
dffeas \registerArray[15][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][5] .is_wysiwyg = "true";
defparam \registerArray[15][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N22
cycloneive_lcell_comb \Mux26~18 (
// Equation(s):
// \Mux26~18_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux26~17_combout  & (\registerArray[15][5]~q )) # (!\Mux26~17_combout  & ((\registerArray[14][5]~q ))))) # (!\my_rf.rsel1[1]~input_o  & (\Mux26~17_combout ))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\Mux26~17_combout ),
	.datac(\registerArray[15][5]~q ),
	.datad(\registerArray[14][5]~q ),
	.cin(gnd),
	.combout(\Mux26~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~18 .lut_mask = 16'hE6C4;
defparam \Mux26~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N24
cycloneive_lcell_comb \Mux26~19 (
// Equation(s):
// \Mux26~19_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux26~16_combout  & ((\Mux26~18_combout ))) # (!\Mux26~16_combout  & (\Mux26~11_combout )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux26~16_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux26~11_combout ),
	.datac(\Mux26~16_combout ),
	.datad(\Mux26~18_combout ),
	.cin(gnd),
	.combout(\Mux26~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~19 .lut_mask = 16'hF858;
defparam \Mux26~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y34_N27
dffeas \registerArray[17][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][5] .is_wysiwyg = "true";
defparam \registerArray[17][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N26
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[25][5]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[17][5]~q )))))

	.dataa(\registerArray[25][5]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[17][5]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hEE30;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N12
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// \Mux26~1_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux26~0_combout  & ((\registerArray[29][5]~q ))) # (!\Mux26~0_combout  & (\registerArray[21][5]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux26~0_combout ))))

	.dataa(\registerArray[21][5]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[29][5]~q ),
	.datad(\Mux26~0_combout ),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hF388;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N7
dffeas \registerArray[28][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][5] .is_wysiwyg = "true";
defparam \registerArray[28][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N18
cycloneive_lcell_comb \Mux26~4 (
// Equation(s):
// \Mux26~4_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[20][5]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[16][5]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[16][5]~q ),
	.datad(\registerArray[20][5]~q ),
	.cin(gnd),
	.combout(\Mux26~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~4 .lut_mask = 16'hDC98;
defparam \Mux26~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N6
cycloneive_lcell_comb \Mux26~5 (
// Equation(s):
// \Mux26~5_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux26~4_combout  & ((\registerArray[28][5]~q ))) # (!\Mux26~4_combout  & (\registerArray[24][5]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux26~4_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[24][5]~q ),
	.datac(\registerArray[28][5]~q ),
	.datad(\Mux26~4_combout ),
	.cin(gnd),
	.combout(\Mux26~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~5 .lut_mask = 16'hF588;
defparam \Mux26~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N8
cycloneive_lcell_comb \Mux26~3 (
// Equation(s):
// \Mux26~3_combout  = (\Mux26~2_combout  & (((\registerArray[30][5]~q )) # (!\my_rf.rsel1[3]~input_o ))) # (!\Mux26~2_combout  & (\my_rf.rsel1[3]~input_o  & ((\registerArray[26][5]~q ))))

	.dataa(\Mux26~2_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[30][5]~q ),
	.datad(\registerArray[26][5]~q ),
	.cin(gnd),
	.combout(\Mux26~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~3 .lut_mask = 16'hE6A2;
defparam \Mux26~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N8
cycloneive_lcell_comb \Mux26~6 (
// Equation(s):
// \Mux26~6_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\Mux26~3_combout ))) # (!\my_rf.rsel1[1]~input_o  & (\Mux26~5_combout ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux26~5_combout ),
	.datac(\Mux26~3_combout ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux26~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~6 .lut_mask = 16'hFA44;
defparam \Mux26~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y32_N15
dffeas \registerArray[31][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][5] .is_wysiwyg = "true";
defparam \registerArray[31][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N13
dffeas \registerArray[19][5] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[5]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][5] .is_wysiwyg = "true";
defparam \registerArray[19][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N12
cycloneive_lcell_comb \Mux26~7 (
// Equation(s):
// \Mux26~7_combout  = (\my_rf.rsel1[2]~input_o  & (\my_rf.rsel1[3]~input_o )) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & ((\registerArray[27][5]~q ))) # (!\my_rf.rsel1[3]~input_o  & (\registerArray[19][5]~q ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[19][5]~q ),
	.datad(\registerArray[27][5]~q ),
	.cin(gnd),
	.combout(\Mux26~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~7 .lut_mask = 16'hDC98;
defparam \Mux26~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N14
cycloneive_lcell_comb \Mux26~8 (
// Equation(s):
// \Mux26~8_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux26~7_combout  & ((\registerArray[31][5]~q ))) # (!\Mux26~7_combout  & (\registerArray[23][5]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux26~7_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[23][5]~q ),
	.datac(\registerArray[31][5]~q ),
	.datad(\Mux26~7_combout ),
	.cin(gnd),
	.combout(\Mux26~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~8 .lut_mask = 16'hF588;
defparam \Mux26~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N10
cycloneive_lcell_comb \Mux26~9 (
// Equation(s):
// \Mux26~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux26~6_combout  & ((\Mux26~8_combout ))) # (!\Mux26~6_combout  & (\Mux26~1_combout )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux26~6_combout ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux26~1_combout ),
	.datac(\Mux26~6_combout ),
	.datad(\Mux26~8_combout ),
	.cin(gnd),
	.combout(\Mux26~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~9 .lut_mask = 16'hF858;
defparam \Mux26~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N2
cycloneive_lcell_comb \Mux26~20 (
// Equation(s):
// \Mux26~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux26~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux26~19_combout ))

	.dataa(gnd),
	.datab(\Mux26~19_combout ),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux26~9_combout ),
	.cin(gnd),
	.combout(\Mux26~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~20 .lut_mask = 16'hFC0C;
defparam \Mux26~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y31_N27
dffeas \registerArray[11][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][6] .is_wysiwyg = "true";
defparam \registerArray[11][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y31_N18
cycloneive_lcell_comb \Mux25~10 (
// Equation(s):
// \Mux25~10_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\registerArray[10][6]~q )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & (\registerArray[8][6]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[8][6]~q ),
	.datad(\registerArray[10][6]~q ),
	.cin(gnd),
	.combout(\Mux25~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~10 .lut_mask = 16'hBA98;
defparam \Mux25~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N26
cycloneive_lcell_comb \Mux25~11 (
// Equation(s):
// \Mux25~11_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux25~10_combout  & ((\registerArray[11][6]~q ))) # (!\Mux25~10_combout  & (\registerArray[9][6]~q )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux25~10_combout ))))

	.dataa(\registerArray[9][6]~q ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[11][6]~q ),
	.datad(\Mux25~10_combout ),
	.cin(gnd),
	.combout(\Mux25~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~11 .lut_mask = 16'hF388;
defparam \Mux25~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N19
dffeas \registerArray[12][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][6] .is_wysiwyg = "true";
defparam \registerArray[12][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N25
dffeas \registerArray[13][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][6] .is_wysiwyg = "true";
defparam \registerArray[13][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N18
cycloneive_lcell_comb \Mux25~17 (
// Equation(s):
// \Mux25~17_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[13][6]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[12][6]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][6]~q ),
	.datad(\registerArray[13][6]~q ),
	.cin(gnd),
	.combout(\Mux25~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~17 .lut_mask = 16'hDC98;
defparam \Mux25~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N9
dffeas \registerArray[15][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][6] .is_wysiwyg = "true";
defparam \registerArray[15][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N13
dffeas \registerArray[14][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][6] .is_wysiwyg = "true";
defparam \registerArray[14][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N8
cycloneive_lcell_comb \Mux25~18 (
// Equation(s):
// \Mux25~18_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux25~17_combout  & (\registerArray[15][6]~q )) # (!\Mux25~17_combout  & ((\registerArray[14][6]~q ))))) # (!\my_rf.rsel1[1]~input_o  & (\Mux25~17_combout ))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\Mux25~17_combout ),
	.datac(\registerArray[15][6]~q ),
	.datad(\registerArray[14][6]~q ),
	.cin(gnd),
	.combout(\Mux25~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~18 .lut_mask = 16'hE6C4;
defparam \Mux25~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N8
cycloneive_lcell_comb \Mux25~19 (
// Equation(s):
// \Mux25~19_combout  = (\Mux25~16_combout  & (((\Mux25~18_combout ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux25~16_combout  & (\Mux25~11_combout  & (\my_rf.rsel1[3]~input_o )))

	.dataa(\Mux25~16_combout ),
	.datab(\Mux25~11_combout ),
	.datac(\my_rf.rsel1[3]~input_o ),
	.datad(\Mux25~18_combout ),
	.cin(gnd),
	.combout(\Mux25~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~19 .lut_mask = 16'hEA4A;
defparam \Mux25~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y0_N3
dffeas \registerArray[25][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[6]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][6] .is_wysiwyg = "true";
defparam \registerArray[25][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y36_N31
dffeas \registerArray[29][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][6] .is_wysiwyg = "true";
defparam \registerArray[29][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N31
dffeas \registerArray[17][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][6] .is_wysiwyg = "true";
defparam \registerArray[17][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N29
dffeas \registerArray[21][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][6] .is_wysiwyg = "true";
defparam \registerArray[21][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N30
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o ) # ((\registerArray[21][6]~q )))) # (!\my_rf.rsel1[2]~input_o  & (!\my_rf.rsel1[3]~input_o  & (\registerArray[17][6]~q )))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[17][6]~q ),
	.datad(\registerArray[21][6]~q ),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hBA98;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N30
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// \Mux25~1_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux25~0_combout  & ((\registerArray[29][6]~q ))) # (!\Mux25~0_combout  & (\registerArray[25][6]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux25~0_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[25][6]~q ),
	.datac(\registerArray[29][6]~q ),
	.datad(\Mux25~0_combout ),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hF588;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N25
dffeas \registerArray[22][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][6] .is_wysiwyg = "true";
defparam \registerArray[22][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y36_N19
dffeas \registerArray[30][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][6] .is_wysiwyg = "true";
defparam \registerArray[30][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y36_N3
dffeas \registerArray[18][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][6] .is_wysiwyg = "true";
defparam \registerArray[18][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y36_N9
dffeas \registerArray[26][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][6] .is_wysiwyg = "true";
defparam \registerArray[26][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N2
cycloneive_lcell_comb \Mux25~2 (
// Equation(s):
// \Mux25~2_combout  = (\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o ) # ((\registerArray[26][6]~q )))) # (!\my_rf.rsel1[3]~input_o  & (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][6]~q )))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][6]~q ),
	.datad(\registerArray[26][6]~q ),
	.cin(gnd),
	.combout(\Mux25~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~2 .lut_mask = 16'hBA98;
defparam \Mux25~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N18
cycloneive_lcell_comb \Mux25~3 (
// Equation(s):
// \Mux25~3_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux25~2_combout  & ((\registerArray[30][6]~q ))) # (!\Mux25~2_combout  & (\registerArray[22][6]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux25~2_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[22][6]~q ),
	.datac(\registerArray[30][6]~q ),
	.datad(\Mux25~2_combout ),
	.cin(gnd),
	.combout(\Mux25~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~3 .lut_mask = 16'hF588;
defparam \Mux25~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y36_N15
dffeas \registerArray[16][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][6] .is_wysiwyg = "true";
defparam \registerArray[16][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N14
cycloneive_lcell_comb \Mux25~4 (
// Equation(s):
// \Mux25~4_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[24][6]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[16][6]~q )))))

	.dataa(\registerArray[24][6]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[16][6]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux25~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~4 .lut_mask = 16'hEE30;
defparam \Mux25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N3
dffeas \registerArray[28][6] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[6]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][6] .is_wysiwyg = "true";
defparam \registerArray[28][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N2
cycloneive_lcell_comb \Mux25~5 (
// Equation(s):
// \Mux25~5_combout  = (\Mux25~4_combout  & (((\registerArray[28][6]~q ) # (!\my_rf.rsel1[2]~input_o )))) # (!\Mux25~4_combout  & (\registerArray[20][6]~q  & ((\my_rf.rsel1[2]~input_o ))))

	.dataa(\registerArray[20][6]~q ),
	.datab(\Mux25~4_combout ),
	.datac(\registerArray[28][6]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux25~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~5 .lut_mask = 16'hE2CC;
defparam \Mux25~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N16
cycloneive_lcell_comb \Mux25~6 (
// Equation(s):
// \Mux25~6_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\Mux25~3_combout )) # (!\my_rf.rsel1[1]~input_o  & ((\Mux25~5_combout )))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux25~3_combout ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\Mux25~5_combout ),
	.cin(gnd),
	.combout(\Mux25~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~6 .lut_mask = 16'hE5E0;
defparam \Mux25~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N2
cycloneive_lcell_comb \Mux25~9 (
// Equation(s):
// \Mux25~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux25~6_combout  & (\Mux25~8_combout )) # (!\Mux25~6_combout  & ((\Mux25~1_combout ))))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux25~6_combout ))))

	.dataa(\Mux25~8_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux25~1_combout ),
	.datad(\Mux25~6_combout ),
	.cin(gnd),
	.combout(\Mux25~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~9 .lut_mask = 16'hBBC0;
defparam \Mux25~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N10
cycloneive_lcell_comb \Mux25~20 (
// Equation(s):
// \Mux25~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux25~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux25~19_combout ))

	.dataa(gnd),
	.datab(\Mux25~19_combout ),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux25~9_combout ),
	.cin(gnd),
	.combout(\Mux25~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~20 .lut_mask = 16'hFC0C;
defparam \Mux25~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N25
dffeas \registerArray[29][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][7] .is_wysiwyg = "true";
defparam \registerArray[29][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y0_N10
dffeas \registerArray[21][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[7]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][7] .is_wysiwyg = "true";
defparam \registerArray[21][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N24
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// \Mux24~1_combout  = (\Mux24~0_combout  & (((\registerArray[29][7]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux24~0_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[21][7]~q ))))

	.dataa(\Mux24~0_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[29][7]~q ),
	.datad(\registerArray[21][7]~q ),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'hE6A2;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N9
dffeas \registerArray[27][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][7] .is_wysiwyg = "true";
defparam \registerArray[27][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N3
dffeas \registerArray[19][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][7] .is_wysiwyg = "true";
defparam \registerArray[19][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N2
cycloneive_lcell_comb \Mux24~7 (
// Equation(s):
// \Mux24~7_combout  = (\my_rf.rsel1[3]~input_o  & ((\registerArray[27][7]~q ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((\registerArray[19][7]~q  & !\my_rf.rsel1[2]~input_o ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[27][7]~q ),
	.datac(\registerArray[19][7]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux24~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~7 .lut_mask = 16'hAAD8;
defparam \Mux24~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N18
cycloneive_lcell_comb \Mux24~8 (
// Equation(s):
// \Mux24~8_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux24~7_combout  & (\registerArray[31][7]~q )) # (!\Mux24~7_combout  & ((\registerArray[23][7]~q ))))) # (!\my_rf.rsel1[2]~input_o  & (\Mux24~7_combout ))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux24~7_combout ),
	.datac(\registerArray[31][7]~q ),
	.datad(\registerArray[23][7]~q ),
	.cin(gnd),
	.combout(\Mux24~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~8 .lut_mask = 16'hE6C4;
defparam \Mux24~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N30
cycloneive_lcell_comb \Mux24~9 (
// Equation(s):
// \Mux24~9_combout  = (\Mux24~6_combout  & (((\Mux24~8_combout ) # (!\my_rf.rsel1[0]~input_o )))) # (!\Mux24~6_combout  & (\Mux24~1_combout  & ((\my_rf.rsel1[0]~input_o ))))

	.dataa(\Mux24~6_combout ),
	.datab(\Mux24~1_combout ),
	.datac(\Mux24~8_combout ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux24~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~9 .lut_mask = 16'hE4AA;
defparam \Mux24~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y29_N11
dffeas \registerArray[7][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][7] .is_wysiwyg = "true";
defparam \registerArray[7][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N10
cycloneive_lcell_comb \Mux24~11 (
// Equation(s):
// \Mux24~11_combout  = (\Mux24~10_combout  & (((\registerArray[7][7]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux24~10_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[6][7]~q ))))

	.dataa(\Mux24~10_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[7][7]~q ),
	.datad(\registerArray[6][7]~q ),
	.cin(gnd),
	.combout(\Mux24~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~11 .lut_mask = 16'hE6A2;
defparam \Mux24~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N26
cycloneive_lcell_comb \Mux24~14 (
// Equation(s):
// \Mux24~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][7]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][7]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[1][7]~q ),
	.datad(\registerArray[3][7]~q ),
	.cin(gnd),
	.combout(\Mux24~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~14 .lut_mask = 16'hC840;
defparam \Mux24~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N8
cycloneive_lcell_comb \Mux24~15 (
// Equation(s):
// \Mux24~15_combout  = (\Mux24~14_combout ) # ((\my_rf.rsel1[1]~input_o  & (\registerArray[2][7]~q  & !\my_rf.rsel1[0]~input_o )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[2][7]~q ),
	.datac(\Mux24~14_combout ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux24~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~15 .lut_mask = 16'hF0F8;
defparam \Mux24~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y31_N15
dffeas \registerArray[11][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][7] .is_wysiwyg = "true";
defparam \registerArray[11][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y31_N29
dffeas \registerArray[9][7] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[7]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][7] .is_wysiwyg = "true";
defparam \registerArray[9][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N14
cycloneive_lcell_comb \Mux24~13 (
// Equation(s):
// \Mux24~13_combout  = (\Mux24~12_combout  & (((\registerArray[11][7]~q )) # (!\my_rf.rsel1[0]~input_o ))) # (!\Mux24~12_combout  & (\my_rf.rsel1[0]~input_o  & ((\registerArray[9][7]~q ))))

	.dataa(\Mux24~12_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[11][7]~q ),
	.datad(\registerArray[9][7]~q ),
	.cin(gnd),
	.combout(\Mux24~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~13 .lut_mask = 16'hE6A2;
defparam \Mux24~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N10
cycloneive_lcell_comb \Mux24~16 (
// Equation(s):
// \Mux24~16_combout  = (\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o ) # ((\Mux24~13_combout )))) # (!\my_rf.rsel1[3]~input_o  & (!\my_rf.rsel1[2]~input_o  & (\Mux24~15_combout )))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux24~15_combout ),
	.datad(\Mux24~13_combout ),
	.cin(gnd),
	.combout(\Mux24~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~16 .lut_mask = 16'hBA98;
defparam \Mux24~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N12
cycloneive_lcell_comb \Mux24~19 (
// Equation(s):
// \Mux24~19_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux24~16_combout  & (\Mux24~18_combout )) # (!\Mux24~16_combout  & ((\Mux24~11_combout ))))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux24~16_combout ))))

	.dataa(\Mux24~18_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux24~11_combout ),
	.datad(\Mux24~16_combout ),
	.cin(gnd),
	.combout(\Mux24~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~19 .lut_mask = 16'hBBC0;
defparam \Mux24~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N14
cycloneive_lcell_comb \Mux24~20 (
// Equation(s):
// \Mux24~20_combout  = (\my_rf.rsel1[4]~input_o  & (\Mux24~9_combout )) # (!\my_rf.rsel1[4]~input_o  & ((\Mux24~19_combout )))

	.dataa(\my_rf.rsel1[4]~input_o ),
	.datab(gnd),
	.datac(\Mux24~9_combout ),
	.datad(\Mux24~19_combout ),
	.cin(gnd),
	.combout(\Mux24~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~20 .lut_mask = 16'hF5A0;
defparam \Mux24~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y33_N7
dffeas \registerArray[31][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][8] .is_wysiwyg = "true";
defparam \registerArray[31][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y33_N21
dffeas \registerArray[19][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][8] .is_wysiwyg = "true";
defparam \registerArray[19][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N20
cycloneive_lcell_comb \Mux23~7 (
// Equation(s):
// \Mux23~7_combout  = (\my_rf.rsel1[2]~input_o  & ((\registerArray[23][8]~q ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\registerArray[19][8]~q  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\registerArray[23][8]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[19][8]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux23~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~7 .lut_mask = 16'hCCB8;
defparam \Mux23~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N6
cycloneive_lcell_comb \Mux23~8 (
// Equation(s):
// \Mux23~8_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux23~7_combout  & ((\registerArray[31][8]~q ))) # (!\Mux23~7_combout  & (\registerArray[27][8]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux23~7_combout ))))

	.dataa(\registerArray[27][8]~q ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[31][8]~q ),
	.datad(\Mux23~7_combout ),
	.cin(gnd),
	.combout(\Mux23~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~8 .lut_mask = 16'hF388;
defparam \Mux23~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N10
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// \Mux23~0_combout  = (\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o ) # ((\registerArray[21][8]~q )))) # (!\my_rf.rsel1[2]~input_o  & (!\my_rf.rsel1[3]~input_o  & (\registerArray[17][8]~q )))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[17][8]~q ),
	.datad(\registerArray[21][8]~q ),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hBA98;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N26
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// \Mux23~1_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux23~0_combout  & (\registerArray[29][8]~q )) # (!\Mux23~0_combout  & ((\registerArray[25][8]~q ))))) # (!\my_rf.rsel1[3]~input_o  & (\Mux23~0_combout ))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux23~0_combout ),
	.datac(\registerArray[29][8]~q ),
	.datad(\registerArray[25][8]~q ),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'hE6C4;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y37_N3
dffeas \registerArray[16][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][8] .is_wysiwyg = "true";
defparam \registerArray[16][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N1
dffeas \registerArray[24][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][8] .is_wysiwyg = "true";
defparam \registerArray[24][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N2
cycloneive_lcell_comb \Mux23~4 (
// Equation(s):
// \Mux23~4_combout  = (\my_rf.rsel1[2]~input_o  & (\my_rf.rsel1[3]~input_o )) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & ((\registerArray[24][8]~q ))) # (!\my_rf.rsel1[3]~input_o  & (\registerArray[16][8]~q ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[16][8]~q ),
	.datad(\registerArray[24][8]~q ),
	.cin(gnd),
	.combout(\Mux23~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~4 .lut_mask = 16'hDC98;
defparam \Mux23~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N2
cycloneive_lcell_comb \Mux23~5 (
// Equation(s):
// \Mux23~5_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux23~4_combout  & ((\registerArray[28][8]~q ))) # (!\Mux23~4_combout  & (\registerArray[20][8]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux23~4_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[20][8]~q ),
	.datac(\registerArray[28][8]~q ),
	.datad(\Mux23~4_combout ),
	.cin(gnd),
	.combout(\Mux23~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~5 .lut_mask = 16'hF588;
defparam \Mux23~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y36_N19
dffeas \registerArray[18][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][8] .is_wysiwyg = "true";
defparam \registerArray[18][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y36_N17
dffeas \registerArray[26][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][8] .is_wysiwyg = "true";
defparam \registerArray[26][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y36_N18
cycloneive_lcell_comb \Mux23~2 (
// Equation(s):
// \Mux23~2_combout  = (\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o ) # ((\registerArray[26][8]~q )))) # (!\my_rf.rsel1[3]~input_o  & (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][8]~q )))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][8]~q ),
	.datad(\registerArray[26][8]~q ),
	.cin(gnd),
	.combout(\Mux23~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~2 .lut_mask = 16'hBA98;
defparam \Mux23~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N26
cycloneive_lcell_comb \Mux23~3 (
// Equation(s):
// \Mux23~3_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux23~2_combout  & ((\registerArray[30][8]~q ))) # (!\Mux23~2_combout  & (\registerArray[22][8]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux23~2_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[22][8]~q ),
	.datac(\registerArray[30][8]~q ),
	.datad(\Mux23~2_combout ),
	.cin(gnd),
	.combout(\Mux23~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~3 .lut_mask = 16'hF588;
defparam \Mux23~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N12
cycloneive_lcell_comb \Mux23~6 (
// Equation(s):
// \Mux23~6_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\Mux23~3_combout ))) # (!\my_rf.rsel1[1]~input_o  & (\Mux23~5_combout ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux23~5_combout ),
	.datac(\Mux23~3_combout ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux23~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~6 .lut_mask = 16'hFA44;
defparam \Mux23~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N6
cycloneive_lcell_comb \Mux23~9 (
// Equation(s):
// \Mux23~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux23~6_combout  & (\Mux23~8_combout )) # (!\Mux23~6_combout  & ((\Mux23~1_combout ))))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux23~6_combout ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux23~8_combout ),
	.datac(\Mux23~1_combout ),
	.datad(\Mux23~6_combout ),
	.cin(gnd),
	.combout(\Mux23~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~9 .lut_mask = 16'hDDA0;
defparam \Mux23~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y37_N27
dffeas \registerArray[11][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][8] .is_wysiwyg = "true";
defparam \registerArray[11][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y37_N26
cycloneive_lcell_comb \Mux23~11 (
// Equation(s):
// \Mux23~11_combout  = (\Mux23~10_combout  & (((\registerArray[11][8]~q )) # (!\my_rf.rsel1[0]~input_o ))) # (!\Mux23~10_combout  & (\my_rf.rsel1[0]~input_o  & ((\registerArray[9][8]~q ))))

	.dataa(\Mux23~10_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[11][8]~q ),
	.datad(\registerArray[9][8]~q ),
	.cin(gnd),
	.combout(\Mux23~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~11 .lut_mask = 16'hE6A2;
defparam \Mux23~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N28
cycloneive_lcell_comb \Mux23~13 (
// Equation(s):
// \Mux23~13_combout  = (\Mux23~12_combout  & (((\registerArray[7][8]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux23~12_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[6][8]~q ))))

	.dataa(\Mux23~12_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[7][8]~q ),
	.datad(\registerArray[6][8]~q ),
	.cin(gnd),
	.combout(\Mux23~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~13 .lut_mask = 16'hE6A2;
defparam \Mux23~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N5
dffeas \registerArray[3][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][8] .is_wysiwyg = "true";
defparam \registerArray[3][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N23
dffeas \registerArray[1][8] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[8]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][8] .is_wysiwyg = "true";
defparam \registerArray[1][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N22
cycloneive_lcell_comb \Mux23~14 (
// Equation(s):
// \Mux23~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\registerArray[3][8]~q )) # (!\my_rf.rsel1[1]~input_o  & ((\registerArray[1][8]~q )))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[3][8]~q ),
	.datac(\registerArray[1][8]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux23~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~14 .lut_mask = 16'hD800;
defparam \Mux23~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N24
cycloneive_lcell_comb \Mux23~15 (
// Equation(s):
// \Mux23~15_combout  = (\Mux23~14_combout ) # ((\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & \registerArray[2][8]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux23~14_combout ),
	.datad(\registerArray[2][8]~q ),
	.cin(gnd),
	.combout(\Mux23~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~15 .lut_mask = 16'hF2F0;
defparam \Mux23~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N2
cycloneive_lcell_comb \Mux23~16 (
// Equation(s):
// \Mux23~16_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & (\Mux23~13_combout )) # (!\my_rf.rsel1[2]~input_o  & ((\Mux23~15_combout )))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux23~13_combout ),
	.datad(\Mux23~15_combout ),
	.cin(gnd),
	.combout(\Mux23~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~16 .lut_mask = 16'hD9C8;
defparam \Mux23~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N28
cycloneive_lcell_comb \Mux23~19 (
// Equation(s):
// \Mux23~19_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux23~16_combout  & (\Mux23~18_combout )) # (!\Mux23~16_combout  & ((\Mux23~11_combout ))))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux23~16_combout ))))

	.dataa(\Mux23~18_combout ),
	.datab(\Mux23~11_combout ),
	.datac(\my_rf.rsel1[3]~input_o ),
	.datad(\Mux23~16_combout ),
	.cin(gnd),
	.combout(\Mux23~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~19 .lut_mask = 16'hAFC0;
defparam \Mux23~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N16
cycloneive_lcell_comb \Mux23~20 (
// Equation(s):
// \Mux23~20_combout  = (\my_rf.rsel1[4]~input_o  & (\Mux23~9_combout )) # (!\my_rf.rsel1[4]~input_o  & ((\Mux23~19_combout )))

	.dataa(\Mux23~9_combout ),
	.datab(gnd),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux23~19_combout ),
	.cin(gnd),
	.combout(\Mux23~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~20 .lut_mask = 16'hAFA0;
defparam \Mux23~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y36_N9
dffeas \registerArray[3][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][9] .is_wysiwyg = "true";
defparam \registerArray[3][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N11
dffeas \registerArray[1][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][9] .is_wysiwyg = "true";
defparam \registerArray[1][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N10
cycloneive_lcell_comb \Mux22~14 (
// Equation(s):
// \Mux22~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\registerArray[3][9]~q )) # (!\my_rf.rsel1[1]~input_o  & ((\registerArray[1][9]~q )))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[3][9]~q ),
	.datac(\registerArray[1][9]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux22~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~14 .lut_mask = 16'hD800;
defparam \Mux22~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N12
cycloneive_lcell_comb \Mux22~15 (
// Equation(s):
// \Mux22~15_combout  = (\Mux22~14_combout ) # ((\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & \registerArray[2][9]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux22~14_combout ),
	.datad(\registerArray[2][9]~q ),
	.cin(gnd),
	.combout(\Mux22~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~15 .lut_mask = 16'hF2F0;
defparam \Mux22~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N14
cycloneive_lcell_comb \Mux22~16 (
// Equation(s):
// \Mux22~16_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux22~13_combout ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((!\my_rf.rsel1[2]~input_o  & \Mux22~15_combout ))))

	.dataa(\Mux22~13_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux22~15_combout ),
	.cin(gnd),
	.combout(\Mux22~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~16 .lut_mask = 16'hCBC8;
defparam \Mux22~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N22
cycloneive_lcell_comb \Mux22~11 (
// Equation(s):
// \Mux22~11_combout  = (\Mux22~10_combout  & (((\registerArray[7][9]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux22~10_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[6][9]~q ))))

	.dataa(\Mux22~10_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[7][9]~q ),
	.datad(\registerArray[6][9]~q ),
	.cin(gnd),
	.combout(\Mux22~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~11 .lut_mask = 16'hE6A2;
defparam \Mux22~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N0
cycloneive_lcell_comb \Mux22~19 (
// Equation(s):
// \Mux22~19_combout  = (\Mux22~16_combout  & ((\Mux22~18_combout ) # ((!\my_rf.rsel1[2]~input_o )))) # (!\Mux22~16_combout  & (((\my_rf.rsel1[2]~input_o  & \Mux22~11_combout ))))

	.dataa(\Mux22~18_combout ),
	.datab(\Mux22~16_combout ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux22~11_combout ),
	.cin(gnd),
	.combout(\Mux22~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~19 .lut_mask = 16'hBC8C;
defparam \Mux22~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y33_N11
dffeas \registerArray[31][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][9] .is_wysiwyg = "true";
defparam \registerArray[31][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N10
cycloneive_lcell_comb \Mux22~8 (
// Equation(s):
// \Mux22~8_combout  = (\Mux22~7_combout  & (((\registerArray[31][9]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux22~7_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[23][9]~q ))))

	.dataa(\Mux22~7_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[31][9]~q ),
	.datad(\registerArray[23][9]~q ),
	.cin(gnd),
	.combout(\Mux22~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~8 .lut_mask = 16'hE6A2;
defparam \Mux22~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N13
dffeas \registerArray[25][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][9] .is_wysiwyg = "true";
defparam \registerArray[25][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y34_N13
dffeas \registerArray[17][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][9] .is_wysiwyg = "true";
defparam \registerArray[17][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y34_N12
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// \Mux22~0_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[25][9]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[17][9]~q )))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[25][9]~q ),
	.datac(\registerArray[17][9]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'hEE50;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N22
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// \Mux22~1_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux22~0_combout  & ((\registerArray[29][9]~q ))) # (!\Mux22~0_combout  & (\registerArray[21][9]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux22~0_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[21][9]~q ),
	.datac(\registerArray[29][9]~q ),
	.datad(\Mux22~0_combout ),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'hF588;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y36_N31
dffeas \registerArray[30][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][9] .is_wysiwyg = "true";
defparam \registerArray[30][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N2
cycloneive_lcell_comb \Mux22~2 (
// Equation(s):
// \Mux22~2_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[22][9]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][9]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][9]~q ),
	.datad(\registerArray[22][9]~q ),
	.cin(gnd),
	.combout(\Mux22~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~2 .lut_mask = 16'hDC98;
defparam \Mux22~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N30
cycloneive_lcell_comb \Mux22~3 (
// Equation(s):
// \Mux22~3_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux22~2_combout  & ((\registerArray[30][9]~q ))) # (!\Mux22~2_combout  & (\registerArray[26][9]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux22~2_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[26][9]~q ),
	.datac(\registerArray[30][9]~q ),
	.datad(\Mux22~2_combout ),
	.cin(gnd),
	.combout(\Mux22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~3 .lut_mask = 16'hF588;
defparam \Mux22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y36_N23
dffeas \registerArray[16][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][9] .is_wysiwyg = "true";
defparam \registerArray[16][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N22
cycloneive_lcell_comb \Mux22~4 (
// Equation(s):
// \Mux22~4_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[20][9]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[16][9]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[16][9]~q ),
	.datad(\registerArray[20][9]~q ),
	.cin(gnd),
	.combout(\Mux22~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~4 .lut_mask = 16'hDC98;
defparam \Mux22~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N5
dffeas \registerArray[28][9] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[9]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][9] .is_wysiwyg = "true";
defparam \registerArray[28][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N4
cycloneive_lcell_comb \Mux22~5 (
// Equation(s):
// \Mux22~5_combout  = (\Mux22~4_combout  & (((\registerArray[28][9]~q ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux22~4_combout  & (\registerArray[24][9]~q  & ((\my_rf.rsel1[3]~input_o ))))

	.dataa(\registerArray[24][9]~q ),
	.datab(\Mux22~4_combout ),
	.datac(\registerArray[28][9]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux22~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~5 .lut_mask = 16'hE2CC;
defparam \Mux22~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N18
cycloneive_lcell_comb \Mux22~6 (
// Equation(s):
// \Mux22~6_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\Mux22~3_combout )) # (!\my_rf.rsel1[1]~input_o  & ((\Mux22~5_combout )))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux22~3_combout ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\Mux22~5_combout ),
	.cin(gnd),
	.combout(\Mux22~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~6 .lut_mask = 16'hE5E0;
defparam \Mux22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N20
cycloneive_lcell_comb \Mux22~9 (
// Equation(s):
// \Mux22~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux22~6_combout  & (\Mux22~8_combout )) # (!\Mux22~6_combout  & ((\Mux22~1_combout ))))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux22~6_combout ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux22~8_combout ),
	.datac(\Mux22~1_combout ),
	.datad(\Mux22~6_combout ),
	.cin(gnd),
	.combout(\Mux22~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~9 .lut_mask = 16'hDDA0;
defparam \Mux22~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N26
cycloneive_lcell_comb \Mux22~20 (
// Equation(s):
// \Mux22~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux22~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux22~19_combout ))

	.dataa(gnd),
	.datab(\Mux22~19_combout ),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux22~9_combout ),
	.cin(gnd),
	.combout(\Mux22~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~20 .lut_mask = 16'hFC0C;
defparam \Mux22~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N23
dffeas \registerArray[12][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][10] .is_wysiwyg = "true";
defparam \registerArray[12][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N22
cycloneive_lcell_comb \Mux21~17 (
// Equation(s):
// \Mux21~17_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o ) # ((\registerArray[13][10]~q )))) # (!\my_rf.rsel1[0]~input_o  & (!\my_rf.rsel1[1]~input_o  & (\registerArray[12][10]~q )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[12][10]~q ),
	.datad(\registerArray[13][10]~q ),
	.cin(gnd),
	.combout(\Mux21~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~17 .lut_mask = 16'hBA98;
defparam \Mux21~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N14
cycloneive_lcell_comb \Mux21~18 (
// Equation(s):
// \Mux21~18_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux21~17_combout  & ((\registerArray[15][10]~q ))) # (!\Mux21~17_combout  & (\registerArray[14][10]~q )))) # (!\my_rf.rsel1[1]~input_o  & (((\Mux21~17_combout ))))

	.dataa(\registerArray[14][10]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][10]~q ),
	.datad(\Mux21~17_combout ),
	.cin(gnd),
	.combout(\Mux21~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~18 .lut_mask = 16'hF388;
defparam \Mux21~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N6
cycloneive_lcell_comb \Mux21~14 (
// Equation(s):
// \Mux21~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][10]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][10]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[1][10]~q ),
	.datad(\registerArray[3][10]~q ),
	.cin(gnd),
	.combout(\Mux21~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~14 .lut_mask = 16'hC840;
defparam \Mux21~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N24
cycloneive_lcell_comb \Mux21~15 (
// Equation(s):
// \Mux21~15_combout  = (\Mux21~14_combout ) # ((\registerArray[2][10]~q  & (\my_rf.rsel1[1]~input_o  & !\my_rf.rsel1[0]~input_o )))

	.dataa(\registerArray[2][10]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\Mux21~14_combout ),
	.cin(gnd),
	.combout(\Mux21~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~15 .lut_mask = 16'hFF08;
defparam \Mux21~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N10
cycloneive_lcell_comb \Mux21~13 (
// Equation(s):
// \Mux21~13_combout  = (\Mux21~12_combout  & (((\registerArray[7][10]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux21~12_combout  & (\registerArray[6][10]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux21~12_combout ),
	.datab(\registerArray[6][10]~q ),
	.datac(\registerArray[7][10]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux21~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~13 .lut_mask = 16'hE4AA;
defparam \Mux21~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N26
cycloneive_lcell_comb \Mux21~16 (
// Equation(s):
// \Mux21~16_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\Mux21~13_combout ))) # (!\my_rf.rsel1[2]~input_o  & (\Mux21~15_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux21~15_combout ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux21~13_combout ),
	.cin(gnd),
	.combout(\Mux21~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~16 .lut_mask = 16'hF4A4;
defparam \Mux21~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y37_N9
dffeas \registerArray[9][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][10] .is_wysiwyg = "true";
defparam \registerArray[9][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y37_N3
dffeas \registerArray[11][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][10] .is_wysiwyg = "true";
defparam \registerArray[11][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y37_N2
cycloneive_lcell_comb \Mux21~11 (
// Equation(s):
// \Mux21~11_combout  = (\Mux21~10_combout  & (((\registerArray[11][10]~q ) # (!\my_rf.rsel1[0]~input_o )))) # (!\Mux21~10_combout  & (\registerArray[9][10]~q  & ((\my_rf.rsel1[0]~input_o ))))

	.dataa(\Mux21~10_combout ),
	.datab(\registerArray[9][10]~q ),
	.datac(\registerArray[11][10]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux21~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~11 .lut_mask = 16'hE4AA;
defparam \Mux21~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N28
cycloneive_lcell_comb \Mux21~19 (
// Equation(s):
// \Mux21~19_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux21~16_combout  & (\Mux21~18_combout )) # (!\Mux21~16_combout  & ((\Mux21~11_combout ))))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux21~16_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux21~18_combout ),
	.datac(\Mux21~16_combout ),
	.datad(\Mux21~11_combout ),
	.cin(gnd),
	.combout(\Mux21~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~19 .lut_mask = 16'hDAD0;
defparam \Mux21~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N22
cycloneive_lcell_comb \Mux21~7 (
// Equation(s):
// \Mux21~7_combout  = (\my_rf.rsel1[2]~input_o  & ((\registerArray[23][10]~q ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\registerArray[19][10]~q  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[23][10]~q ),
	.datac(\registerArray[19][10]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux21~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~7 .lut_mask = 16'hAAD8;
defparam \Mux21~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N22
cycloneive_lcell_comb \Mux21~8 (
// Equation(s):
// \Mux21~8_combout  = (\Mux21~7_combout  & (((\registerArray[31][10]~q ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux21~7_combout  & (\registerArray[27][10]~q  & ((\my_rf.rsel1[3]~input_o ))))

	.dataa(\registerArray[27][10]~q ),
	.datab(\Mux21~7_combout ),
	.datac(\registerArray[31][10]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux21~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~8 .lut_mask = 16'hE2CC;
defparam \Mux21~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N7
dffeas \registerArray[28][10] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[10]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][10] .is_wysiwyg = "true";
defparam \registerArray[28][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N14
cycloneive_lcell_comb \Mux21~4 (
// Equation(s):
// \Mux21~4_combout  = (\my_rf.rsel1[2]~input_o  & (\my_rf.rsel1[3]~input_o )) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & ((\registerArray[24][10]~q ))) # (!\my_rf.rsel1[3]~input_o  & (\registerArray[16][10]~q ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[16][10]~q ),
	.datad(\registerArray[24][10]~q ),
	.cin(gnd),
	.combout(\Mux21~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~4 .lut_mask = 16'hDC98;
defparam \Mux21~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N6
cycloneive_lcell_comb \Mux21~5 (
// Equation(s):
// \Mux21~5_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux21~4_combout  & ((\registerArray[28][10]~q ))) # (!\Mux21~4_combout  & (\registerArray[20][10]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux21~4_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[20][10]~q ),
	.datac(\registerArray[28][10]~q ),
	.datad(\Mux21~4_combout ),
	.cin(gnd),
	.combout(\Mux21~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~5 .lut_mask = 16'hF588;
defparam \Mux21~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N20
cycloneive_lcell_comb \Mux21~6 (
// Equation(s):
// \Mux21~6_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux21~3_combout ) # ((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & (((!\my_rf.rsel1[0]~input_o  & \Mux21~5_combout ))))

	.dataa(\Mux21~3_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\Mux21~5_combout ),
	.cin(gnd),
	.combout(\Mux21~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~6 .lut_mask = 16'hCBC8;
defparam \Mux21~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N6
cycloneive_lcell_comb \Mux21~9 (
// Equation(s):
// \Mux21~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux21~6_combout  & ((\Mux21~8_combout ))) # (!\Mux21~6_combout  & (\Mux21~1_combout )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux21~6_combout ))))

	.dataa(\Mux21~1_combout ),
	.datab(\Mux21~8_combout ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\Mux21~6_combout ),
	.cin(gnd),
	.combout(\Mux21~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~9 .lut_mask = 16'hCFA0;
defparam \Mux21~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N30
cycloneive_lcell_comb \Mux21~20 (
// Equation(s):
// \Mux21~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux21~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux21~19_combout ))

	.dataa(gnd),
	.datab(\Mux21~19_combout ),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux21~9_combout ),
	.cin(gnd),
	.combout(\Mux21~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~20 .lut_mask = 16'hFC0C;
defparam \Mux21~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N27
dffeas \registerArray[15][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][11] .is_wysiwyg = "true";
defparam \registerArray[15][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N17
dffeas \registerArray[14][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][11] .is_wysiwyg = "true";
defparam \registerArray[14][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N26
cycloneive_lcell_comb \Mux20~18 (
// Equation(s):
// \Mux20~18_combout  = (\Mux20~17_combout  & (((\registerArray[15][11]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux20~17_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[14][11]~q ))))

	.dataa(\Mux20~17_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][11]~q ),
	.datad(\registerArray[14][11]~q ),
	.cin(gnd),
	.combout(\Mux20~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~18 .lut_mask = 16'hE6A2;
defparam \Mux20~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N6
cycloneive_lcell_comb \Mux20~11 (
// Equation(s):
// \Mux20~11_combout  = (\Mux20~10_combout  & (((\registerArray[7][11]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux20~10_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[6][11]~q ))))

	.dataa(\Mux20~10_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[7][11]~q ),
	.datad(\registerArray[6][11]~q ),
	.cin(gnd),
	.combout(\Mux20~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~11 .lut_mask = 16'hE6A2;
defparam \Mux20~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N4
cycloneive_lcell_comb \Mux20~19 (
// Equation(s):
// \Mux20~19_combout  = (\Mux20~16_combout  & ((\Mux20~18_combout ) # ((!\my_rf.rsel1[2]~input_o )))) # (!\Mux20~16_combout  & (((\my_rf.rsel1[2]~input_o  & \Mux20~11_combout ))))

	.dataa(\Mux20~16_combout ),
	.datab(\Mux20~18_combout ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux20~11_combout ),
	.cin(gnd),
	.combout(\Mux20~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~19 .lut_mask = 16'hDA8A;
defparam \Mux20~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N29
dffeas \registerArray[29][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][11] .is_wysiwyg = "true";
defparam \registerArray[29][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N5
dffeas \registerArray[17][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][11] .is_wysiwyg = "true";
defparam \registerArray[17][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N4
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// \Mux20~0_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[25][11]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[17][11]~q )))))

	.dataa(\registerArray[25][11]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[17][11]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'hEE30;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N28
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// \Mux20~1_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux20~0_combout  & ((\registerArray[29][11]~q ))) # (!\Mux20~0_combout  & (\registerArray[21][11]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux20~0_combout ))))

	.dataa(\registerArray[21][11]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[29][11]~q ),
	.datad(\Mux20~0_combout ),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'hF388;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y36_N27
dffeas \registerArray[18][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][11] .is_wysiwyg = "true";
defparam \registerArray[18][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N26
cycloneive_lcell_comb \Mux20~2 (
// Equation(s):
// \Mux20~2_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & (\registerArray[22][11]~q )) # (!\my_rf.rsel1[2]~input_o  & ((\registerArray[18][11]~q )))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[22][11]~q ),
	.datac(\registerArray[18][11]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux20~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~2 .lut_mask = 16'hEE50;
defparam \Mux20~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y36_N23
dffeas \registerArray[30][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][11] .is_wysiwyg = "true";
defparam \registerArray[30][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y36_N22
cycloneive_lcell_comb \Mux20~3 (
// Equation(s):
// \Mux20~3_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux20~2_combout  & (\registerArray[30][11]~q )) # (!\Mux20~2_combout  & ((\registerArray[26][11]~q ))))) # (!\my_rf.rsel1[3]~input_o  & (\Mux20~2_combout ))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux20~2_combout ),
	.datac(\registerArray[30][11]~q ),
	.datad(\registerArray[26][11]~q ),
	.cin(gnd),
	.combout(\Mux20~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~3 .lut_mask = 16'hE6C4;
defparam \Mux20~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N27
dffeas \registerArray[28][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][11] .is_wysiwyg = "true";
defparam \registerArray[28][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y37_N11
dffeas \registerArray[16][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][11] .is_wysiwyg = "true";
defparam \registerArray[16][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y37_N1
dffeas \registerArray[20][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][11] .is_wysiwyg = "true";
defparam \registerArray[20][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N10
cycloneive_lcell_comb \Mux20~4 (
// Equation(s):
// \Mux20~4_combout  = (\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o ) # ((\registerArray[20][11]~q )))) # (!\my_rf.rsel1[2]~input_o  & (!\my_rf.rsel1[3]~input_o  & (\registerArray[16][11]~q )))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[16][11]~q ),
	.datad(\registerArray[20][11]~q ),
	.cin(gnd),
	.combout(\Mux20~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~4 .lut_mask = 16'hBA98;
defparam \Mux20~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N26
cycloneive_lcell_comb \Mux20~5 (
// Equation(s):
// \Mux20~5_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux20~4_combout  & ((\registerArray[28][11]~q ))) # (!\Mux20~4_combout  & (\registerArray[24][11]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux20~4_combout ))))

	.dataa(\registerArray[24][11]~q ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[28][11]~q ),
	.datad(\Mux20~4_combout ),
	.cin(gnd),
	.combout(\Mux20~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~5 .lut_mask = 16'hF388;
defparam \Mux20~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N8
cycloneive_lcell_comb \Mux20~6 (
// Equation(s):
// \Mux20~6_combout  = (\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o )) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\Mux20~3_combout )) # (!\my_rf.rsel1[1]~input_o  & ((\Mux20~5_combout )))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\Mux20~3_combout ),
	.datad(\Mux20~5_combout ),
	.cin(gnd),
	.combout(\Mux20~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~6 .lut_mask = 16'hD9C8;
defparam \Mux20~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y33_N27
dffeas \registerArray[31][11] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[11]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][11] .is_wysiwyg = "true";
defparam \registerArray[31][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N26
cycloneive_lcell_comb \Mux20~8 (
// Equation(s):
// \Mux20~8_combout  = (\Mux20~7_combout  & (((\registerArray[31][11]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux20~7_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[23][11]~q ))))

	.dataa(\Mux20~7_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[31][11]~q ),
	.datad(\registerArray[23][11]~q ),
	.cin(gnd),
	.combout(\Mux20~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~8 .lut_mask = 16'hE6A2;
defparam \Mux20~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N2
cycloneive_lcell_comb \Mux20~9 (
// Equation(s):
// \Mux20~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux20~6_combout  & ((\Mux20~8_combout ))) # (!\Mux20~6_combout  & (\Mux20~1_combout )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux20~6_combout ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux20~1_combout ),
	.datac(\Mux20~6_combout ),
	.datad(\Mux20~8_combout ),
	.cin(gnd),
	.combout(\Mux20~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~9 .lut_mask = 16'hF858;
defparam \Mux20~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N14
cycloneive_lcell_comb \Mux20~20 (
// Equation(s):
// \Mux20~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux20~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux20~19_combout ))

	.dataa(gnd),
	.datab(\Mux20~19_combout ),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux20~9_combout ),
	.cin(gnd),
	.combout(\Mux20~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~20 .lut_mask = 16'hFC0C;
defparam \Mux20~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y32_N17
dffeas \registerArray[17][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][12] .is_wysiwyg = "true";
defparam \registerArray[17][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N16
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (\my_rf.rsel1[2]~input_o  & ((\registerArray[21][12]~q ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\registerArray[17][12]~q  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\registerArray[21][12]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[17][12]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'hCCB8;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N26
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// \Mux19~1_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux19~0_combout  & ((\registerArray[29][12]~q ))) # (!\Mux19~0_combout  & (\registerArray[25][12]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux19~0_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[25][12]~q ),
	.datac(\registerArray[29][12]~q ),
	.datad(\Mux19~0_combout ),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'hF588;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y33_N1
dffeas \registerArray[27][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][12] .is_wysiwyg = "true";
defparam \registerArray[27][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y32_N29
dffeas \registerArray[31][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][12] .is_wysiwyg = "true";
defparam \registerArray[31][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y33_N27
dffeas \registerArray[19][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][12] .is_wysiwyg = "true";
defparam \registerArray[19][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N26
cycloneive_lcell_comb \Mux19~7 (
// Equation(s):
// \Mux19~7_combout  = (\my_rf.rsel1[2]~input_o  & ((\registerArray[23][12]~q ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\registerArray[19][12]~q  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\registerArray[23][12]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[19][12]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux19~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~7 .lut_mask = 16'hCCB8;
defparam \Mux19~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N28
cycloneive_lcell_comb \Mux19~8 (
// Equation(s):
// \Mux19~8_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux19~7_combout  & ((\registerArray[31][12]~q ))) # (!\Mux19~7_combout  & (\registerArray[27][12]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux19~7_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[27][12]~q ),
	.datac(\registerArray[31][12]~q ),
	.datad(\Mux19~7_combout ),
	.cin(gnd),
	.combout(\Mux19~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~8 .lut_mask = 16'hF588;
defparam \Mux19~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N0
cycloneive_lcell_comb \Mux19~9 (
// Equation(s):
// \Mux19~9_combout  = (\Mux19~6_combout  & (((\Mux19~8_combout )) # (!\my_rf.rsel1[0]~input_o ))) # (!\Mux19~6_combout  & (\my_rf.rsel1[0]~input_o  & (\Mux19~1_combout )))

	.dataa(\Mux19~6_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux19~1_combout ),
	.datad(\Mux19~8_combout ),
	.cin(gnd),
	.combout(\Mux19~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~9 .lut_mask = 16'hEA62;
defparam \Mux19~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N13
dffeas \registerArray[2][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][12] .is_wysiwyg = "true";
defparam \registerArray[2][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N23
dffeas \registerArray[1][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][12] .is_wysiwyg = "true";
defparam \registerArray[1][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N21
dffeas \registerArray[3][12] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[12]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][12] .is_wysiwyg = "true";
defparam \registerArray[3][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N22
cycloneive_lcell_comb \Mux19~14 (
// Equation(s):
// \Mux19~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][12]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][12]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[1][12]~q ),
	.datad(\registerArray[3][12]~q ),
	.cin(gnd),
	.combout(\Mux19~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~14 .lut_mask = 16'hC840;
defparam \Mux19~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N2
cycloneive_lcell_comb \Mux19~15 (
// Equation(s):
// \Mux19~15_combout  = (\Mux19~14_combout ) # ((\my_rf.rsel1[1]~input_o  & (\registerArray[2][12]~q  & !\my_rf.rsel1[0]~input_o )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[2][12]~q ),
	.datac(\Mux19~14_combout ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux19~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~15 .lut_mask = 16'hF0F8;
defparam \Mux19~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N20
cycloneive_lcell_comb \Mux19~16 (
// Equation(s):
// \Mux19~16_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux19~13_combout ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((!\my_rf.rsel1[3]~input_o  & \Mux19~15_combout ))))

	.dataa(\Mux19~13_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\my_rf.rsel1[3]~input_o ),
	.datad(\Mux19~15_combout ),
	.cin(gnd),
	.combout(\Mux19~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~16 .lut_mask = 16'hCBC8;
defparam \Mux19~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N30
cycloneive_lcell_comb \Mux19~17 (
// Equation(s):
// \Mux19~17_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[13][12]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[12][12]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[12][12]~q ),
	.datad(\registerArray[13][12]~q ),
	.cin(gnd),
	.combout(\Mux19~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~17 .lut_mask = 16'hDC98;
defparam \Mux19~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N0
cycloneive_lcell_comb \Mux19~18 (
// Equation(s):
// \Mux19~18_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux19~17_combout  & ((\registerArray[15][12]~q ))) # (!\Mux19~17_combout  & (\registerArray[14][12]~q )))) # (!\my_rf.rsel1[1]~input_o  & (((\Mux19~17_combout ))))

	.dataa(\registerArray[14][12]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][12]~q ),
	.datad(\Mux19~17_combout ),
	.cin(gnd),
	.combout(\Mux19~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~18 .lut_mask = 16'hF388;
defparam \Mux19~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N6
cycloneive_lcell_comb \Mux19~19 (
// Equation(s):
// \Mux19~19_combout  = (\Mux19~16_combout  & (((\Mux19~18_combout ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux19~16_combout  & (\Mux19~11_combout  & ((\my_rf.rsel1[3]~input_o ))))

	.dataa(\Mux19~11_combout ),
	.datab(\Mux19~16_combout ),
	.datac(\Mux19~18_combout ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux19~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~19 .lut_mask = 16'hE2CC;
defparam \Mux19~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N8
cycloneive_lcell_comb \Mux19~20 (
// Equation(s):
// \Mux19~20_combout  = (\my_rf.rsel1[4]~input_o  & (\Mux19~9_combout )) # (!\my_rf.rsel1[4]~input_o  & ((\Mux19~19_combout )))

	.dataa(gnd),
	.datab(\Mux19~9_combout ),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux19~19_combout ),
	.cin(gnd),
	.combout(\Mux19~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~20 .lut_mask = 16'hCFC0;
defparam \Mux19~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N31
dffeas \registerArray[7][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][13] .is_wysiwyg = "true";
defparam \registerArray[7][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N30
cycloneive_lcell_comb \Mux18~11 (
// Equation(s):
// \Mux18~11_combout  = (\Mux18~10_combout  & (((\registerArray[7][13]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux18~10_combout  & (\registerArray[6][13]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux18~10_combout ),
	.datab(\registerArray[6][13]~q ),
	.datac(\registerArray[7][13]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux18~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~11 .lut_mask = 16'hE4AA;
defparam \Mux18~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y36_N26
cycloneive_lcell_comb \Mux18~17 (
// Equation(s):
// \Mux18~17_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[13][13]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[12][13]~q )))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[13][13]~q ),
	.datac(\registerArray[12][13]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux18~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~17 .lut_mask = 16'hEE50;
defparam \Mux18~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N28
cycloneive_lcell_comb \Mux18~18 (
// Equation(s):
// \Mux18~18_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux18~17_combout  & ((\registerArray[15][13]~q ))) # (!\Mux18~17_combout  & (\registerArray[14][13]~q )))) # (!\my_rf.rsel1[1]~input_o  & (((\Mux18~17_combout ))))

	.dataa(\registerArray[14][13]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][13]~q ),
	.datad(\Mux18~17_combout ),
	.cin(gnd),
	.combout(\Mux18~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~18 .lut_mask = 16'hF388;
defparam \Mux18~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N22
cycloneive_lcell_comb \Mux18~19 (
// Equation(s):
// \Mux18~19_combout  = (\Mux18~16_combout  & (((\Mux18~18_combout ) # (!\my_rf.rsel1[2]~input_o )))) # (!\Mux18~16_combout  & (\Mux18~11_combout  & (\my_rf.rsel1[2]~input_o )))

	.dataa(\Mux18~16_combout ),
	.datab(\Mux18~11_combout ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux18~18_combout ),
	.cin(gnd),
	.combout(\Mux18~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~19 .lut_mask = 16'hEA4A;
defparam \Mux18~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y37_N19
dffeas \registerArray[28][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][13] .is_wysiwyg = "true";
defparam \registerArray[28][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N27
dffeas \registerArray[16][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][13] .is_wysiwyg = "true";
defparam \registerArray[16][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y37_N9
dffeas \registerArray[20][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][13] .is_wysiwyg = "true";
defparam \registerArray[20][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N26
cycloneive_lcell_comb \Mux18~4 (
// Equation(s):
// \Mux18~4_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[20][13]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[16][13]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[16][13]~q ),
	.datad(\registerArray[20][13]~q ),
	.cin(gnd),
	.combout(\Mux18~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~4 .lut_mask = 16'hDC98;
defparam \Mux18~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N18
cycloneive_lcell_comb \Mux18~5 (
// Equation(s):
// \Mux18~5_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux18~4_combout  & ((\registerArray[28][13]~q ))) # (!\Mux18~4_combout  & (\registerArray[24][13]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux18~4_combout ))))

	.dataa(\registerArray[24][13]~q ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[28][13]~q ),
	.datad(\Mux18~4_combout ),
	.cin(gnd),
	.combout(\Mux18~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~5 .lut_mask = 16'hF388;
defparam \Mux18~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y36_N11
dffeas \registerArray[18][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][13] .is_wysiwyg = "true";
defparam \registerArray[18][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y36_N25
dffeas \registerArray[22][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][13] .is_wysiwyg = "true";
defparam \registerArray[22][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N10
cycloneive_lcell_comb \Mux18~2 (
// Equation(s):
// \Mux18~2_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[22][13]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][13]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][13]~q ),
	.datad(\registerArray[22][13]~q ),
	.cin(gnd),
	.combout(\Mux18~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~2 .lut_mask = 16'hDC98;
defparam \Mux18~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N26
cycloneive_lcell_comb \Mux18~3 (
// Equation(s):
// \Mux18~3_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux18~2_combout  & ((\registerArray[30][13]~q ))) # (!\Mux18~2_combout  & (\registerArray[26][13]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux18~2_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[26][13]~q ),
	.datac(\registerArray[30][13]~q ),
	.datad(\Mux18~2_combout ),
	.cin(gnd),
	.combout(\Mux18~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~3 .lut_mask = 16'hF588;
defparam \Mux18~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N2
cycloneive_lcell_comb \Mux18~6 (
// Equation(s):
// \Mux18~6_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\Mux18~3_combout ))) # (!\my_rf.rsel1[1]~input_o  & (\Mux18~5_combout ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux18~5_combout ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\Mux18~3_combout ),
	.cin(gnd),
	.combout(\Mux18~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~6 .lut_mask = 16'hF4A4;
defparam \Mux18~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y34_N11
dffeas \registerArray[29][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][13] .is_wysiwyg = "true";
defparam \registerArray[29][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y0_N10
dffeas \registerArray[21][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[13]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][13] .is_wysiwyg = "true";
defparam \registerArray[21][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N10
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// \Mux18~1_combout  = (\Mux18~0_combout  & (((\registerArray[29][13]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux18~0_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[21][13]~q ))))

	.dataa(\Mux18~0_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[29][13]~q ),
	.datad(\registerArray[21][13]~q ),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'hE6A2;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y33_N31
dffeas \registerArray[31][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][13] .is_wysiwyg = "true";
defparam \registerArray[31][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y33_N29
dffeas \registerArray[19][13] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[13]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][13] .is_wysiwyg = "true";
defparam \registerArray[19][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N28
cycloneive_lcell_comb \Mux18~7 (
// Equation(s):
// \Mux18~7_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[27][13]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[19][13]~q )))))

	.dataa(\registerArray[27][13]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[19][13]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux18~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~7 .lut_mask = 16'hEE30;
defparam \Mux18~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N30
cycloneive_lcell_comb \Mux18~8 (
// Equation(s):
// \Mux18~8_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux18~7_combout  & ((\registerArray[31][13]~q ))) # (!\Mux18~7_combout  & (\registerArray[23][13]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux18~7_combout ))))

	.dataa(\registerArray[23][13]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[31][13]~q ),
	.datad(\Mux18~7_combout ),
	.cin(gnd),
	.combout(\Mux18~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~8 .lut_mask = 16'hF388;
defparam \Mux18~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N12
cycloneive_lcell_comb \Mux18~9 (
// Equation(s):
// \Mux18~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux18~6_combout  & ((\Mux18~8_combout ))) # (!\Mux18~6_combout  & (\Mux18~1_combout )))) # (!\my_rf.rsel1[0]~input_o  & (\Mux18~6_combout ))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux18~6_combout ),
	.datac(\Mux18~1_combout ),
	.datad(\Mux18~8_combout ),
	.cin(gnd),
	.combout(\Mux18~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~9 .lut_mask = 16'hEC64;
defparam \Mux18~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N8
cycloneive_lcell_comb \Mux18~20 (
// Equation(s):
// \Mux18~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux18~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux18~19_combout ))

	.dataa(gnd),
	.datab(\my_rf.rsel1[4]~input_o ),
	.datac(\Mux18~19_combout ),
	.datad(\Mux18~9_combout ),
	.cin(gnd),
	.combout(\Mux18~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~20 .lut_mask = 16'hFC30;
defparam \Mux18~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N23
dffeas \registerArray[15][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][14] .is_wysiwyg = "true";
defparam \registerArray[15][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N22
cycloneive_lcell_comb \Mux17~18 (
// Equation(s):
// \Mux17~18_combout  = (\Mux17~17_combout  & (((\registerArray[15][14]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux17~17_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[14][14]~q ))))

	.dataa(\Mux17~17_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][14]~q ),
	.datad(\registerArray[14][14]~q ),
	.cin(gnd),
	.combout(\Mux17~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~18 .lut_mask = 16'hE6A2;
defparam \Mux17~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y37_N19
dffeas \registerArray[8][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][14] .is_wysiwyg = "true";
defparam \registerArray[8][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y37_N17
dffeas \registerArray[10][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][14] .is_wysiwyg = "true";
defparam \registerArray[10][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y37_N18
cycloneive_lcell_comb \Mux17~10 (
// Equation(s):
// \Mux17~10_combout  = (\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o )) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[10][14]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[8][14]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[8][14]~q ),
	.datad(\registerArray[10][14]~q ),
	.cin(gnd),
	.combout(\Mux17~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~10 .lut_mask = 16'hDC98;
defparam \Mux17~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y37_N18
cycloneive_lcell_comb \Mux17~11 (
// Equation(s):
// \Mux17~11_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux17~10_combout  & (\registerArray[11][14]~q )) # (!\Mux17~10_combout  & ((\registerArray[9][14]~q ))))) # (!\my_rf.rsel1[0]~input_o  & (\Mux17~10_combout ))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux17~10_combout ),
	.datac(\registerArray[11][14]~q ),
	.datad(\registerArray[9][14]~q ),
	.cin(gnd),
	.combout(\Mux17~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~11 .lut_mask = 16'hE6C4;
defparam \Mux17~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N23
dffeas \registerArray[2][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][14] .is_wysiwyg = "true";
defparam \registerArray[2][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N5
dffeas \registerArray[3][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][14] .is_wysiwyg = "true";
defparam \registerArray[3][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y36_N15
dffeas \registerArray[1][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][14] .is_wysiwyg = "true";
defparam \registerArray[1][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y36_N14
cycloneive_lcell_comb \Mux17~14 (
// Equation(s):
// \Mux17~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\registerArray[3][14]~q )) # (!\my_rf.rsel1[1]~input_o  & ((\registerArray[1][14]~q )))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[3][14]~q ),
	.datac(\registerArray[1][14]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux17~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~14 .lut_mask = 16'hD800;
defparam \Mux17~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y38_N14
cycloneive_lcell_comb \Mux17~15 (
// Equation(s):
// \Mux17~15_combout  = (\Mux17~14_combout ) # ((\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & \registerArray[2][14]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[2][14]~q ),
	.datad(\Mux17~14_combout ),
	.cin(gnd),
	.combout(\Mux17~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~15 .lut_mask = 16'hFF20;
defparam \Mux17~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N1
dffeas \registerArray[6][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][14] .is_wysiwyg = "true";
defparam \registerArray[6][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N19
dffeas \registerArray[7][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][14] .is_wysiwyg = "true";
defparam \registerArray[7][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N18
cycloneive_lcell_comb \Mux17~13 (
// Equation(s):
// \Mux17~13_combout  = (\Mux17~12_combout  & (((\registerArray[7][14]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux17~12_combout  & (\registerArray[6][14]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux17~12_combout ),
	.datab(\registerArray[6][14]~q ),
	.datac(\registerArray[7][14]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux17~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~13 .lut_mask = 16'hE4AA;
defparam \Mux17~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y38_N0
cycloneive_lcell_comb \Mux17~16 (
// Equation(s):
// \Mux17~16_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\Mux17~13_combout ))) # (!\my_rf.rsel1[2]~input_o  & (\Mux17~15_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux17~15_combout ),
	.datad(\Mux17~13_combout ),
	.cin(gnd),
	.combout(\Mux17~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~16 .lut_mask = 16'hDC98;
defparam \Mux17~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y38_N2
cycloneive_lcell_comb \Mux17~19 (
// Equation(s):
// \Mux17~19_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux17~16_combout  & (\Mux17~18_combout )) # (!\Mux17~16_combout  & ((\Mux17~11_combout ))))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux17~16_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux17~18_combout ),
	.datac(\Mux17~11_combout ),
	.datad(\Mux17~16_combout ),
	.cin(gnd),
	.combout(\Mux17~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~19 .lut_mask = 16'hDDA0;
defparam \Mux17~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N8
cycloneive_lcell_comb \Mux17~8 (
// Equation(s):
// \Mux17~8_combout  = (\Mux17~7_combout  & (((\registerArray[31][14]~q )) # (!\my_rf.rsel1[3]~input_o ))) # (!\Mux17~7_combout  & (\my_rf.rsel1[3]~input_o  & ((\registerArray[27][14]~q ))))

	.dataa(\Mux17~7_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[31][14]~q ),
	.datad(\registerArray[27][14]~q ),
	.cin(gnd),
	.combout(\Mux17~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~8 .lut_mask = 16'hE6A2;
defparam \Mux17~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y32_N23
dffeas \registerArray[17][14] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[14]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][14] .is_wysiwyg = "true";
defparam \registerArray[17][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N22
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// \Mux17~0_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[21][14]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[17][14]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[17][14]~q ),
	.datad(\registerArray[21][14]~q ),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'hDC98;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N16
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// \Mux17~1_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux17~0_combout  & (\registerArray[29][14]~q )) # (!\Mux17~0_combout  & ((\registerArray[25][14]~q ))))) # (!\my_rf.rsel1[3]~input_o  & (\Mux17~0_combout ))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux17~0_combout ),
	.datac(\registerArray[29][14]~q ),
	.datad(\registerArray[25][14]~q ),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hE6C4;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y38_N12
cycloneive_lcell_comb \Mux17~9 (
// Equation(s):
// \Mux17~9_combout  = (\Mux17~6_combout  & (((\Mux17~8_combout )) # (!\my_rf.rsel1[0]~input_o ))) # (!\Mux17~6_combout  & (\my_rf.rsel1[0]~input_o  & ((\Mux17~1_combout ))))

	.dataa(\Mux17~6_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux17~8_combout ),
	.datad(\Mux17~1_combout ),
	.cin(gnd),
	.combout(\Mux17~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~9 .lut_mask = 16'hE6A2;
defparam \Mux17~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y38_N28
cycloneive_lcell_comb \Mux17~20 (
// Equation(s):
// \Mux17~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux17~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux17~19_combout ))

	.dataa(gnd),
	.datab(\Mux17~19_combout ),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux17~9_combout ),
	.cin(gnd),
	.combout(\Mux17~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~20 .lut_mask = 16'hFC0C;
defparam \Mux17~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y36_N19
dffeas \registerArray[18][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][15] .is_wysiwyg = "true";
defparam \registerArray[18][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y36_N1
dffeas \registerArray[22][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][15] .is_wysiwyg = "true";
defparam \registerArray[22][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y36_N18
cycloneive_lcell_comb \Mux16~2 (
// Equation(s):
// \Mux16~2_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[22][15]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][15]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][15]~q ),
	.datad(\registerArray[22][15]~q ),
	.cin(gnd),
	.combout(\Mux16~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~2 .lut_mask = 16'hDC98;
defparam \Mux16~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N28
cycloneive_lcell_comb \Mux16~3 (
// Equation(s):
// \Mux16~3_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux16~2_combout  & (\registerArray[30][15]~q )) # (!\Mux16~2_combout  & ((\registerArray[26][15]~q ))))) # (!\my_rf.rsel1[3]~input_o  & (\Mux16~2_combout ))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux16~2_combout ),
	.datac(\registerArray[30][15]~q ),
	.datad(\registerArray[26][15]~q ),
	.cin(gnd),
	.combout(\Mux16~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~3 .lut_mask = 16'hE6C4;
defparam \Mux16~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y36_N14
cycloneive_lcell_comb \Mux16~6 (
// Equation(s):
// \Mux16~6_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\Mux16~3_combout ))) # (!\my_rf.rsel1[1]~input_o  & (\Mux16~5_combout ))))

	.dataa(\Mux16~5_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\Mux16~3_combout ),
	.cin(gnd),
	.combout(\Mux16~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~6 .lut_mask = 16'hF2C2;
defparam \Mux16~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N0
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// \Mux16~0_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[25][15]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[17][15]~q )))))

	.dataa(\registerArray[25][15]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[17][15]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'hEE30;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N16
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// \Mux16~1_combout  = (\Mux16~0_combout  & (((\registerArray[29][15]~q ) # (!\my_rf.rsel1[2]~input_o )))) # (!\Mux16~0_combout  & (\registerArray[21][15]~q  & ((\my_rf.rsel1[2]~input_o ))))

	.dataa(\registerArray[21][15]~q ),
	.datab(\Mux16~0_combout ),
	.datac(\registerArray[29][15]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hE2CC;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y36_N16
cycloneive_lcell_comb \Mux16~9 (
// Equation(s):
// \Mux16~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux16~6_combout  & (\Mux16~8_combout )) # (!\Mux16~6_combout  & ((\Mux16~1_combout ))))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux16~6_combout ))))

	.dataa(\Mux16~8_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux16~6_combout ),
	.datad(\Mux16~1_combout ),
	.cin(gnd),
	.combout(\Mux16~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~9 .lut_mask = 16'hBCB0;
defparam \Mux16~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N7
dffeas \registerArray[4][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][15] .is_wysiwyg = "true";
defparam \registerArray[4][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N6
cycloneive_lcell_comb \Mux16~10 (
// Equation(s):
// \Mux16~10_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[5][15]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[4][15]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[4][15]~q ),
	.datad(\registerArray[5][15]~q ),
	.cin(gnd),
	.combout(\Mux16~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~10 .lut_mask = 16'hDC98;
defparam \Mux16~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N4
cycloneive_lcell_comb \Mux16~11 (
// Equation(s):
// \Mux16~11_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux16~10_combout  & ((\registerArray[7][15]~q ))) # (!\Mux16~10_combout  & (\registerArray[6][15]~q )))) # (!\my_rf.rsel1[1]~input_o  & (((\Mux16~10_combout ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[6][15]~q ),
	.datac(\registerArray[7][15]~q ),
	.datad(\Mux16~10_combout ),
	.cin(gnd),
	.combout(\Mux16~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~11 .lut_mask = 16'hF588;
defparam \Mux16~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N5
dffeas \registerArray[14][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][15] .is_wysiwyg = "true";
defparam \registerArray[14][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y35_N15
dffeas \registerArray[15][15] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[15]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][15] .is_wysiwyg = "true";
defparam \registerArray[15][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N14
cycloneive_lcell_comb \Mux16~18 (
// Equation(s):
// \Mux16~18_combout  = (\Mux16~17_combout  & (((\registerArray[15][15]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux16~17_combout  & (\registerArray[14][15]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux16~17_combout ),
	.datab(\registerArray[14][15]~q ),
	.datac(\registerArray[15][15]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux16~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~18 .lut_mask = 16'hE4AA;
defparam \Mux16~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y38_N24
cycloneive_lcell_comb \Mux16~19 (
// Equation(s):
// \Mux16~19_combout  = (\Mux16~16_combout  & (((\Mux16~18_combout )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux16~16_combout  & (\my_rf.rsel1[2]~input_o  & (\Mux16~11_combout )))

	.dataa(\Mux16~16_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux16~11_combout ),
	.datad(\Mux16~18_combout ),
	.cin(gnd),
	.combout(\Mux16~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~19 .lut_mask = 16'hEA62;
defparam \Mux16~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y38_N10
cycloneive_lcell_comb \Mux16~20 (
// Equation(s):
// \Mux16~20_combout  = (\my_rf.rsel1[4]~input_o  & (\Mux16~9_combout )) # (!\my_rf.rsel1[4]~input_o  & ((\Mux16~19_combout )))

	.dataa(gnd),
	.datab(\Mux16~9_combout ),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux16~19_combout ),
	.cin(gnd),
	.combout(\Mux16~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~20 .lut_mask = 16'hCFC0;
defparam \Mux16~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N21
dffeas \registerArray[29][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][16] .is_wysiwyg = "true";
defparam \registerArray[29][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N28
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// \Mux15~0_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\registerArray[21][16]~q ))) # (!\my_rf.rsel1[2]~input_o  & (\registerArray[17][16]~q ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[17][16]~q ),
	.datad(\registerArray[21][16]~q ),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hDC98;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N20
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// \Mux15~1_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux15~0_combout  & ((\registerArray[29][16]~q ))) # (!\Mux15~0_combout  & (\registerArray[25][16]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux15~0_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[25][16]~q ),
	.datac(\registerArray[29][16]~q ),
	.datad(\Mux15~0_combout ),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'hF588;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y38_N15
dffeas \registerArray[26][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][16] .is_wysiwyg = "true";
defparam \registerArray[26][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y38_N17
dffeas \registerArray[18][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][16] .is_wysiwyg = "true";
defparam \registerArray[18][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N16
cycloneive_lcell_comb \Mux15~2 (
// Equation(s):
// \Mux15~2_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[26][16]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[18][16]~q )))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[26][16]~q ),
	.datac(\registerArray[18][16]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux15~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~2 .lut_mask = 16'hEE50;
defparam \Mux15~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N30
cycloneive_lcell_comb \Mux15~3 (
// Equation(s):
// \Mux15~3_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux15~2_combout  & (\registerArray[30][16]~q )) # (!\Mux15~2_combout  & ((\registerArray[22][16]~q ))))) # (!\my_rf.rsel1[2]~input_o  & (\Mux15~2_combout ))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux15~2_combout ),
	.datac(\registerArray[30][16]~q ),
	.datad(\registerArray[22][16]~q ),
	.cin(gnd),
	.combout(\Mux15~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~3 .lut_mask = 16'hE6C4;
defparam \Mux15~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y35_N21
dffeas \registerArray[28][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][16] .is_wysiwyg = "true";
defparam \registerArray[28][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y35_N9
dffeas \registerArray[20][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][16] .is_wysiwyg = "true";
defparam \registerArray[20][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N20
cycloneive_lcell_comb \Mux15~5 (
// Equation(s):
// \Mux15~5_combout  = (\Mux15~4_combout  & (((\registerArray[28][16]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux15~4_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[20][16]~q ))))

	.dataa(\Mux15~4_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[28][16]~q ),
	.datad(\registerArray[20][16]~q ),
	.cin(gnd),
	.combout(\Mux15~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~5 .lut_mask = 16'hE6A2;
defparam \Mux15~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N18
cycloneive_lcell_comb \Mux15~6 (
// Equation(s):
// \Mux15~6_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux15~3_combout ) # ((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & (((!\my_rf.rsel1[0]~input_o  & \Mux15~5_combout ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\Mux15~3_combout ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\Mux15~5_combout ),
	.cin(gnd),
	.combout(\Mux15~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~6 .lut_mask = 16'hADA8;
defparam \Mux15~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N28
cycloneive_lcell_comb \Mux15~9 (
// Equation(s):
// \Mux15~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux15~6_combout  & (\Mux15~8_combout )) # (!\Mux15~6_combout  & ((\Mux15~1_combout ))))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux15~6_combout ))))

	.dataa(\Mux15~8_combout ),
	.datab(\Mux15~1_combout ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\Mux15~6_combout ),
	.cin(gnd),
	.combout(\Mux15~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~9 .lut_mask = 16'hAFC0;
defparam \Mux15~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N1
dffeas \registerArray[2][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][16] .is_wysiwyg = "true";
defparam \registerArray[2][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y32_N19
dffeas \registerArray[1][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][16] .is_wysiwyg = "true";
defparam \registerArray[1][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y32_N9
dffeas \registerArray[3][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][16] .is_wysiwyg = "true";
defparam \registerArray[3][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N18
cycloneive_lcell_comb \Mux15~14 (
// Equation(s):
// \Mux15~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][16]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][16]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[1][16]~q ),
	.datad(\registerArray[3][16]~q ),
	.cin(gnd),
	.combout(\Mux15~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~14 .lut_mask = 16'hC840;
defparam \Mux15~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N22
cycloneive_lcell_comb \Mux15~15 (
// Equation(s):
// \Mux15~15_combout  = (\Mux15~14_combout ) # ((!\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o  & \registerArray[2][16]~q )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[2][16]~q ),
	.datad(\Mux15~14_combout ),
	.cin(gnd),
	.combout(\Mux15~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~15 .lut_mask = 16'hFF40;
defparam \Mux15~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N16
cycloneive_lcell_comb \Mux15~16 (
// Equation(s):
// \Mux15~16_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux15~13_combout ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux15~15_combout  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\Mux15~13_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux15~15_combout ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux15~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~16 .lut_mask = 16'hCCB8;
defparam \Mux15~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y39_N7
dffeas \registerArray[8][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][16] .is_wysiwyg = "true";
defparam \registerArray[8][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y39_N29
dffeas \registerArray[10][16] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[16]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][16] .is_wysiwyg = "true";
defparam \registerArray[10][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N6
cycloneive_lcell_comb \Mux15~10 (
// Equation(s):
// \Mux15~10_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\registerArray[10][16]~q )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & (\registerArray[8][16]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[8][16]~q ),
	.datad(\registerArray[10][16]~q ),
	.cin(gnd),
	.combout(\Mux15~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~10 .lut_mask = 16'hBA98;
defparam \Mux15~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N14
cycloneive_lcell_comb \Mux15~11 (
// Equation(s):
// \Mux15~11_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux15~10_combout  & ((\registerArray[11][16]~q ))) # (!\Mux15~10_combout  & (\registerArray[9][16]~q )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux15~10_combout ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\registerArray[9][16]~q ),
	.datac(\registerArray[11][16]~q ),
	.datad(\Mux15~10_combout ),
	.cin(gnd),
	.combout(\Mux15~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~11 .lut_mask = 16'hF588;
defparam \Mux15~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N10
cycloneive_lcell_comb \Mux15~19 (
// Equation(s):
// \Mux15~19_combout  = (\Mux15~16_combout  & ((\Mux15~18_combout ) # ((!\my_rf.rsel1[3]~input_o )))) # (!\Mux15~16_combout  & (((\Mux15~11_combout  & \my_rf.rsel1[3]~input_o ))))

	.dataa(\Mux15~18_combout ),
	.datab(\Mux15~16_combout ),
	.datac(\Mux15~11_combout ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux15~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~19 .lut_mask = 16'hB8CC;
defparam \Mux15~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N12
cycloneive_lcell_comb \Mux15~20 (
// Equation(s):
// \Mux15~20_combout  = (\my_rf.rsel1[4]~input_o  & (\Mux15~9_combout )) # (!\my_rf.rsel1[4]~input_o  & ((\Mux15~19_combout )))

	.dataa(gnd),
	.datab(\Mux15~9_combout ),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux15~19_combout ),
	.cin(gnd),
	.combout(\Mux15~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~20 .lut_mask = 16'hCFC0;
defparam \Mux15~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y32_N23
dffeas \registerArray[1][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][17] .is_wysiwyg = "true";
defparam \registerArray[1][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N22
cycloneive_lcell_comb \Mux14~14 (
// Equation(s):
// \Mux14~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\registerArray[3][17]~q )) # (!\my_rf.rsel1[1]~input_o  & ((\registerArray[1][17]~q )))))

	.dataa(\registerArray[3][17]~q ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[1][17]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux14~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~14 .lut_mask = 16'h88C0;
defparam \Mux14~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N3
dffeas \registerArray[2][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][17] .is_wysiwyg = "true";
defparam \registerArray[2][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N18
cycloneive_lcell_comb \Mux14~15 (
// Equation(s):
// \Mux14~15_combout  = (\Mux14~14_combout ) # ((\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & \registerArray[2][17]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\Mux14~14_combout ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\registerArray[2][17]~q ),
	.cin(gnd),
	.combout(\Mux14~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~15 .lut_mask = 16'hCECC;
defparam \Mux14~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N14
cycloneive_lcell_comb \Mux14~16 (
// Equation(s):
// \Mux14~16_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\Mux14~13_combout )) # (!\my_rf.rsel1[3]~input_o  & ((\Mux14~15_combout )))))

	.dataa(\Mux14~13_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux14~15_combout ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux14~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~16 .lut_mask = 16'hEE30;
defparam \Mux14~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N28
cycloneive_lcell_comb \Mux14~18 (
// Equation(s):
// \Mux14~18_combout  = (\Mux14~17_combout  & (((\registerArray[15][17]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux14~17_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[14][17]~q ))))

	.dataa(\Mux14~17_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][17]~q ),
	.datad(\registerArray[14][17]~q ),
	.cin(gnd),
	.combout(\Mux14~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~18 .lut_mask = 16'hE6A2;
defparam \Mux14~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N0
cycloneive_lcell_comb \Mux14~19 (
// Equation(s):
// \Mux14~19_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux14~16_combout  & ((\Mux14~18_combout ))) # (!\Mux14~16_combout  & (\Mux14~11_combout )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux14~16_combout ))))

	.dataa(\Mux14~11_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux14~16_combout ),
	.datad(\Mux14~18_combout ),
	.cin(gnd),
	.combout(\Mux14~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~19 .lut_mask = 16'hF838;
defparam \Mux14~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y35_N5
dffeas \registerArray[20][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][17] .is_wysiwyg = "true";
defparam \registerArray[20][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y35_N7
dffeas \registerArray[16][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][17] .is_wysiwyg = "true";
defparam \registerArray[16][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N6
cycloneive_lcell_comb \Mux14~4 (
// Equation(s):
// \Mux14~4_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & (\registerArray[20][17]~q )) # (!\my_rf.rsel1[2]~input_o  & ((\registerArray[16][17]~q )))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[20][17]~q ),
	.datac(\registerArray[16][17]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux14~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~4 .lut_mask = 16'hEE50;
defparam \Mux14~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y35_N29
dffeas \registerArray[28][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][17] .is_wysiwyg = "true";
defparam \registerArray[28][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y35_N19
dffeas \registerArray[24][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][17] .is_wysiwyg = "true";
defparam \registerArray[24][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N28
cycloneive_lcell_comb \Mux14~5 (
// Equation(s):
// \Mux14~5_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux14~4_combout  & (\registerArray[28][17]~q )) # (!\Mux14~4_combout  & ((\registerArray[24][17]~q ))))) # (!\my_rf.rsel1[3]~input_o  & (\Mux14~4_combout ))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux14~4_combout ),
	.datac(\registerArray[28][17]~q ),
	.datad(\registerArray[24][17]~q ),
	.cin(gnd),
	.combout(\Mux14~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~5 .lut_mask = 16'hE6C4;
defparam \Mux14~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y37_N5
dffeas \registerArray[30][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][17] .is_wysiwyg = "true";
defparam \registerArray[30][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N2
cycloneive_lcell_comb \Mux14~2 (
// Equation(s):
// \Mux14~2_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & (\registerArray[22][17]~q )) # (!\my_rf.rsel1[2]~input_o  & ((\registerArray[18][17]~q )))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[22][17]~q ),
	.datac(\registerArray[18][17]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux14~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~2 .lut_mask = 16'hEE50;
defparam \Mux14~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y37_N4
cycloneive_lcell_comb \Mux14~3 (
// Equation(s):
// \Mux14~3_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux14~2_combout  & ((\registerArray[30][17]~q ))) # (!\Mux14~2_combout  & (\registerArray[26][17]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux14~2_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[26][17]~q ),
	.datac(\registerArray[30][17]~q ),
	.datad(\Mux14~2_combout ),
	.cin(gnd),
	.combout(\Mux14~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~3 .lut_mask = 16'hF588;
defparam \Mux14~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y36_N4
cycloneive_lcell_comb \Mux14~6 (
// Equation(s):
// \Mux14~6_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\Mux14~3_combout )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & (\Mux14~5_combout )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux14~5_combout ),
	.datad(\Mux14~3_combout ),
	.cin(gnd),
	.combout(\Mux14~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~6 .lut_mask = 16'hBA98;
defparam \Mux14~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y33_N11
dffeas \registerArray[31][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][17] .is_wysiwyg = "true";
defparam \registerArray[31][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y33_N25
dffeas \registerArray[23][17] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[17]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][17] .is_wysiwyg = "true";
defparam \registerArray[23][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N10
cycloneive_lcell_comb \Mux14~8 (
// Equation(s):
// \Mux14~8_combout  = (\Mux14~7_combout  & (((\registerArray[31][17]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux14~7_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[23][17]~q ))))

	.dataa(\Mux14~7_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[31][17]~q ),
	.datad(\registerArray[23][17]~q ),
	.cin(gnd),
	.combout(\Mux14~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~8 .lut_mask = 16'hE6A2;
defparam \Mux14~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y36_N22
cycloneive_lcell_comb \Mux14~9 (
// Equation(s):
// \Mux14~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux14~6_combout  & ((\Mux14~8_combout ))) # (!\Mux14~6_combout  & (\Mux14~1_combout )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux14~6_combout ))))

	.dataa(\Mux14~1_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux14~6_combout ),
	.datad(\Mux14~8_combout ),
	.cin(gnd),
	.combout(\Mux14~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~9 .lut_mask = 16'hF838;
defparam \Mux14~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N2
cycloneive_lcell_comb \Mux14~20 (
// Equation(s):
// \Mux14~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux14~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux14~19_combout ))

	.dataa(\my_rf.rsel1[4]~input_o ),
	.datab(\Mux14~19_combout ),
	.datac(gnd),
	.datad(\Mux14~9_combout ),
	.cin(gnd),
	.combout(\Mux14~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~20 .lut_mask = 16'hEE44;
defparam \Mux14~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N18
cycloneive_lcell_comb \Mux13~11 (
// Equation(s):
// \Mux13~11_combout  = (\Mux13~10_combout  & (((\registerArray[11][18]~q ) # (!\my_rf.rsel1[0]~input_o )))) # (!\Mux13~10_combout  & (\registerArray[9][18]~q  & ((\my_rf.rsel1[0]~input_o ))))

	.dataa(\Mux13~10_combout ),
	.datab(\registerArray[9][18]~q ),
	.datac(\registerArray[11][18]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux13~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~11 .lut_mask = 16'hE4AA;
defparam \Mux13~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N6
cycloneive_lcell_comb \Mux13~18 (
// Equation(s):
// \Mux13~18_combout  = (\Mux13~17_combout  & (((\registerArray[15][18]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux13~17_combout  & (\registerArray[14][18]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux13~17_combout ),
	.datab(\registerArray[14][18]~q ),
	.datac(\registerArray[15][18]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux13~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~18 .lut_mask = 16'hE4AA;
defparam \Mux13~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N12
cycloneive_lcell_comb \Mux13~19 (
// Equation(s):
// \Mux13~19_combout  = (\Mux13~16_combout  & (((\Mux13~18_combout )) # (!\my_rf.rsel1[3]~input_o ))) # (!\Mux13~16_combout  & (\my_rf.rsel1[3]~input_o  & (\Mux13~11_combout )))

	.dataa(\Mux13~16_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\Mux13~11_combout ),
	.datad(\Mux13~18_combout ),
	.cin(gnd),
	.combout(\Mux13~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~19 .lut_mask = 16'hEA62;
defparam \Mux13~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N8
cycloneive_lcell_comb \Mux13~7 (
// Equation(s):
// \Mux13~7_combout  = (\my_rf.rsel1[2]~input_o  & ((\registerArray[23][18]~q ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\registerArray[19][18]~q  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[23][18]~q ),
	.datac(\registerArray[19][18]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux13~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~7 .lut_mask = 16'hAAD8;
defparam \Mux13~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y32_N23
dffeas \registerArray[31][18] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[18]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][18] .is_wysiwyg = "true";
defparam \registerArray[31][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N22
cycloneive_lcell_comb \Mux13~8 (
// Equation(s):
// \Mux13~8_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux13~7_combout  & (\registerArray[31][18]~q )) # (!\Mux13~7_combout  & ((\registerArray[27][18]~q ))))) # (!\my_rf.rsel1[3]~input_o  & (\Mux13~7_combout ))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux13~7_combout ),
	.datac(\registerArray[31][18]~q ),
	.datad(\registerArray[27][18]~q ),
	.cin(gnd),
	.combout(\Mux13~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~8 .lut_mask = 16'hE6C4;
defparam \Mux13~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N28
cycloneive_lcell_comb \Mux13~2 (
// Equation(s):
// \Mux13~2_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[26][18]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[18][18]~q )))))

	.dataa(\registerArray[26][18]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][18]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux13~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~2 .lut_mask = 16'hEE30;
defparam \Mux13~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y37_N30
cycloneive_lcell_comb \Mux13~3 (
// Equation(s):
// \Mux13~3_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux13~2_combout  & ((\registerArray[30][18]~q ))) # (!\Mux13~2_combout  & (\registerArray[22][18]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux13~2_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[22][18]~q ),
	.datac(\registerArray[30][18]~q ),
	.datad(\Mux13~2_combout ),
	.cin(gnd),
	.combout(\Mux13~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~3 .lut_mask = 16'hF588;
defparam \Mux13~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N20
cycloneive_lcell_comb \Mux13~5 (
// Equation(s):
// \Mux13~5_combout  = (\Mux13~4_combout  & (((\registerArray[28][18]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux13~4_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[20][18]~q ))))

	.dataa(\Mux13~4_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[28][18]~q ),
	.datad(\registerArray[20][18]~q ),
	.cin(gnd),
	.combout(\Mux13~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~5 .lut_mask = 16'hE6A2;
defparam \Mux13~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N28
cycloneive_lcell_comb \Mux13~6 (
// Equation(s):
// \Mux13~6_combout  = (\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o )) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\Mux13~3_combout )) # (!\my_rf.rsel1[1]~input_o  & ((\Mux13~5_combout )))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\Mux13~3_combout ),
	.datad(\Mux13~5_combout ),
	.cin(gnd),
	.combout(\Mux13~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~6 .lut_mask = 16'hD9C8;
defparam \Mux13~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N6
cycloneive_lcell_comb \Mux13~9 (
// Equation(s):
// \Mux13~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux13~6_combout  & ((\Mux13~8_combout ))) # (!\Mux13~6_combout  & (\Mux13~1_combout )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux13~6_combout ))))

	.dataa(\Mux13~1_combout ),
	.datab(\Mux13~8_combout ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\Mux13~6_combout ),
	.cin(gnd),
	.combout(\Mux13~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~9 .lut_mask = 16'hCFA0;
defparam \Mux13~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N30
cycloneive_lcell_comb \Mux13~20 (
// Equation(s):
// \Mux13~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux13~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux13~19_combout ))

	.dataa(\my_rf.rsel1[4]~input_o ),
	.datab(\Mux13~19_combout ),
	.datac(gnd),
	.datad(\Mux13~9_combout ),
	.cin(gnd),
	.combout(\Mux13~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~20 .lut_mask = 16'hEE44;
defparam \Mux13~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N27
dffeas \registerArray[4][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][19] .is_wysiwyg = "true";
defparam \registerArray[4][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N26
cycloneive_lcell_comb \Mux12~10 (
// Equation(s):
// \Mux12~10_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[5][19]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[4][19]~q )))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[5][19]~q ),
	.datac(\registerArray[4][19]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux12~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~10 .lut_mask = 16'hEE50;
defparam \Mux12~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N14
cycloneive_lcell_comb \Mux12~11 (
// Equation(s):
// \Mux12~11_combout  = (\Mux12~10_combout  & (((\registerArray[7][19]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux12~10_combout  & (\registerArray[6][19]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\registerArray[6][19]~q ),
	.datab(\Mux12~10_combout ),
	.datac(\registerArray[7][19]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux12~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~11 .lut_mask = 16'hE2CC;
defparam \Mux12~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N14
cycloneive_lcell_comb \Mux12~15 (
// Equation(s):
// \Mux12~15_combout  = (\Mux12~14_combout ) # ((!\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o  & \registerArray[2][19]~q )))

	.dataa(\Mux12~14_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\registerArray[2][19]~q ),
	.cin(gnd),
	.combout(\Mux12~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~15 .lut_mask = 16'hBAAA;
defparam \Mux12~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N16
cycloneive_lcell_comb \Mux12~16 (
// Equation(s):
// \Mux12~16_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\Mux12~13_combout )) # (!\my_rf.rsel1[3]~input_o  & ((\Mux12~15_combout )))))

	.dataa(\Mux12~13_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux12~15_combout ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux12~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~16 .lut_mask = 16'hEE30;
defparam \Mux12~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N10
cycloneive_lcell_comb \Mux12~19 (
// Equation(s):
// \Mux12~19_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux12~16_combout  & (\Mux12~18_combout )) # (!\Mux12~16_combout  & ((\Mux12~11_combout ))))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux12~16_combout ))))

	.dataa(\Mux12~18_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux12~11_combout ),
	.datad(\Mux12~16_combout ),
	.cin(gnd),
	.combout(\Mux12~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~19 .lut_mask = 16'hBBC0;
defparam \Mux12~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y32_N31
dffeas \registerArray[29][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][19] .is_wysiwyg = "true";
defparam \registerArray[29][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N30
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// \Mux12~1_combout  = (\Mux12~0_combout  & (((\registerArray[29][19]~q ) # (!\my_rf.rsel1[2]~input_o )))) # (!\Mux12~0_combout  & (\registerArray[21][19]~q  & ((\my_rf.rsel1[2]~input_o ))))

	.dataa(\Mux12~0_combout ),
	.datab(\registerArray[21][19]~q ),
	.datac(\registerArray[29][19]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hE4AA;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y35_N25
dffeas \registerArray[28][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][19] .is_wysiwyg = "true";
defparam \registerArray[28][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N5
dffeas \registerArray[20][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][19] .is_wysiwyg = "true";
defparam \registerArray[20][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N7
dffeas \registerArray[16][19] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[19]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][19] .is_wysiwyg = "true";
defparam \registerArray[16][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N6
cycloneive_lcell_comb \Mux12~4 (
// Equation(s):
// \Mux12~4_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & (\registerArray[20][19]~q )) # (!\my_rf.rsel1[2]~input_o  & ((\registerArray[16][19]~q )))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[20][19]~q ),
	.datac(\registerArray[16][19]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux12~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~4 .lut_mask = 16'hEE50;
defparam \Mux12~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N24
cycloneive_lcell_comb \Mux12~5 (
// Equation(s):
// \Mux12~5_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux12~4_combout  & ((\registerArray[28][19]~q ))) # (!\Mux12~4_combout  & (\registerArray[24][19]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux12~4_combout ))))

	.dataa(\registerArray[24][19]~q ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[28][19]~q ),
	.datad(\Mux12~4_combout ),
	.cin(gnd),
	.combout(\Mux12~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~5 .lut_mask = 16'hF388;
defparam \Mux12~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N18
cycloneive_lcell_comb \Mux12~6 (
// Equation(s):
// \Mux12~6_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\Mux12~3_combout )) # (!\my_rf.rsel1[1]~input_o  & ((\Mux12~5_combout )))))

	.dataa(\Mux12~3_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\Mux12~5_combout ),
	.cin(gnd),
	.combout(\Mux12~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~6 .lut_mask = 16'hE3E0;
defparam \Mux12~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N12
cycloneive_lcell_comb \Mux12~9 (
// Equation(s):
// \Mux12~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux12~6_combout  & (\Mux12~8_combout )) # (!\Mux12~6_combout  & ((\Mux12~1_combout ))))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux12~6_combout ))))

	.dataa(\Mux12~8_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux12~1_combout ),
	.datad(\Mux12~6_combout ),
	.cin(gnd),
	.combout(\Mux12~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~9 .lut_mask = 16'hBBC0;
defparam \Mux12~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N4
cycloneive_lcell_comb \Mux12~20 (
// Equation(s):
// \Mux12~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux12~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux12~19_combout ))

	.dataa(\Mux12~19_combout ),
	.datab(gnd),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux12~9_combout ),
	.cin(gnd),
	.combout(\Mux12~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~20 .lut_mask = 16'hFA0A;
defparam \Mux12~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N12
cycloneive_lcell_comb \Mux11~7 (
// Equation(s):
// \Mux11~7_combout  = (\my_rf.rsel1[2]~input_o  & ((\registerArray[23][20]~q ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\registerArray[19][20]~q  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\registerArray[23][20]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[19][20]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux11~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~7 .lut_mask = 16'hCCB8;
defparam \Mux11~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N30
cycloneive_lcell_comb \Mux11~8 (
// Equation(s):
// \Mux11~8_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux11~7_combout  & (\registerArray[31][20]~q )) # (!\Mux11~7_combout  & ((\registerArray[27][20]~q ))))) # (!\my_rf.rsel1[3]~input_o  & (\Mux11~7_combout ))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux11~7_combout ),
	.datac(\registerArray[31][20]~q ),
	.datad(\registerArray[27][20]~q ),
	.cin(gnd),
	.combout(\Mux11~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~8 .lut_mask = 16'hE6C4;
defparam \Mux11~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y34_N1
dffeas \registerArray[28][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][20] .is_wysiwyg = "true";
defparam \registerArray[28][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N9
dffeas \registerArray[24][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][20] .is_wysiwyg = "true";
defparam \registerArray[24][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N11
dffeas \registerArray[16][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][20] .is_wysiwyg = "true";
defparam \registerArray[16][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N10
cycloneive_lcell_comb \Mux11~4 (
// Equation(s):
// \Mux11~4_combout  = (\my_rf.rsel1[3]~input_o  & ((\registerArray[24][20]~q ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((\registerArray[16][20]~q  & !\my_rf.rsel1[2]~input_o ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\registerArray[24][20]~q ),
	.datac(\registerArray[16][20]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~4 .lut_mask = 16'hAAD8;
defparam \Mux11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N0
cycloneive_lcell_comb \Mux11~5 (
// Equation(s):
// \Mux11~5_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux11~4_combout  & ((\registerArray[28][20]~q ))) # (!\Mux11~4_combout  & (\registerArray[20][20]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux11~4_combout ))))

	.dataa(\registerArray[20][20]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[28][20]~q ),
	.datad(\Mux11~4_combout ),
	.cin(gnd),
	.combout(\Mux11~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~5 .lut_mask = 16'hF388;
defparam \Mux11~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y37_N25
dffeas \registerArray[30][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][20] .is_wysiwyg = "true";
defparam \registerArray[30][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y38_N21
dffeas \registerArray[22][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][20] .is_wysiwyg = "true";
defparam \registerArray[22][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y37_N24
cycloneive_lcell_comb \Mux11~3 (
// Equation(s):
// \Mux11~3_combout  = (\Mux11~2_combout  & (((\registerArray[30][20]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux11~2_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[22][20]~q ))))

	.dataa(\Mux11~2_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[30][20]~q ),
	.datad(\registerArray[22][20]~q ),
	.cin(gnd),
	.combout(\Mux11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~3 .lut_mask = 16'hE6A2;
defparam \Mux11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N18
cycloneive_lcell_comb \Mux11~6 (
// Equation(s):
// \Mux11~6_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\Mux11~3_combout ))) # (!\my_rf.rsel1[1]~input_o  & (\Mux11~5_combout ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux11~5_combout ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\Mux11~3_combout ),
	.cin(gnd),
	.combout(\Mux11~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~6 .lut_mask = 16'hF4A4;
defparam \Mux11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N4
cycloneive_lcell_comb \Mux11~9 (
// Equation(s):
// \Mux11~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux11~6_combout  & ((\Mux11~8_combout ))) # (!\Mux11~6_combout  & (\Mux11~1_combout )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux11~6_combout ))))

	.dataa(\Mux11~1_combout ),
	.datab(\Mux11~8_combout ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\Mux11~6_combout ),
	.cin(gnd),
	.combout(\Mux11~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~9 .lut_mask = 16'hCFA0;
defparam \Mux11~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N27
dffeas \registerArray[15][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][20] .is_wysiwyg = "true";
defparam \registerArray[15][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y35_N1
dffeas \registerArray[14][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][20] .is_wysiwyg = "true";
defparam \registerArray[14][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N26
cycloneive_lcell_comb \Mux11~18 (
// Equation(s):
// \Mux11~18_combout  = (\Mux11~17_combout  & (((\registerArray[15][20]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux11~17_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[14][20]~q ))))

	.dataa(\Mux11~17_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][20]~q ),
	.datad(\registerArray[14][20]~q ),
	.cin(gnd),
	.combout(\Mux11~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~18 .lut_mask = 16'hE6A2;
defparam \Mux11~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y39_N23
dffeas \registerArray[8][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][20] .is_wysiwyg = "true";
defparam \registerArray[8][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N22
cycloneive_lcell_comb \Mux11~10 (
// Equation(s):
// \Mux11~10_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\registerArray[10][20]~q )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & (\registerArray[8][20]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[8][20]~q ),
	.datad(\registerArray[10][20]~q ),
	.cin(gnd),
	.combout(\Mux11~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~10 .lut_mask = 16'hBA98;
defparam \Mux11~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N7
dffeas \registerArray[11][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][20] .is_wysiwyg = "true";
defparam \registerArray[11][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N6
cycloneive_lcell_comb \Mux11~11 (
// Equation(s):
// \Mux11~11_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux11~10_combout  & (\registerArray[11][20]~q )) # (!\Mux11~10_combout  & ((\registerArray[9][20]~q ))))) # (!\my_rf.rsel1[0]~input_o  & (\Mux11~10_combout ))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux11~10_combout ),
	.datac(\registerArray[11][20]~q ),
	.datad(\registerArray[9][20]~q ),
	.cin(gnd),
	.combout(\Mux11~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~11 .lut_mask = 16'hE6C4;
defparam \Mux11~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N31
dffeas \registerArray[2][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][20] .is_wysiwyg = "true";
defparam \registerArray[2][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N4
cycloneive_lcell_comb \Mux11~15 (
// Equation(s):
// \Mux11~15_combout  = (\Mux11~14_combout ) # ((\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & \registerArray[2][20]~q )))

	.dataa(\Mux11~14_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\registerArray[2][20]~q ),
	.cin(gnd),
	.combout(\Mux11~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~15 .lut_mask = 16'hAEAA;
defparam \Mux11~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y31_N28
cycloneive_lcell_comb \Mux11~12 (
// Equation(s):
// \Mux11~12_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[5][20]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[4][20]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[4][20]~q ),
	.datad(\registerArray[5][20]~q ),
	.cin(gnd),
	.combout(\Mux11~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~12 .lut_mask = 16'hDC98;
defparam \Mux11~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y37_N31
dffeas \registerArray[7][20] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[20]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][20] .is_wysiwyg = "true";
defparam \registerArray[7][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N30
cycloneive_lcell_comb \Mux11~13 (
// Equation(s):
// \Mux11~13_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux11~12_combout  & (\registerArray[7][20]~q )) # (!\Mux11~12_combout  & ((\registerArray[6][20]~q ))))) # (!\my_rf.rsel1[1]~input_o  & (\Mux11~12_combout ))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\Mux11~12_combout ),
	.datac(\registerArray[7][20]~q ),
	.datad(\registerArray[6][20]~q ),
	.cin(gnd),
	.combout(\Mux11~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~13 .lut_mask = 16'hE6C4;
defparam \Mux11~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N6
cycloneive_lcell_comb \Mux11~16 (
// Equation(s):
// \Mux11~16_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\Mux11~13_combout ))) # (!\my_rf.rsel1[2]~input_o  & (\Mux11~15_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux11~15_combout ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux11~13_combout ),
	.cin(gnd),
	.combout(\Mux11~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~16 .lut_mask = 16'hF4A4;
defparam \Mux11~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N24
cycloneive_lcell_comb \Mux11~19 (
// Equation(s):
// \Mux11~19_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux11~16_combout  & (\Mux11~18_combout )) # (!\Mux11~16_combout  & ((\Mux11~11_combout ))))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux11~16_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux11~18_combout ),
	.datac(\Mux11~11_combout ),
	.datad(\Mux11~16_combout ),
	.cin(gnd),
	.combout(\Mux11~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~19 .lut_mask = 16'hDDA0;
defparam \Mux11~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N26
cycloneive_lcell_comb \Mux11~20 (
// Equation(s):
// \Mux11~20_combout  = (\my_rf.rsel1[4]~input_o  & (\Mux11~9_combout )) # (!\my_rf.rsel1[4]~input_o  & ((\Mux11~19_combout )))

	.dataa(gnd),
	.datab(\my_rf.rsel1[4]~input_o ),
	.datac(\Mux11~9_combout ),
	.datad(\Mux11~19_combout ),
	.cin(gnd),
	.combout(\Mux11~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~20 .lut_mask = 16'hF3C0;
defparam \Mux11~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y32_N19
dffeas \registerArray[17][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][21] .is_wysiwyg = "true";
defparam \registerArray[17][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y32_N15
dffeas \registerArray[25][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][21] .is_wysiwyg = "true";
defparam \registerArray[25][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N18
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// \Mux10~0_combout  = (\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o ) # ((\registerArray[25][21]~q )))) # (!\my_rf.rsel1[3]~input_o  & (!\my_rf.rsel1[2]~input_o  & (\registerArray[17][21]~q )))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[17][21]~q ),
	.datad(\registerArray[25][21]~q ),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hBA98;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N1
dffeas \registerArray[29][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][21] .is_wysiwyg = "true";
defparam \registerArray[29][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N0
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// \Mux10~1_combout  = (\Mux10~0_combout  & (((\registerArray[29][21]~q ) # (!\my_rf.rsel1[2]~input_o )))) # (!\Mux10~0_combout  & (\registerArray[21][21]~q  & ((\my_rf.rsel1[2]~input_o ))))

	.dataa(\registerArray[21][21]~q ),
	.datab(\Mux10~0_combout ),
	.datac(\registerArray[29][21]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'hE2CC;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y35_N21
dffeas \registerArray[20][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][21] .is_wysiwyg = "true";
defparam \registerArray[20][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y35_N15
dffeas \registerArray[16][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][21] .is_wysiwyg = "true";
defparam \registerArray[16][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N14
cycloneive_lcell_comb \Mux10~4 (
// Equation(s):
// \Mux10~4_combout  = (\my_rf.rsel1[2]~input_o  & ((\registerArray[20][21]~q ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\registerArray[16][21]~q  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[20][21]~q ),
	.datac(\registerArray[16][21]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~4 .lut_mask = 16'hAAD8;
defparam \Mux10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y35_N25
dffeas \registerArray[28][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][21] .is_wysiwyg = "true";
defparam \registerArray[28][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N24
cycloneive_lcell_comb \Mux10~5 (
// Equation(s):
// \Mux10~5_combout  = (\Mux10~4_combout  & (((\registerArray[28][21]~q ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux10~4_combout  & (\registerArray[24][21]~q  & ((\my_rf.rsel1[3]~input_o ))))

	.dataa(\registerArray[24][21]~q ),
	.datab(\Mux10~4_combout ),
	.datac(\registerArray[28][21]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux10~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~5 .lut_mask = 16'hE2CC;
defparam \Mux10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y38_N12
cycloneive_lcell_comb \Mux10~2 (
// Equation(s):
// \Mux10~2_combout  = (\my_rf.rsel1[2]~input_o  & ((\registerArray[22][21]~q ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\registerArray[18][21]~q  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\registerArray[22][21]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][21]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~2 .lut_mask = 16'hCCB8;
defparam \Mux10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y37_N19
dffeas \registerArray[30][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][21] .is_wysiwyg = "true";
defparam \registerArray[30][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y37_N18
cycloneive_lcell_comb \Mux10~3 (
// Equation(s):
// \Mux10~3_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux10~2_combout  & (\registerArray[30][21]~q )) # (!\Mux10~2_combout  & ((\registerArray[26][21]~q ))))) # (!\my_rf.rsel1[3]~input_o  & (\Mux10~2_combout ))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux10~2_combout ),
	.datac(\registerArray[30][21]~q ),
	.datad(\registerArray[26][21]~q ),
	.cin(gnd),
	.combout(\Mux10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~3 .lut_mask = 16'hE6C4;
defparam \Mux10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N16
cycloneive_lcell_comb \Mux10~6 (
// Equation(s):
// \Mux10~6_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\Mux10~3_combout )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & (\Mux10~5_combout )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux10~5_combout ),
	.datad(\Mux10~3_combout ),
	.cin(gnd),
	.combout(\Mux10~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~6 .lut_mask = 16'hBA98;
defparam \Mux10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N26
cycloneive_lcell_comb \Mux10~9 (
// Equation(s):
// \Mux10~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux10~6_combout  & (\Mux10~8_combout )) # (!\Mux10~6_combout  & ((\Mux10~1_combout ))))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux10~6_combout ))))

	.dataa(\Mux10~8_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux10~1_combout ),
	.datad(\Mux10~6_combout ),
	.cin(gnd),
	.combout(\Mux10~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~9 .lut_mask = 16'hBBC0;
defparam \Mux10~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y31_N11
dffeas \registerArray[7][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][21] .is_wysiwyg = "true";
defparam \registerArray[7][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y31_N10
cycloneive_lcell_comb \Mux10~11 (
// Equation(s):
// \Mux10~11_combout  = (\Mux10~10_combout  & (((\registerArray[7][21]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux10~10_combout  & (\registerArray[6][21]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux10~10_combout ),
	.datab(\registerArray[6][21]~q ),
	.datac(\registerArray[7][21]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux10~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~11 .lut_mask = 16'hE4AA;
defparam \Mux10~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N6
cycloneive_lcell_comb \Mux10~18 (
// Equation(s):
// \Mux10~18_combout  = (\Mux10~17_combout  & (((\registerArray[15][21]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux10~17_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[14][21]~q ))))

	.dataa(\Mux10~17_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][21]~q ),
	.datad(\registerArray[14][21]~q ),
	.cin(gnd),
	.combout(\Mux10~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~18 .lut_mask = 16'hE6A2;
defparam \Mux10~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y32_N15
dffeas \registerArray[1][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][21] .is_wysiwyg = "true";
defparam \registerArray[1][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y32_N29
dffeas \registerArray[3][21] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[21]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][21] .is_wysiwyg = "true";
defparam \registerArray[3][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N14
cycloneive_lcell_comb \Mux10~14 (
// Equation(s):
// \Mux10~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][21]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][21]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[1][21]~q ),
	.datad(\registerArray[3][21]~q ),
	.cin(gnd),
	.combout(\Mux10~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~14 .lut_mask = 16'hC840;
defparam \Mux10~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N6
cycloneive_lcell_comb \Mux10~15 (
// Equation(s):
// \Mux10~15_combout  = (\Mux10~14_combout ) # ((\registerArray[2][21]~q  & (!\my_rf.rsel1[0]~input_o  & \my_rf.rsel1[1]~input_o )))

	.dataa(\registerArray[2][21]~q ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux10~14_combout ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux10~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~15 .lut_mask = 16'hF2F0;
defparam \Mux10~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N28
cycloneive_lcell_comb \Mux10~16 (
// Equation(s):
// \Mux10~16_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux10~13_combout ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux10~15_combout  & !\my_rf.rsel1[2]~input_o ))))

	.dataa(\Mux10~13_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\Mux10~15_combout ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux10~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~16 .lut_mask = 16'hCCB8;
defparam \Mux10~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N22
cycloneive_lcell_comb \Mux10~19 (
// Equation(s):
// \Mux10~19_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux10~16_combout  & ((\Mux10~18_combout ))) # (!\Mux10~16_combout  & (\Mux10~11_combout )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux10~16_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux10~11_combout ),
	.datac(\Mux10~18_combout ),
	.datad(\Mux10~16_combout ),
	.cin(gnd),
	.combout(\Mux10~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~19 .lut_mask = 16'hF588;
defparam \Mux10~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N28
cycloneive_lcell_comb \Mux10~20 (
// Equation(s):
// \Mux10~20_combout  = (\my_rf.rsel1[4]~input_o  & (\Mux10~9_combout )) # (!\my_rf.rsel1[4]~input_o  & ((\Mux10~19_combout )))

	.dataa(\Mux10~9_combout ),
	.datab(gnd),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux10~19_combout ),
	.cin(gnd),
	.combout(\Mux10~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~20 .lut_mask = 16'hAFA0;
defparam \Mux10~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y31_N4
cycloneive_lcell_comb \Mux9~13 (
// Equation(s):
// \Mux9~13_combout  = (\Mux9~12_combout  & (((\registerArray[7][22]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux9~12_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[6][22]~q ))))

	.dataa(\Mux9~12_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[7][22]~q ),
	.datad(\registerArray[6][22]~q ),
	.cin(gnd),
	.combout(\Mux9~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~13 .lut_mask = 16'hE6A2;
defparam \Mux9~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N24
cycloneive_lcell_comb \Mux9~16 (
// Equation(s):
// \Mux9~16_combout  = (\my_rf.rsel1[2]~input_o  & (((\Mux9~13_combout ) # (\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (\Mux9~15_combout  & ((!\my_rf.rsel1[3]~input_o ))))

	.dataa(\Mux9~15_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux9~13_combout ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux9~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~16 .lut_mask = 16'hCCE2;
defparam \Mux9~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N30
cycloneive_lcell_comb \Mux9~10 (
// Equation(s):
// \Mux9~10_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\registerArray[10][22]~q )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & (\registerArray[8][22]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[8][22]~q ),
	.datad(\registerArray[10][22]~q ),
	.cin(gnd),
	.combout(\Mux9~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~10 .lut_mask = 16'hBA98;
defparam \Mux9~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N23
dffeas \registerArray[11][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][22] .is_wysiwyg = "true";
defparam \registerArray[11][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N22
cycloneive_lcell_comb \Mux9~11 (
// Equation(s):
// \Mux9~11_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux9~10_combout  & (\registerArray[11][22]~q )) # (!\Mux9~10_combout  & ((\registerArray[9][22]~q ))))) # (!\my_rf.rsel1[0]~input_o  & (\Mux9~10_combout ))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux9~10_combout ),
	.datac(\registerArray[11][22]~q ),
	.datad(\registerArray[9][22]~q ),
	.cin(gnd),
	.combout(\Mux9~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~11 .lut_mask = 16'hE6C4;
defparam \Mux9~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N18
cycloneive_lcell_comb \Mux9~19 (
// Equation(s):
// \Mux9~19_combout  = (\Mux9~16_combout  & ((\Mux9~18_combout ) # ((!\my_rf.rsel1[3]~input_o )))) # (!\Mux9~16_combout  & (((\Mux9~11_combout  & \my_rf.rsel1[3]~input_o ))))

	.dataa(\Mux9~18_combout ),
	.datab(\Mux9~16_combout ),
	.datac(\Mux9~11_combout ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux9~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~19 .lut_mask = 16'hB8CC;
defparam \Mux9~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y33_N21
dffeas \registerArray[31][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][22] .is_wysiwyg = "true";
defparam \registerArray[31][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N20
cycloneive_lcell_comb \Mux9~8 (
// Equation(s):
// \Mux9~8_combout  = (\Mux9~7_combout  & (((\registerArray[31][22]~q ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux9~7_combout  & (\registerArray[27][22]~q  & ((\my_rf.rsel1[3]~input_o ))))

	.dataa(\Mux9~7_combout ),
	.datab(\registerArray[27][22]~q ),
	.datac(\registerArray[31][22]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux9~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~8 .lut_mask = 16'hE4AA;
defparam \Mux9~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N23
dffeas \registerArray[17][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][22] .is_wysiwyg = "true";
defparam \registerArray[17][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N22
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// \Mux9~0_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & (\registerArray[21][22]~q )) # (!\my_rf.rsel1[2]~input_o  & ((\registerArray[17][22]~q )))))

	.dataa(\registerArray[21][22]~q ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[17][22]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hEE30;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y36_N29
dffeas \registerArray[29][22] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[22]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][22] .is_wysiwyg = "true";
defparam \registerArray[29][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N28
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// \Mux9~1_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux9~0_combout  & (\registerArray[29][22]~q )) # (!\Mux9~0_combout  & ((\registerArray[25][22]~q ))))) # (!\my_rf.rsel1[3]~input_o  & (\Mux9~0_combout ))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux9~0_combout ),
	.datac(\registerArray[29][22]~q ),
	.datad(\registerArray[25][22]~q ),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'hE6C4;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N12
cycloneive_lcell_comb \Mux9~9 (
// Equation(s):
// \Mux9~9_combout  = (\Mux9~6_combout  & (((\Mux9~8_combout )) # (!\my_rf.rsel1[0]~input_o ))) # (!\Mux9~6_combout  & (\my_rf.rsel1[0]~input_o  & ((\Mux9~1_combout ))))

	.dataa(\Mux9~6_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux9~8_combout ),
	.datad(\Mux9~1_combout ),
	.cin(gnd),
	.combout(\Mux9~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~9 .lut_mask = 16'hE6A2;
defparam \Mux9~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N28
cycloneive_lcell_comb \Mux9~20 (
// Equation(s):
// \Mux9~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux9~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux9~19_combout ))

	.dataa(gnd),
	.datab(\Mux9~19_combout ),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux9~9_combout ),
	.cin(gnd),
	.combout(\Mux9~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~20 .lut_mask = 16'hFC0C;
defparam \Mux9~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N10
cycloneive_lcell_comb \Mux8~18 (
// Equation(s):
// \Mux8~18_combout  = (\Mux8~17_combout  & (((\registerArray[15][23]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux8~17_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[14][23]~q ))))

	.dataa(\Mux8~17_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][23]~q ),
	.datad(\registerArray[14][23]~q ),
	.cin(gnd),
	.combout(\Mux8~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~18 .lut_mask = 16'hE6A2;
defparam \Mux8~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y39_N25
dffeas \registerArray[9][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][23] .is_wysiwyg = "true";
defparam \registerArray[9][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y39_N27
dffeas \registerArray[11][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][23] .is_wysiwyg = "true";
defparam \registerArray[11][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y39_N11
dffeas \registerArray[8][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][23] .is_wysiwyg = "true";
defparam \registerArray[8][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y39_N1
dffeas \registerArray[10][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][23] .is_wysiwyg = "true";
defparam \registerArray[10][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y39_N10
cycloneive_lcell_comb \Mux8~12 (
// Equation(s):
// \Mux8~12_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\registerArray[10][23]~q )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & (\registerArray[8][23]~q )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[8][23]~q ),
	.datad(\registerArray[10][23]~q ),
	.cin(gnd),
	.combout(\Mux8~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~12 .lut_mask = 16'hBA98;
defparam \Mux8~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y39_N26
cycloneive_lcell_comb \Mux8~13 (
// Equation(s):
// \Mux8~13_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux8~12_combout  & ((\registerArray[11][23]~q ))) # (!\Mux8~12_combout  & (\registerArray[9][23]~q )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux8~12_combout ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\registerArray[9][23]~q ),
	.datac(\registerArray[11][23]~q ),
	.datad(\Mux8~12_combout ),
	.cin(gnd),
	.combout(\Mux8~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~13 .lut_mask = 16'hF588;
defparam \Mux8~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N16
cycloneive_lcell_comb \Mux8~16 (
// Equation(s):
// \Mux8~16_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & ((\Mux8~13_combout ))) # (!\my_rf.rsel1[3]~input_o  & (\Mux8~15_combout ))))

	.dataa(\Mux8~15_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux8~13_combout ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux8~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~16 .lut_mask = 16'hFC22;
defparam \Mux8~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y38_N26
cycloneive_lcell_comb \Mux8~19 (
// Equation(s):
// \Mux8~19_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux8~16_combout  & ((\Mux8~18_combout ))) # (!\Mux8~16_combout  & (\Mux8~11_combout )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux8~16_combout ))))

	.dataa(\Mux8~11_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux8~18_combout ),
	.datad(\Mux8~16_combout ),
	.cin(gnd),
	.combout(\Mux8~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~19 .lut_mask = 16'hF388;
defparam \Mux8~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y37_N15
dffeas \registerArray[30][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][23] .is_wysiwyg = "true";
defparam \registerArray[30][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y37_N21
dffeas \registerArray[26][23] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[23]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][23] .is_wysiwyg = "true";
defparam \registerArray[26][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y37_N14
cycloneive_lcell_comb \Mux8~3 (
// Equation(s):
// \Mux8~3_combout  = (\Mux8~2_combout  & (((\registerArray[30][23]~q )) # (!\my_rf.rsel1[3]~input_o ))) # (!\Mux8~2_combout  & (\my_rf.rsel1[3]~input_o  & ((\registerArray[26][23]~q ))))

	.dataa(\Mux8~2_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[30][23]~q ),
	.datad(\registerArray[26][23]~q ),
	.cin(gnd),
	.combout(\Mux8~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~3 .lut_mask = 16'hE6A2;
defparam \Mux8~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N6
cycloneive_lcell_comb \Mux8~6 (
// Equation(s):
// \Mux8~6_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\Mux8~3_combout ))) # (!\my_rf.rsel1[1]~input_o  & (\Mux8~5_combout ))))

	.dataa(\Mux8~5_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\Mux8~3_combout ),
	.cin(gnd),
	.combout(\Mux8~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~6 .lut_mask = 16'hF2C2;
defparam \Mux8~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N2
cycloneive_lcell_comb \Mux8~7 (
// Equation(s):
// \Mux8~7_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[27][23]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[19][23]~q )))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[27][23]~q ),
	.datac(\registerArray[19][23]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux8~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~7 .lut_mask = 16'hEE50;
defparam \Mux8~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y33_N8
cycloneive_lcell_comb \Mux8~8 (
// Equation(s):
// \Mux8~8_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux8~7_combout  & ((\registerArray[31][23]~q ))) # (!\Mux8~7_combout  & (\registerArray[23][23]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux8~7_combout ))))

	.dataa(\registerArray[23][23]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[31][23]~q ),
	.datad(\Mux8~7_combout ),
	.cin(gnd),
	.combout(\Mux8~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~8 .lut_mask = 16'hF388;
defparam \Mux8~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N0
cycloneive_lcell_comb \Mux8~9 (
// Equation(s):
// \Mux8~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux8~6_combout  & ((\Mux8~8_combout ))) # (!\Mux8~6_combout  & (\Mux8~1_combout )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux8~6_combout ))))

	.dataa(\Mux8~1_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux8~6_combout ),
	.datad(\Mux8~8_combout ),
	.cin(gnd),
	.combout(\Mux8~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~9 .lut_mask = 16'hF838;
defparam \Mux8~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N10
cycloneive_lcell_comb \Mux8~20 (
// Equation(s):
// \Mux8~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux8~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux8~19_combout ))

	.dataa(gnd),
	.datab(\Mux8~19_combout ),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux8~9_combout ),
	.cin(gnd),
	.combout(\Mux8~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~20 .lut_mask = 16'hFC0C;
defparam \Mux8~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y36_N29
dffeas \registerArray[14][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][24] .is_wysiwyg = "true";
defparam \registerArray[14][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y36_N23
dffeas \registerArray[15][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][24] .is_wysiwyg = "true";
defparam \registerArray[15][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y36_N22
cycloneive_lcell_comb \Mux7~18 (
// Equation(s):
// \Mux7~18_combout  = (\Mux7~17_combout  & (((\registerArray[15][24]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux7~17_combout  & (\registerArray[14][24]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux7~17_combout ),
	.datab(\registerArray[14][24]~q ),
	.datac(\registerArray[15][24]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux7~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~18 .lut_mask = 16'hE4AA;
defparam \Mux7~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y33_N2
cycloneive_lcell_comb \Mux7~11 (
// Equation(s):
// \Mux7~11_combout  = (\Mux7~10_combout  & (((\registerArray[11][24]~q )) # (!\my_rf.rsel1[0]~input_o ))) # (!\Mux7~10_combout  & (\my_rf.rsel1[0]~input_o  & ((\registerArray[9][24]~q ))))

	.dataa(\Mux7~10_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[11][24]~q ),
	.datad(\registerArray[9][24]~q ),
	.cin(gnd),
	.combout(\Mux7~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~11 .lut_mask = 16'hE6A2;
defparam \Mux7~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y34_N11
dffeas \registerArray[1][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][24] .is_wysiwyg = "true";
defparam \registerArray[1][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y34_N1
dffeas \registerArray[3][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][24] .is_wysiwyg = "true";
defparam \registerArray[3][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N10
cycloneive_lcell_comb \Mux7~14 (
// Equation(s):
// \Mux7~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][24]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][24]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[1][24]~q ),
	.datad(\registerArray[3][24]~q ),
	.cin(gnd),
	.combout(\Mux7~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~14 .lut_mask = 16'hA820;
defparam \Mux7~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N21
dffeas \registerArray[2][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][24] .is_wysiwyg = "true";
defparam \registerArray[2][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N14
cycloneive_lcell_comb \Mux7~15 (
// Equation(s):
// \Mux7~15_combout  = (\Mux7~14_combout ) # ((!\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o  & \registerArray[2][24]~q )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux7~14_combout ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\registerArray[2][24]~q ),
	.cin(gnd),
	.combout(\Mux7~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~15 .lut_mask = 16'hDCCC;
defparam \Mux7~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N11
dffeas \registerArray[7][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][24] .is_wysiwyg = "true";
defparam \registerArray[7][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N10
cycloneive_lcell_comb \Mux7~13 (
// Equation(s):
// \Mux7~13_combout  = (\Mux7~12_combout  & (((\registerArray[7][24]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux7~12_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[6][24]~q ))))

	.dataa(\Mux7~12_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[7][24]~q ),
	.datad(\registerArray[6][24]~q ),
	.cin(gnd),
	.combout(\Mux7~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~13 .lut_mask = 16'hE6A2;
defparam \Mux7~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N16
cycloneive_lcell_comb \Mux7~16 (
// Equation(s):
// \Mux7~16_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\Mux7~13_combout ))) # (!\my_rf.rsel1[2]~input_o  & (\Mux7~15_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux7~15_combout ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux7~13_combout ),
	.cin(gnd),
	.combout(\Mux7~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~16 .lut_mask = 16'hF4A4;
defparam \Mux7~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N10
cycloneive_lcell_comb \Mux7~19 (
// Equation(s):
// \Mux7~19_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux7~16_combout  & (\Mux7~18_combout )) # (!\Mux7~16_combout  & ((\Mux7~11_combout ))))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux7~16_combout ))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux7~18_combout ),
	.datac(\Mux7~11_combout ),
	.datad(\Mux7~16_combout ),
	.cin(gnd),
	.combout(\Mux7~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~19 .lut_mask = 16'hDDA0;
defparam \Mux7~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N9
dffeas \registerArray[21][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][24] .is_wysiwyg = "true";
defparam \registerArray[21][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N19
dffeas \registerArray[17][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][24] .is_wysiwyg = "true";
defparam \registerArray[17][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N18
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (\my_rf.rsel1[2]~input_o  & ((\registerArray[21][24]~q ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\registerArray[17][24]~q  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[21][24]~q ),
	.datac(\registerArray[17][24]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hAAD8;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N0
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// \Mux7~1_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux7~0_combout  & ((\registerArray[29][24]~q ))) # (!\Mux7~0_combout  & (\registerArray[25][24]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux7~0_combout ))))

	.dataa(\registerArray[25][24]~q ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[29][24]~q ),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hF388;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y33_N13
dffeas \registerArray[27][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][24] .is_wysiwyg = "true";
defparam \registerArray[27][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y33_N5
dffeas \registerArray[31][24] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[24]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][24] .is_wysiwyg = "true";
defparam \registerArray[31][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N4
cycloneive_lcell_comb \Mux7~8 (
// Equation(s):
// \Mux7~8_combout  = (\Mux7~7_combout  & (((\registerArray[31][24]~q ) # (!\my_rf.rsel1[3]~input_o )))) # (!\Mux7~7_combout  & (\registerArray[27][24]~q  & ((\my_rf.rsel1[3]~input_o ))))

	.dataa(\Mux7~7_combout ),
	.datab(\registerArray[27][24]~q ),
	.datac(\registerArray[31][24]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux7~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~8 .lut_mask = 16'hE4AA;
defparam \Mux7~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N20
cycloneive_lcell_comb \Mux7~9 (
// Equation(s):
// \Mux7~9_combout  = (\Mux7~6_combout  & (((\Mux7~8_combout ) # (!\my_rf.rsel1[0]~input_o )))) # (!\Mux7~6_combout  & (\Mux7~1_combout  & (\my_rf.rsel1[0]~input_o )))

	.dataa(\Mux7~6_combout ),
	.datab(\Mux7~1_combout ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\Mux7~8_combout ),
	.cin(gnd),
	.combout(\Mux7~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~9 .lut_mask = 16'hEA4A;
defparam \Mux7~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N28
cycloneive_lcell_comb \Mux7~20 (
// Equation(s):
// \Mux7~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux7~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux7~19_combout ))

	.dataa(\Mux7~19_combout ),
	.datab(\my_rf.rsel1[4]~input_o ),
	.datac(gnd),
	.datad(\Mux7~9_combout ),
	.cin(gnd),
	.combout(\Mux7~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~20 .lut_mask = 16'hEE22;
defparam \Mux7~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N23
dffeas \registerArray[7][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][25] .is_wysiwyg = "true";
defparam \registerArray[7][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N22
cycloneive_lcell_comb \Mux6~11 (
// Equation(s):
// \Mux6~11_combout  = (\Mux6~10_combout  & (((\registerArray[7][25]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux6~10_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[6][25]~q ))))

	.dataa(\Mux6~10_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[7][25]~q ),
	.datad(\registerArray[6][25]~q ),
	.cin(gnd),
	.combout(\Mux6~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~11 .lut_mask = 16'hE6A2;
defparam \Mux6~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N14
cycloneive_lcell_comb \Mux6~14 (
// Equation(s):
// \Mux6~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][25]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][25]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[1][25]~q ),
	.datad(\registerArray[3][25]~q ),
	.cin(gnd),
	.combout(\Mux6~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~14 .lut_mask = 16'hA820;
defparam \Mux6~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y38_N22
cycloneive_lcell_comb \Mux6~15 (
// Equation(s):
// \Mux6~15_combout  = (\Mux6~14_combout ) # ((\my_rf.rsel1[1]~input_o  & (\registerArray[2][25]~q  & !\my_rf.rsel1[0]~input_o )))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[2][25]~q ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\Mux6~14_combout ),
	.cin(gnd),
	.combout(\Mux6~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~15 .lut_mask = 16'hFF08;
defparam \Mux6~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y38_N16
cycloneive_lcell_comb \Mux6~16 (
// Equation(s):
// \Mux6~16_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux6~13_combout ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux6~15_combout  & !\my_rf.rsel1[2]~input_o ))))

	.dataa(\Mux6~13_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\Mux6~15_combout ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux6~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~16 .lut_mask = 16'hCCB8;
defparam \Mux6~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y38_N26
cycloneive_lcell_comb \Mux6~19 (
// Equation(s):
// \Mux6~19_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux6~16_combout  & (\Mux6~18_combout )) # (!\Mux6~16_combout  & ((\Mux6~11_combout ))))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux6~16_combout ))))

	.dataa(\Mux6~18_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux6~11_combout ),
	.datad(\Mux6~16_combout ),
	.cin(gnd),
	.combout(\Mux6~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~19 .lut_mask = 16'hBBC0;
defparam \Mux6~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y32_N31
dffeas \registerArray[23][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][25] .is_wysiwyg = "true";
defparam \registerArray[23][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y33_N27
dffeas \registerArray[31][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][25] .is_wysiwyg = "true";
defparam \registerArray[31][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N15
dffeas \registerArray[27][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][25] .is_wysiwyg = "true";
defparam \registerArray[27][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N1
dffeas \registerArray[19][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][25] .is_wysiwyg = "true";
defparam \registerArray[19][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N0
cycloneive_lcell_comb \Mux6~7 (
// Equation(s):
// \Mux6~7_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[27][25]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[19][25]~q )))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[27][25]~q ),
	.datac(\registerArray[19][25]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux6~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~7 .lut_mask = 16'hEE50;
defparam \Mux6~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N26
cycloneive_lcell_comb \Mux6~8 (
// Equation(s):
// \Mux6~8_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux6~7_combout  & ((\registerArray[31][25]~q ))) # (!\Mux6~7_combout  & (\registerArray[23][25]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux6~7_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[23][25]~q ),
	.datac(\registerArray[31][25]~q ),
	.datad(\Mux6~7_combout ),
	.cin(gnd),
	.combout(\Mux6~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~8 .lut_mask = 16'hF588;
defparam \Mux6~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N20
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// \Mux6~0_combout  = (\my_rf.rsel1[2]~input_o  & (\my_rf.rsel1[3]~input_o )) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & ((\registerArray[25][25]~q ))) # (!\my_rf.rsel1[3]~input_o  & (\registerArray[17][25]~q ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[17][25]~q ),
	.datad(\registerArray[25][25]~q ),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'hDC98;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X0_Y33_N24
dffeas \registerArray[21][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[25]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][25] .is_wysiwyg = "true";
defparam \registerArray[21][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N22
cycloneive_lcell_comb \Mux6~1 (
// Equation(s):
// \Mux6~1_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux6~0_combout  & (\registerArray[29][25]~q )) # (!\Mux6~0_combout  & ((\registerArray[21][25]~q ))))) # (!\my_rf.rsel1[2]~input_o  & (\Mux6~0_combout ))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux6~0_combout ),
	.datac(\registerArray[29][25]~q ),
	.datad(\registerArray[21][25]~q ),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~1 .lut_mask = 16'hE6C4;
defparam \Mux6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y38_N19
dffeas \registerArray[30][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][25] .is_wysiwyg = "true";
defparam \registerArray[30][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y38_N18
cycloneive_lcell_comb \Mux6~3 (
// Equation(s):
// \Mux6~3_combout  = (\Mux6~2_combout  & (((\registerArray[30][25]~q )) # (!\my_rf.rsel1[3]~input_o ))) # (!\Mux6~2_combout  & (\my_rf.rsel1[3]~input_o  & ((\registerArray[26][25]~q ))))

	.dataa(\Mux6~2_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[30][25]~q ),
	.datad(\registerArray[26][25]~q ),
	.cin(gnd),
	.combout(\Mux6~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~3 .lut_mask = 16'hE6A2;
defparam \Mux6~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y35_N9
dffeas \registerArray[28][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][25] .is_wysiwyg = "true";
defparam \registerArray[28][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N3
dffeas \registerArray[24][25] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[25]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][25] .is_wysiwyg = "true";
defparam \registerArray[24][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N8
cycloneive_lcell_comb \Mux6~5 (
// Equation(s):
// \Mux6~5_combout  = (\Mux6~4_combout  & (((\registerArray[28][25]~q )) # (!\my_rf.rsel1[3]~input_o ))) # (!\Mux6~4_combout  & (\my_rf.rsel1[3]~input_o  & ((\registerArray[24][25]~q ))))

	.dataa(\Mux6~4_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[28][25]~q ),
	.datad(\registerArray[24][25]~q ),
	.cin(gnd),
	.combout(\Mux6~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~5 .lut_mask = 16'hE6A2;
defparam \Mux6~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y38_N10
cycloneive_lcell_comb \Mux6~6 (
// Equation(s):
// \Mux6~6_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux6~3_combout ) # ((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & (((!\my_rf.rsel1[0]~input_o  & \Mux6~5_combout ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\Mux6~3_combout ),
	.datac(\my_rf.rsel1[0]~input_o ),
	.datad(\Mux6~5_combout ),
	.cin(gnd),
	.combout(\Mux6~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~6 .lut_mask = 16'hADA8;
defparam \Mux6~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y38_N12
cycloneive_lcell_comb \Mux6~9 (
// Equation(s):
// \Mux6~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux6~6_combout  & (\Mux6~8_combout )) # (!\Mux6~6_combout  & ((\Mux6~1_combout ))))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux6~6_combout ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux6~8_combout ),
	.datac(\Mux6~1_combout ),
	.datad(\Mux6~6_combout ),
	.cin(gnd),
	.combout(\Mux6~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~9 .lut_mask = 16'hDDA0;
defparam \Mux6~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y38_N20
cycloneive_lcell_comb \Mux6~20 (
// Equation(s):
// \Mux6~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux6~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux6~19_combout ))

	.dataa(gnd),
	.datab(\Mux6~19_combout ),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux6~9_combout ),
	.cin(gnd),
	.combout(\Mux6~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~20 .lut_mask = 16'hFC0C;
defparam \Mux6~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y34_N27
dffeas \registerArray[15][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][26] .is_wysiwyg = "true";
defparam \registerArray[15][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y34_N26
cycloneive_lcell_comb \Mux5~18 (
// Equation(s):
// \Mux5~18_combout  = (\Mux5~17_combout  & (((\registerArray[15][26]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux5~17_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[14][26]~q ))))

	.dataa(\Mux5~17_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][26]~q ),
	.datad(\registerArray[14][26]~q ),
	.cin(gnd),
	.combout(\Mux5~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~18 .lut_mask = 16'hE6A2;
defparam \Mux5~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N7
dffeas \registerArray[7][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][26] .is_wysiwyg = "true";
defparam \registerArray[7][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N6
cycloneive_lcell_comb \Mux5~13 (
// Equation(s):
// \Mux5~13_combout  = (\Mux5~12_combout  & (((\registerArray[7][26]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux5~12_combout  & (\registerArray[6][26]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux5~12_combout ),
	.datab(\registerArray[6][26]~q ),
	.datac(\registerArray[7][26]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux5~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~13 .lut_mask = 16'hE4AA;
defparam \Mux5~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N16
cycloneive_lcell_comb \Mux5~14 (
// Equation(s):
// \Mux5~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][26]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][26]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[1][26]~q ),
	.datad(\registerArray[3][26]~q ),
	.cin(gnd),
	.combout(\Mux5~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~14 .lut_mask = 16'hA820;
defparam \Mux5~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N24
cycloneive_lcell_comb \Mux5~15 (
// Equation(s):
// \Mux5~15_combout  = (\Mux5~14_combout ) # ((!\my_rf.rsel1[0]~input_o  & (\registerArray[2][26]~q  & \my_rf.rsel1[1]~input_o )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux5~14_combout ),
	.datac(\registerArray[2][26]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux5~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~15 .lut_mask = 16'hDCCC;
defparam \Mux5~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N18
cycloneive_lcell_comb \Mux5~16 (
// Equation(s):
// \Mux5~16_combout  = (\my_rf.rsel1[3]~input_o  & (\my_rf.rsel1[2]~input_o )) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & (\Mux5~13_combout )) # (!\my_rf.rsel1[2]~input_o  & ((\Mux5~15_combout )))))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux5~13_combout ),
	.datad(\Mux5~15_combout ),
	.cin(gnd),
	.combout(\Mux5~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~16 .lut_mask = 16'hD9C8;
defparam \Mux5~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N4
cycloneive_lcell_comb \Mux5~19 (
// Equation(s):
// \Mux5~19_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux5~16_combout  & ((\Mux5~18_combout ))) # (!\Mux5~16_combout  & (\Mux5~11_combout )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux5~16_combout ))))

	.dataa(\Mux5~11_combout ),
	.datab(\Mux5~18_combout ),
	.datac(\my_rf.rsel1[3]~input_o ),
	.datad(\Mux5~16_combout ),
	.cin(gnd),
	.combout(\Mux5~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~19 .lut_mask = 16'hCFA0;
defparam \Mux5~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y35_N21
dffeas \registerArray[28][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][26] .is_wysiwyg = "true";
defparam \registerArray[28][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y35_N27
dffeas \registerArray[20][26] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[26]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][26] .is_wysiwyg = "true";
defparam \registerArray[20][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N20
cycloneive_lcell_comb \Mux5~5 (
// Equation(s):
// \Mux5~5_combout  = (\Mux5~4_combout  & (((\registerArray[28][26]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux5~4_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[20][26]~q ))))

	.dataa(\Mux5~4_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[28][26]~q ),
	.datad(\registerArray[20][26]~q ),
	.cin(gnd),
	.combout(\Mux5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~5 .lut_mask = 16'hE6A2;
defparam \Mux5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N14
cycloneive_lcell_comb \Mux5~6 (
// Equation(s):
// \Mux5~6_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\Mux5~3_combout )) # (!\my_rf.rsel1[1]~input_o  & ((\Mux5~5_combout )))))

	.dataa(\Mux5~3_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux5~5_combout ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux5~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~6 .lut_mask = 16'hEE30;
defparam \Mux5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N12
cycloneive_lcell_comb \Mux5~8 (
// Equation(s):
// \Mux5~8_combout  = (\Mux5~7_combout  & (((\registerArray[31][26]~q )) # (!\my_rf.rsel1[3]~input_o ))) # (!\Mux5~7_combout  & (\my_rf.rsel1[3]~input_o  & ((\registerArray[27][26]~q ))))

	.dataa(\Mux5~7_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[31][26]~q ),
	.datad(\registerArray[27][26]~q ),
	.cin(gnd),
	.combout(\Mux5~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~8 .lut_mask = 16'hE6A2;
defparam \Mux5~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N0
cycloneive_lcell_comb \Mux5~9 (
// Equation(s):
// \Mux5~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux5~6_combout  & ((\Mux5~8_combout ))) # (!\Mux5~6_combout  & (\Mux5~1_combout )))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux5~6_combout ))))

	.dataa(\Mux5~1_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux5~6_combout ),
	.datad(\Mux5~8_combout ),
	.cin(gnd),
	.combout(\Mux5~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~9 .lut_mask = 16'hF838;
defparam \Mux5~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N30
cycloneive_lcell_comb \Mux5~20 (
// Equation(s):
// \Mux5~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux5~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux5~19_combout ))

	.dataa(gnd),
	.datab(\Mux5~19_combout ),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux5~9_combout ),
	.cin(gnd),
	.combout(\Mux5~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~20 .lut_mask = 16'hFC0C;
defparam \Mux5~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N3
dffeas \registerArray[17][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][27] .is_wysiwyg = "true";
defparam \registerArray[17][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N2
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// \Mux4~0_combout  = (\my_rf.rsel1[3]~input_o  & ((\registerArray[25][27]~q ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((\registerArray[17][27]~q  & !\my_rf.rsel1[2]~input_o ))))

	.dataa(\registerArray[25][27]~q ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[17][27]~q ),
	.datad(\my_rf.rsel1[2]~input_o ),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'hCCB8;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N30
cycloneive_lcell_comb \Mux4~1 (
// Equation(s):
// \Mux4~1_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux4~0_combout  & ((\registerArray[29][27]~q ))) # (!\Mux4~0_combout  & (\registerArray[21][27]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux4~0_combout ))))

	.dataa(\registerArray[21][27]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[29][27]~q ),
	.datad(\Mux4~0_combout ),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~1 .lut_mask = 16'hF388;
defparam \Mux4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y32_N27
dffeas \registerArray[23][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][27] .is_wysiwyg = "true";
defparam \registerArray[23][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y33_N3
dffeas \registerArray[31][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][27] .is_wysiwyg = "true";
defparam \registerArray[31][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y31_N9
dffeas \registerArray[19][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][27] .is_wysiwyg = "true";
defparam \registerArray[19][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N31
dffeas \registerArray[27][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~20_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][27] .is_wysiwyg = "true";
defparam \registerArray[27][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N8
cycloneive_lcell_comb \Mux4~7 (
// Equation(s):
// \Mux4~7_combout  = (\my_rf.rsel1[2]~input_o  & (\my_rf.rsel1[3]~input_o )) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & ((\registerArray[27][27]~q ))) # (!\my_rf.rsel1[3]~input_o  & (\registerArray[19][27]~q ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[19][27]~q ),
	.datad(\registerArray[27][27]~q ),
	.cin(gnd),
	.combout(\Mux4~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~7 .lut_mask = 16'hDC98;
defparam \Mux4~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N2
cycloneive_lcell_comb \Mux4~8 (
// Equation(s):
// \Mux4~8_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux4~7_combout  & ((\registerArray[31][27]~q ))) # (!\Mux4~7_combout  & (\registerArray[23][27]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux4~7_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[23][27]~q ),
	.datac(\registerArray[31][27]~q ),
	.datad(\Mux4~7_combout ),
	.cin(gnd),
	.combout(\Mux4~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~8 .lut_mask = 16'hF588;
defparam \Mux4~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N12
cycloneive_lcell_comb \Mux4~9 (
// Equation(s):
// \Mux4~9_combout  = (\Mux4~6_combout  & (((\Mux4~8_combout )) # (!\my_rf.rsel1[0]~input_o ))) # (!\Mux4~6_combout  & (\my_rf.rsel1[0]~input_o  & (\Mux4~1_combout )))

	.dataa(\Mux4~6_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux4~1_combout ),
	.datad(\Mux4~8_combout ),
	.cin(gnd),
	.combout(\Mux4~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~9 .lut_mask = 16'hEA62;
defparam \Mux4~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y34_N5
dffeas \registerArray[13][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][27] .is_wysiwyg = "true";
defparam \registerArray[13][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y34_N23
dffeas \registerArray[12][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][27] .is_wysiwyg = "true";
defparam \registerArray[12][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N22
cycloneive_lcell_comb \Mux4~17 (
// Equation(s):
// \Mux4~17_combout  = (\my_rf.rsel1[1]~input_o  & (((\my_rf.rsel1[0]~input_o )))) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & (\registerArray[13][27]~q )) # (!\my_rf.rsel1[0]~input_o  & ((\registerArray[12][27]~q )))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\registerArray[13][27]~q ),
	.datac(\registerArray[12][27]~q ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux4~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~17 .lut_mask = 16'hEE50;
defparam \Mux4~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y34_N14
cycloneive_lcell_comb \Mux4~18 (
// Equation(s):
// \Mux4~18_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux4~17_combout  & ((\registerArray[15][27]~q ))) # (!\Mux4~17_combout  & (\registerArray[14][27]~q )))) # (!\my_rf.rsel1[1]~input_o  & (((\Mux4~17_combout ))))

	.dataa(\registerArray[14][27]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][27]~q ),
	.datad(\Mux4~17_combout ),
	.cin(gnd),
	.combout(\Mux4~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~18 .lut_mask = 16'hF388;
defparam \Mux4~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N22
cycloneive_lcell_comb \Mux4~14 (
// Equation(s):
// \Mux4~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & ((\registerArray[3][27]~q ))) # (!\my_rf.rsel1[1]~input_o  & (\registerArray[1][27]~q ))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[1][27]~q ),
	.datad(\registerArray[3][27]~q ),
	.cin(gnd),
	.combout(\Mux4~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~14 .lut_mask = 16'hA820;
defparam \Mux4~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N26
cycloneive_lcell_comb \Mux4~15 (
// Equation(s):
// \Mux4~15_combout  = (\Mux4~14_combout ) # ((!\my_rf.rsel1[0]~input_o  & (\registerArray[2][27]~q  & \my_rf.rsel1[1]~input_o )))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\Mux4~14_combout ),
	.datac(\registerArray[2][27]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux4~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~15 .lut_mask = 16'hDCCC;
defparam \Mux4~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N14
cycloneive_lcell_comb \Mux4~16 (
// Equation(s):
// \Mux4~16_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux4~13_combout ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((!\my_rf.rsel1[2]~input_o  & \Mux4~15_combout ))))

	.dataa(\Mux4~13_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux4~15_combout ),
	.cin(gnd),
	.combout(\Mux4~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~16 .lut_mask = 16'hCBC8;
defparam \Mux4~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N31
dffeas \registerArray[4][27] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[27]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][27] .is_wysiwyg = "true";
defparam \registerArray[4][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N30
cycloneive_lcell_comb \Mux4~10 (
// Equation(s):
// \Mux4~10_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[5][27]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[4][27]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[4][27]~q ),
	.datad(\registerArray[5][27]~q ),
	.cin(gnd),
	.combout(\Mux4~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~10 .lut_mask = 16'hDC98;
defparam \Mux4~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N2
cycloneive_lcell_comb \Mux4~11 (
// Equation(s):
// \Mux4~11_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux4~10_combout  & (\registerArray[7][27]~q )) # (!\Mux4~10_combout  & ((\registerArray[6][27]~q ))))) # (!\my_rf.rsel1[1]~input_o  & (\Mux4~10_combout ))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\Mux4~10_combout ),
	.datac(\registerArray[7][27]~q ),
	.datad(\registerArray[6][27]~q ),
	.cin(gnd),
	.combout(\Mux4~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~11 .lut_mask = 16'hE6C4;
defparam \Mux4~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N0
cycloneive_lcell_comb \Mux4~19 (
// Equation(s):
// \Mux4~19_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux4~16_combout  & (\Mux4~18_combout )) # (!\Mux4~16_combout  & ((\Mux4~11_combout ))))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux4~16_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux4~18_combout ),
	.datac(\Mux4~16_combout ),
	.datad(\Mux4~11_combout ),
	.cin(gnd),
	.combout(\Mux4~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~19 .lut_mask = 16'hDAD0;
defparam \Mux4~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N18
cycloneive_lcell_comb \Mux4~20 (
// Equation(s):
// \Mux4~20_combout  = (\my_rf.rsel1[4]~input_o  & (\Mux4~9_combout )) # (!\my_rf.rsel1[4]~input_o  & ((\Mux4~19_combout )))

	.dataa(\Mux4~9_combout ),
	.datab(\my_rf.rsel1[4]~input_o ),
	.datac(gnd),
	.datad(\Mux4~19_combout ),
	.cin(gnd),
	.combout(\Mux4~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~20 .lut_mask = 16'hBB88;
defparam \Mux4~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y37_N9
dffeas \registerArray[22][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][28] .is_wysiwyg = "true";
defparam \registerArray[22][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y35_N15
dffeas \registerArray[30][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][28] .is_wysiwyg = "true";
defparam \registerArray[30][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y37_N19
dffeas \registerArray[18][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][28] .is_wysiwyg = "true";
defparam \registerArray[18][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y36_N1
dffeas \registerArray[26][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][28] .is_wysiwyg = "true";
defparam \registerArray[26][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y37_N18
cycloneive_lcell_comb \Mux3~2 (
// Equation(s):
// \Mux3~2_combout  = (\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o ) # ((\registerArray[26][28]~q )))) # (!\my_rf.rsel1[3]~input_o  & (!\my_rf.rsel1[2]~input_o  & (\registerArray[18][28]~q )))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[18][28]~q ),
	.datad(\registerArray[26][28]~q ),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~2 .lut_mask = 16'hBA98;
defparam \Mux3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N14
cycloneive_lcell_comb \Mux3~3 (
// Equation(s):
// \Mux3~3_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux3~2_combout  & ((\registerArray[30][28]~q ))) # (!\Mux3~2_combout  & (\registerArray[22][28]~q )))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux3~2_combout ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[22][28]~q ),
	.datac(\registerArray[30][28]~q ),
	.datad(\Mux3~2_combout ),
	.cin(gnd),
	.combout(\Mux3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~3 .lut_mask = 16'hF588;
defparam \Mux3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N12
cycloneive_lcell_comb \Mux3~4 (
// Equation(s):
// \Mux3~4_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[24][28]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[16][28]~q )))))

	.dataa(\registerArray[24][28]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[16][28]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~4 .lut_mask = 16'hEE30;
defparam \Mux3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N16
cycloneive_lcell_comb \Mux3~5 (
// Equation(s):
// \Mux3~5_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux3~4_combout  & (\registerArray[28][28]~q )) # (!\Mux3~4_combout  & ((\registerArray[20][28]~q ))))) # (!\my_rf.rsel1[2]~input_o  & (\Mux3~4_combout ))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux3~4_combout ),
	.datac(\registerArray[28][28]~q ),
	.datad(\registerArray[20][28]~q ),
	.cin(gnd),
	.combout(\Mux3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~5 .lut_mask = 16'hE6C4;
defparam \Mux3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N4
cycloneive_lcell_comb \Mux3~6 (
// Equation(s):
// \Mux3~6_combout  = (\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o ) # ((\Mux3~3_combout )))) # (!\my_rf.rsel1[1]~input_o  & (!\my_rf.rsel1[0]~input_o  & ((\Mux3~5_combout ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux3~3_combout ),
	.datad(\Mux3~5_combout ),
	.cin(gnd),
	.combout(\Mux3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~6 .lut_mask = 16'hB9A8;
defparam \Mux3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N15
dffeas \registerArray[17][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][28] .is_wysiwyg = "true";
defparam \registerArray[17][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N13
dffeas \registerArray[21][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][28] .is_wysiwyg = "true";
defparam \registerArray[21][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N14
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o ) # ((\registerArray[21][28]~q )))) # (!\my_rf.rsel1[2]~input_o  & (!\my_rf.rsel1[3]~input_o  & (\registerArray[17][28]~q )))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[17][28]~q ),
	.datad(\registerArray[21][28]~q ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hBA98;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N20
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// \Mux3~1_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux3~0_combout  & ((\registerArray[29][28]~q ))) # (!\Mux3~0_combout  & (\registerArray[25][28]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux3~0_combout ))))

	.dataa(\registerArray[25][28]~q ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[29][28]~q ),
	.datad(\Mux3~0_combout ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'hF388;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N30
cycloneive_lcell_comb \Mux3~9 (
// Equation(s):
// \Mux3~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux3~6_combout  & (\Mux3~8_combout )) # (!\Mux3~6_combout  & ((\Mux3~1_combout ))))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux3~6_combout ))))

	.dataa(\Mux3~8_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux3~6_combout ),
	.datad(\Mux3~1_combout ),
	.cin(gnd),
	.combout(\Mux3~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~9 .lut_mask = 16'hBCB0;
defparam \Mux3~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N20
cycloneive_lcell_comb \Mux3~15 (
// Equation(s):
// \Mux3~15_combout  = (\Mux3~14_combout ) # ((!\my_rf.rsel1[0]~input_o  & (\registerArray[2][28]~q  & \my_rf.rsel1[1]~input_o )))

	.dataa(\Mux3~14_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[2][28]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux3~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~15 .lut_mask = 16'hBAAA;
defparam \Mux3~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N22
cycloneive_lcell_comb \Mux3~16 (
// Equation(s):
// \Mux3~16_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & (\Mux3~13_combout )) # (!\my_rf.rsel1[2]~input_o  & ((\Mux3~15_combout )))))

	.dataa(\Mux3~13_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux3~15_combout ),
	.cin(gnd),
	.combout(\Mux3~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~16 .lut_mask = 16'hE3E0;
defparam \Mux3~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y31_N31
dffeas \registerArray[11][28] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[28]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][28] .is_wysiwyg = "true";
defparam \registerArray[11][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y31_N30
cycloneive_lcell_comb \Mux3~11 (
// Equation(s):
// \Mux3~11_combout  = (\Mux3~10_combout  & (((\registerArray[11][28]~q )) # (!\my_rf.rsel1[0]~input_o ))) # (!\Mux3~10_combout  & (\my_rf.rsel1[0]~input_o  & ((\registerArray[9][28]~q ))))

	.dataa(\Mux3~10_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[11][28]~q ),
	.datad(\registerArray[9][28]~q ),
	.cin(gnd),
	.combout(\Mux3~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~11 .lut_mask = 16'hE6A2;
defparam \Mux3~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N16
cycloneive_lcell_comb \Mux3~19 (
// Equation(s):
// \Mux3~19_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux3~16_combout  & (\Mux3~18_combout )) # (!\Mux3~16_combout  & ((\Mux3~11_combout ))))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux3~16_combout ))))

	.dataa(\Mux3~18_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\Mux3~16_combout ),
	.datad(\Mux3~11_combout ),
	.cin(gnd),
	.combout(\Mux3~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~19 .lut_mask = 16'hBCB0;
defparam \Mux3~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y38_N2
cycloneive_lcell_comb \Mux3~20 (
// Equation(s):
// \Mux3~20_combout  = (\my_rf.rsel1[4]~input_o  & (\Mux3~9_combout )) # (!\my_rf.rsel1[4]~input_o  & ((\Mux3~19_combout )))

	.dataa(gnd),
	.datab(\my_rf.rsel1[4]~input_o ),
	.datac(\Mux3~9_combout ),
	.datad(\Mux3~19_combout ),
	.cin(gnd),
	.combout(\Mux3~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~20 .lut_mask = 16'hF3C0;
defparam \Mux3~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N30
cycloneive_lcell_comb \Mux2~14 (
// Equation(s):
// \Mux2~14_combout  = (\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\registerArray[3][29]~q )) # (!\my_rf.rsel1[1]~input_o  & ((\registerArray[1][29]~q )))))

	.dataa(\my_rf.rsel1[0]~input_o ),
	.datab(\registerArray[3][29]~q ),
	.datac(\registerArray[1][29]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux2~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~14 .lut_mask = 16'h88A0;
defparam \Mux2~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N18
cycloneive_lcell_comb \Mux2~15 (
// Equation(s):
// \Mux2~15_combout  = (\Mux2~14_combout ) # ((\registerArray[2][29]~q  & (\my_rf.rsel1[1]~input_o  & !\my_rf.rsel1[0]~input_o )))

	.dataa(\registerArray[2][29]~q ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\Mux2~14_combout ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux2~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~15 .lut_mask = 16'hF0F8;
defparam \Mux2~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N28
cycloneive_lcell_comb \Mux2~16 (
// Equation(s):
// \Mux2~16_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux2~13_combout ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((!\my_rf.rsel1[2]~input_o  & \Mux2~15_combout ))))

	.dataa(\Mux2~13_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux2~15_combout ),
	.cin(gnd),
	.combout(\Mux2~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~16 .lut_mask = 16'hCBC8;
defparam \Mux2~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N31
dffeas \registerArray[7][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][29] .is_wysiwyg = "true";
defparam \registerArray[7][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N30
cycloneive_lcell_comb \Mux2~11 (
// Equation(s):
// \Mux2~11_combout  = (\Mux2~10_combout  & (((\registerArray[7][29]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux2~10_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[6][29]~q ))))

	.dataa(\Mux2~10_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[7][29]~q ),
	.datad(\registerArray[6][29]~q ),
	.cin(gnd),
	.combout(\Mux2~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~11 .lut_mask = 16'hE6A2;
defparam \Mux2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N30
cycloneive_lcell_comb \Mux2~19 (
// Equation(s):
// \Mux2~19_combout  = (\Mux2~16_combout  & ((\Mux2~18_combout ) # ((!\my_rf.rsel1[2]~input_o )))) # (!\Mux2~16_combout  & (((\my_rf.rsel1[2]~input_o  & \Mux2~11_combout ))))

	.dataa(\Mux2~18_combout ),
	.datab(\Mux2~16_combout ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux2~11_combout ),
	.cin(gnd),
	.combout(\Mux2~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~19 .lut_mask = 16'hBC8C;
defparam \Mux2~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N9
dffeas \registerArray[25][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][29] .is_wysiwyg = "true";
defparam \registerArray[25][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y33_N9
dffeas \registerArray[17][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][29] .is_wysiwyg = "true";
defparam \registerArray[17][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N8
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// \Mux2~0_combout  = (\my_rf.rsel1[2]~input_o  & (((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o  & (\registerArray[25][29]~q )) # (!\my_rf.rsel1[3]~input_o  & ((\registerArray[17][29]~q )))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[25][29]~q ),
	.datac(\registerArray[17][29]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'hEE50;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y33_N27
dffeas \registerArray[29][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][29] .is_wysiwyg = "true";
defparam \registerArray[29][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X0_Y33_N17
dffeas \registerArray[21][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[29]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][29] .is_wysiwyg = "true";
defparam \registerArray[21][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N26
cycloneive_lcell_comb \Mux2~1 (
// Equation(s):
// \Mux2~1_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux2~0_combout  & (\registerArray[29][29]~q )) # (!\Mux2~0_combout  & ((\registerArray[21][29]~q ))))) # (!\my_rf.rsel1[2]~input_o  & (\Mux2~0_combout ))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\Mux2~0_combout ),
	.datac(\registerArray[29][29]~q ),
	.datad(\registerArray[21][29]~q ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~1 .lut_mask = 16'hE6C4;
defparam \Mux2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y35_N1
dffeas \registerArray[16][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][29] .is_wysiwyg = "true";
defparam \registerArray[16][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y35_N0
cycloneive_lcell_comb \Mux2~4 (
// Equation(s):
// \Mux2~4_combout  = (\my_rf.rsel1[2]~input_o  & ((\registerArray[20][29]~q ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\registerArray[16][29]~q  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\registerArray[20][29]~q ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[16][29]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~4 .lut_mask = 16'hCCB8;
defparam \Mux2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y35_N5
dffeas \registerArray[28][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][29] .is_wysiwyg = "true";
defparam \registerArray[28][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y35_N11
dffeas \registerArray[24][29] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[29]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][29] .is_wysiwyg = "true";
defparam \registerArray[24][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N4
cycloneive_lcell_comb \Mux2~5 (
// Equation(s):
// \Mux2~5_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux2~4_combout  & (\registerArray[28][29]~q )) # (!\Mux2~4_combout  & ((\registerArray[24][29]~q ))))) # (!\my_rf.rsel1[3]~input_o  & (\Mux2~4_combout ))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux2~4_combout ),
	.datac(\registerArray[28][29]~q ),
	.datad(\registerArray[24][29]~q ),
	.cin(gnd),
	.combout(\Mux2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~5 .lut_mask = 16'hE6C4;
defparam \Mux2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N22
cycloneive_lcell_comb \Mux2~6 (
// Equation(s):
// \Mux2~6_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\Mux2~3_combout )) # (!\my_rf.rsel1[1]~input_o  & ((\Mux2~5_combout )))))

	.dataa(\Mux2~3_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux2~5_combout ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~6 .lut_mask = 16'hEE30;
defparam \Mux2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N0
cycloneive_lcell_comb \Mux2~9 (
// Equation(s):
// \Mux2~9_combout  = (\my_rf.rsel1[0]~input_o  & ((\Mux2~6_combout  & (\Mux2~8_combout )) # (!\Mux2~6_combout  & ((\Mux2~1_combout ))))) # (!\my_rf.rsel1[0]~input_o  & (((\Mux2~6_combout ))))

	.dataa(\Mux2~8_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\Mux2~1_combout ),
	.datad(\Mux2~6_combout ),
	.cin(gnd),
	.combout(\Mux2~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~9 .lut_mask = 16'hBBC0;
defparam \Mux2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y33_N24
cycloneive_lcell_comb \Mux2~20 (
// Equation(s):
// \Mux2~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux2~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux2~19_combout ))

	.dataa(\my_rf.rsel1[4]~input_o ),
	.datab(gnd),
	.datac(\Mux2~19_combout ),
	.datad(\Mux2~9_combout ),
	.cin(gnd),
	.combout(\Mux2~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~20 .lut_mask = 16'hFA50;
defparam \Mux2~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N31
dffeas \registerArray[15][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][30] .is_wysiwyg = "true";
defparam \registerArray[15][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N30
cycloneive_lcell_comb \Mux1~18 (
// Equation(s):
// \Mux1~18_combout  = (\Mux1~17_combout  & (((\registerArray[15][30]~q )) # (!\my_rf.rsel1[1]~input_o ))) # (!\Mux1~17_combout  & (\my_rf.rsel1[1]~input_o  & ((\registerArray[14][30]~q ))))

	.dataa(\Mux1~17_combout ),
	.datab(\my_rf.rsel1[1]~input_o ),
	.datac(\registerArray[15][30]~q ),
	.datad(\registerArray[14][30]~q ),
	.cin(gnd),
	.combout(\Mux1~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~18 .lut_mask = 16'hE6A2;
defparam \Mux1~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y31_N3
dffeas \registerArray[6][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][30] .is_wysiwyg = "true";
defparam \registerArray[6][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y31_N29
dffeas \registerArray[7][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][30] .is_wysiwyg = "true";
defparam \registerArray[7][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y31_N28
cycloneive_lcell_comb \Mux1~13 (
// Equation(s):
// \Mux1~13_combout  = (\Mux1~12_combout  & (((\registerArray[7][30]~q ) # (!\my_rf.rsel1[1]~input_o )))) # (!\Mux1~12_combout  & (\registerArray[6][30]~q  & ((\my_rf.rsel1[1]~input_o ))))

	.dataa(\Mux1~12_combout ),
	.datab(\registerArray[6][30]~q ),
	.datac(\registerArray[7][30]~q ),
	.datad(\my_rf.rsel1[1]~input_o ),
	.cin(gnd),
	.combout(\Mux1~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~13 .lut_mask = 16'hE4AA;
defparam \Mux1~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N12
cycloneive_lcell_comb \Mux1~16 (
// Equation(s):
// \Mux1~16_combout  = (\my_rf.rsel1[3]~input_o  & (((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & ((\my_rf.rsel1[2]~input_o  & ((\Mux1~13_combout ))) # (!\my_rf.rsel1[2]~input_o  & (\Mux1~15_combout ))))

	.dataa(\Mux1~15_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux1~13_combout ),
	.cin(gnd),
	.combout(\Mux1~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~16 .lut_mask = 16'hF2C2;
defparam \Mux1~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N30
cycloneive_lcell_comb \Mux1~19 (
// Equation(s):
// \Mux1~19_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux1~16_combout  & ((\Mux1~18_combout ))) # (!\Mux1~16_combout  & (\Mux1~11_combout )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux1~16_combout ))))

	.dataa(\Mux1~11_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\Mux1~18_combout ),
	.datad(\Mux1~16_combout ),
	.cin(gnd),
	.combout(\Mux1~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~19 .lut_mask = 16'hF388;
defparam \Mux1~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N25
dffeas \registerArray[29][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~5_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][30] .is_wysiwyg = "true";
defparam \registerArray[29][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y0_N17
dffeas \registerArray[25][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(\my_rf.wdat[30]~input_o ),
	.asdata(vcc),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][30] .is_wysiwyg = "true";
defparam \registerArray[25][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N24
cycloneive_lcell_comb \Mux1~1 (
// Equation(s):
// \Mux1~1_combout  = (\Mux1~0_combout  & (((\registerArray[29][30]~q )) # (!\my_rf.rsel1[3]~input_o ))) # (!\Mux1~0_combout  & (\my_rf.rsel1[3]~input_o  & ((\registerArray[25][30]~q ))))

	.dataa(\Mux1~0_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[29][30]~q ),
	.datad(\registerArray[25][30]~q ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~1 .lut_mask = 16'hE6A2;
defparam \Mux1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N15
dffeas \registerArray[31][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][30] .is_wysiwyg = "true";
defparam \registerArray[31][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y31_N7
dffeas \registerArray[19][30] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[30]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][30] .is_wysiwyg = "true";
defparam \registerArray[19][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y31_N6
cycloneive_lcell_comb \Mux1~7 (
// Equation(s):
// \Mux1~7_combout  = (\my_rf.rsel1[2]~input_o  & ((\my_rf.rsel1[3]~input_o ) # ((\registerArray[23][30]~q )))) # (!\my_rf.rsel1[2]~input_o  & (!\my_rf.rsel1[3]~input_o  & (\registerArray[19][30]~q )))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[19][30]~q ),
	.datad(\registerArray[23][30]~q ),
	.cin(gnd),
	.combout(\Mux1~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~7 .lut_mask = 16'hBA98;
defparam \Mux1~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N14
cycloneive_lcell_comb \Mux1~8 (
// Equation(s):
// \Mux1~8_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux1~7_combout  & ((\registerArray[31][30]~q ))) # (!\Mux1~7_combout  & (\registerArray[27][30]~q )))) # (!\my_rf.rsel1[3]~input_o  & (((\Mux1~7_combout ))))

	.dataa(\registerArray[27][30]~q ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\registerArray[31][30]~q ),
	.datad(\Mux1~7_combout ),
	.cin(gnd),
	.combout(\Mux1~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~8 .lut_mask = 16'hF388;
defparam \Mux1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N8
cycloneive_lcell_comb \Mux1~9 (
// Equation(s):
// \Mux1~9_combout  = (\Mux1~6_combout  & (((\Mux1~8_combout ) # (!\my_rf.rsel1[0]~input_o )))) # (!\Mux1~6_combout  & (\Mux1~1_combout  & ((\my_rf.rsel1[0]~input_o ))))

	.dataa(\Mux1~6_combout ),
	.datab(\Mux1~1_combout ),
	.datac(\Mux1~8_combout ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux1~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~9 .lut_mask = 16'hE4AA;
defparam \Mux1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N16
cycloneive_lcell_comb \Mux1~20 (
// Equation(s):
// \Mux1~20_combout  = (\my_rf.rsel1[4]~input_o  & ((\Mux1~9_combout ))) # (!\my_rf.rsel1[4]~input_o  & (\Mux1~19_combout ))

	.dataa(\Mux1~19_combout ),
	.datab(\my_rf.rsel1[4]~input_o ),
	.datac(\Mux1~9_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux1~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~20 .lut_mask = 16'hE2E2;
defparam \Mux1~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y35_N17
dffeas \registerArray[20][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][31] .is_wysiwyg = "true";
defparam \registerArray[20][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y35_N19
dffeas \registerArray[16][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][31] .is_wysiwyg = "true";
defparam \registerArray[16][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N18
cycloneive_lcell_comb \Mux0~4 (
// Equation(s):
// \Mux0~4_combout  = (\my_rf.rsel1[2]~input_o  & ((\registerArray[20][31]~q ) # ((\my_rf.rsel1[3]~input_o )))) # (!\my_rf.rsel1[2]~input_o  & (((\registerArray[16][31]~q  & !\my_rf.rsel1[3]~input_o ))))

	.dataa(\my_rf.rsel1[2]~input_o ),
	.datab(\registerArray[20][31]~q ),
	.datac(\registerArray[16][31]~q ),
	.datad(\my_rf.rsel1[3]~input_o ),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~4 .lut_mask = 16'hAAD8;
defparam \Mux0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N11
dffeas \registerArray[28][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][31] .is_wysiwyg = "true";
defparam \registerArray[28][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N25
dffeas \registerArray[24][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][31] .is_wysiwyg = "true";
defparam \registerArray[24][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N10
cycloneive_lcell_comb \Mux0~5 (
// Equation(s):
// \Mux0~5_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux0~4_combout  & (\registerArray[28][31]~q )) # (!\Mux0~4_combout  & ((\registerArray[24][31]~q ))))) # (!\my_rf.rsel1[3]~input_o  & (\Mux0~4_combout ))

	.dataa(\my_rf.rsel1[3]~input_o ),
	.datab(\Mux0~4_combout ),
	.datac(\registerArray[28][31]~q ),
	.datad(\registerArray[24][31]~q ),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~5 .lut_mask = 16'hE6C4;
defparam \Mux0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N24
cycloneive_lcell_comb \Mux0~6 (
// Equation(s):
// \Mux0~6_combout  = (\my_rf.rsel1[0]~input_o  & (((\my_rf.rsel1[1]~input_o )))) # (!\my_rf.rsel1[0]~input_o  & ((\my_rf.rsel1[1]~input_o  & (\Mux0~3_combout )) # (!\my_rf.rsel1[1]~input_o  & ((\Mux0~5_combout )))))

	.dataa(\Mux0~3_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\Mux0~5_combout ),
	.cin(gnd),
	.combout(\Mux0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~6 .lut_mask = 16'hE3E0;
defparam \Mux0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N20
cycloneive_lcell_comb \Mux0~8 (
// Equation(s):
// \Mux0~8_combout  = (\Mux0~7_combout  & (((\registerArray[31][31]~q )) # (!\my_rf.rsel1[2]~input_o ))) # (!\Mux0~7_combout  & (\my_rf.rsel1[2]~input_o  & ((\registerArray[23][31]~q ))))

	.dataa(\Mux0~7_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\registerArray[31][31]~q ),
	.datad(\registerArray[23][31]~q ),
	.cin(gnd),
	.combout(\Mux0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~8 .lut_mask = 16'hE6A2;
defparam \Mux0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N2
cycloneive_lcell_comb \Mux0~9 (
// Equation(s):
// \Mux0~9_combout  = (\Mux0~6_combout  & (((\Mux0~8_combout ) # (!\my_rf.rsel1[0]~input_o )))) # (!\Mux0~6_combout  & (\Mux0~1_combout  & ((\my_rf.rsel1[0]~input_o ))))

	.dataa(\Mux0~1_combout ),
	.datab(\Mux0~6_combout ),
	.datac(\Mux0~8_combout ),
	.datad(\my_rf.rsel1[0]~input_o ),
	.cin(gnd),
	.combout(\Mux0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~9 .lut_mask = 16'hE2CC;
defparam \Mux0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N12
cycloneive_lcell_comb \Mux0~15 (
// Equation(s):
// \Mux0~15_combout  = (\Mux0~14_combout ) # ((!\my_rf.rsel1[0]~input_o  & (\my_rf.rsel1[1]~input_o  & \registerArray[2][31]~q )))

	.dataa(\Mux0~14_combout ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\my_rf.rsel1[1]~input_o ),
	.datad(\registerArray[2][31]~q ),
	.cin(gnd),
	.combout(\Mux0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~15 .lut_mask = 16'hBAAA;
defparam \Mux0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N14
cycloneive_lcell_comb \Mux0~16 (
// Equation(s):
// \Mux0~16_combout  = (\my_rf.rsel1[3]~input_o  & ((\Mux0~13_combout ) # ((\my_rf.rsel1[2]~input_o )))) # (!\my_rf.rsel1[3]~input_o  & (((!\my_rf.rsel1[2]~input_o  & \Mux0~15_combout ))))

	.dataa(\Mux0~13_combout ),
	.datab(\my_rf.rsel1[3]~input_o ),
	.datac(\my_rf.rsel1[2]~input_o ),
	.datad(\Mux0~15_combout ),
	.cin(gnd),
	.combout(\Mux0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~16 .lut_mask = 16'hCBC8;
defparam \Mux0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y37_N23
dffeas \registerArray[4][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][31] .is_wysiwyg = "true";
defparam \registerArray[4][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y37_N13
dffeas \registerArray[5][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][31] .is_wysiwyg = "true";
defparam \registerArray[5][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y37_N22
cycloneive_lcell_comb \Mux0~10 (
// Equation(s):
// \Mux0~10_combout  = (\my_rf.rsel1[1]~input_o  & (\my_rf.rsel1[0]~input_o )) # (!\my_rf.rsel1[1]~input_o  & ((\my_rf.rsel1[0]~input_o  & ((\registerArray[5][31]~q ))) # (!\my_rf.rsel1[0]~input_o  & (\registerArray[4][31]~q ))))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\my_rf.rsel1[0]~input_o ),
	.datac(\registerArray[4][31]~q ),
	.datad(\registerArray[5][31]~q ),
	.cin(gnd),
	.combout(\Mux0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~10 .lut_mask = 16'hDC98;
defparam \Mux0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y37_N21
dffeas \registerArray[7][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][31] .is_wysiwyg = "true";
defparam \registerArray[7][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y37_N11
dffeas \registerArray[6][31] (
	.clk(\clk~inputclkctrl_outclk ),
	.d(gnd),
	.asdata(\my_rf.wdat[31]~input_o ),
	.clrn(\n_rst~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][31] .is_wysiwyg = "true";
defparam \registerArray[6][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y37_N20
cycloneive_lcell_comb \Mux0~11 (
// Equation(s):
// \Mux0~11_combout  = (\my_rf.rsel1[1]~input_o  & ((\Mux0~10_combout  & (\registerArray[7][31]~q )) # (!\Mux0~10_combout  & ((\registerArray[6][31]~q ))))) # (!\my_rf.rsel1[1]~input_o  & (\Mux0~10_combout ))

	.dataa(\my_rf.rsel1[1]~input_o ),
	.datab(\Mux0~10_combout ),
	.datac(\registerArray[7][31]~q ),
	.datad(\registerArray[6][31]~q ),
	.cin(gnd),
	.combout(\Mux0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~11 .lut_mask = 16'hE6C4;
defparam \Mux0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N0
cycloneive_lcell_comb \Mux0~19 (
// Equation(s):
// \Mux0~19_combout  = (\my_rf.rsel1[2]~input_o  & ((\Mux0~16_combout  & (\Mux0~18_combout )) # (!\Mux0~16_combout  & ((\Mux0~11_combout ))))) # (!\my_rf.rsel1[2]~input_o  & (((\Mux0~16_combout ))))

	.dataa(\Mux0~18_combout ),
	.datab(\my_rf.rsel1[2]~input_o ),
	.datac(\Mux0~16_combout ),
	.datad(\Mux0~11_combout ),
	.cin(gnd),
	.combout(\Mux0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~19 .lut_mask = 16'hBCB0;
defparam \Mux0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y38_N10
cycloneive_lcell_comb \Mux0~20 (
// Equation(s):
// \Mux0~20_combout  = (\my_rf.rsel1[4]~input_o  & (\Mux0~9_combout )) # (!\my_rf.rsel1[4]~input_o  & ((\Mux0~19_combout )))

	.dataa(gnd),
	.datab(\Mux0~9_combout ),
	.datac(\my_rf.rsel1[4]~input_o ),
	.datad(\Mux0~19_combout ),
	.cin(gnd),
	.combout(\Mux0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~20 .lut_mask = 16'hCFC0;
defparam \Mux0~20 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule
