// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 64-Bit"
// VERSION "Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"

// DATE "10/04/2017 17:56:17"

// 
// Device: Altera EP4CE115F29C8 Package FBGA780
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module system (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	CLK,
	nRST,
	\syif.halt ,
	\syif.load ,
	\syif.addr ,
	\syif.store ,
	\syif.REN ,
	\syif.WEN ,
	\syif.tbCTRL );
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	CLK;
input 	nRST;
output 	\syif.halt ;
output 	[31:0] \syif.load ;
input 	[31:0] \syif.addr ;
input 	[31:0] \syif.store ;
input 	\syif.REN ;
input 	\syif.WEN ;
input 	\syif.tbCTRL ;

// Design Ports Information
// syif.halt	=>  Location: PIN_AD12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[0]	=>  Location: PIN_AC15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[1]	=>  Location: PIN_AC14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[2]	=>  Location: PIN_J15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[3]	=>  Location: PIN_AH17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[4]	=>  Location: PIN_AB10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[5]	=>  Location: PIN_AE16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[6]	=>  Location: PIN_Y14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[7]	=>  Location: PIN_C15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[8]	=>  Location: PIN_R25,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[9]	=>  Location: PIN_V1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[10]	=>  Location: PIN_J16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[11]	=>  Location: PIN_AG17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[12]	=>  Location: PIN_AE17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[13]	=>  Location: PIN_U27,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[14]	=>  Location: PIN_AD15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[15]	=>  Location: PIN_B17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[16]	=>  Location: PIN_F15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[17]	=>  Location: PIN_AG19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[18]	=>  Location: PIN_AF15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[19]	=>  Location: PIN_C12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[20]	=>  Location: PIN_AH19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[21]	=>  Location: PIN_H16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[22]	=>  Location: PIN_D16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[23]	=>  Location: PIN_H15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[24]	=>  Location: PIN_AF16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[25]	=>  Location: PIN_AA16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[26]	=>  Location: PIN_AA15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[27]	=>  Location: PIN_V2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[28]	=>  Location: PIN_AE15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[29]	=>  Location: PIN_C16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[30]	=>  Location: PIN_A17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[31]	=>  Location: PIN_A10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// nRST	=>  Location: PIN_Y2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.tbCTRL	=>  Location: PIN_AG15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[1]	=>  Location: PIN_AH15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[0]	=>  Location: PIN_AG12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[3]	=>  Location: PIN_AB15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[2]	=>  Location: PIN_Y15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[5]	=>  Location: PIN_AF13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[4]	=>  Location: PIN_AB14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[7]	=>  Location: PIN_D15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[6]	=>  Location: PIN_V3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[9]	=>  Location: PIN_D14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[8]	=>  Location: PIN_H14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[11]	=>  Location: PIN_A11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[10]	=>  Location: PIN_AF11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[13]	=>  Location: PIN_T26,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[12]	=>  Location: PIN_AF14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[15]	=>  Location: PIN_J14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[14]	=>  Location: PIN_T3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[17]	=>  Location: PIN_AE11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[16]	=>  Location: PIN_AE13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[19]	=>  Location: PIN_H17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[18]	=>  Location: PIN_G14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[21]	=>  Location: PIN_E17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[20]	=>  Location: PIN_AE12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[23]	=>  Location: PIN_B11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[22]	=>  Location: PIN_D13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[25]	=>  Location: PIN_J12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[24]	=>  Location: PIN_AC12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[27]	=>  Location: PIN_AC11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[26]	=>  Location: PIN_AH11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[29]	=>  Location: PIN_AD11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[28]	=>  Location: PIN_AH12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[31]	=>  Location: PIN_D12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[30]	=>  Location: PIN_AD17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.WEN	=>  Location: PIN_AD14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.REN	=>  Location: PIN_U24,	 I/O Standard: 2.5 V,	 Current Strength: Default
// CLK	=>  Location: PIN_J1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[0]	=>  Location: PIN_C14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[1]	=>  Location: PIN_F14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[2]	=>  Location: PIN_Y22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[3]	=>  Location: PIN_R5,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[4]	=>  Location: PIN_Y12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[5]	=>  Location: PIN_AB12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[6]	=>  Location: PIN_C13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[7]	=>  Location: PIN_AC10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[8]	=>  Location: PIN_AE14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[9]	=>  Location: PIN_J13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[10]	=>  Location: PIN_AB16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[11]	=>  Location: PIN_AG11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[12]	=>  Location: PIN_G15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[13]	=>  Location: PIN_AG18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[14]	=>  Location: PIN_AB13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[15]	=>  Location: PIN_V4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[16]	=>  Location: PIN_AA12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[17]	=>  Location: PIN_R1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[18]	=>  Location: PIN_Y13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[19]	=>  Location: PIN_AH18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[20]	=>  Location: PIN_G13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[21]	=>  Location: PIN_E15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[22]	=>  Location: PIN_R23,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[23]	=>  Location: PIN_W22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[24]	=>  Location: PIN_AF17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[25]	=>  Location: PIN_AA13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[26]	=>  Location: PIN_A12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[27]	=>  Location: PIN_AF10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[28]	=>  Location: PIN_R2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[29]	=>  Location: PIN_E14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[30]	=>  Location: PIN_F17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[31]	=>  Location: PIN_AA14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tms	=>  Location: PIN_P8,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tck	=>  Location: PIN_P5,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdi	=>  Location: PIN_P7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdo	=>  Location: PIN_P6,	 I/O Standard: 2.5 V,	 Current Strength: Default


wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ;
wire \RAM|ramif.ramload[0]~0_combout ;
wire \CPU|DP|EXMEM|exmem_if.dWEN_o~q ;
wire \CPU|DP|EXMEM|exmem_if.dREN_o~q ;
wire \ramaddr~0_combout ;
wire \ramaddr~1_combout ;
wire \ramaddr~2_combout ;
wire \ramaddr~3_combout ;
wire \ramaddr~4_combout ;
wire \ramaddr~5_combout ;
wire \ramaddr~6_combout ;
wire \ramaddr~7_combout ;
wire \ramaddr~8_combout ;
wire \ramaddr~9_combout ;
wire \ramaddr~10_combout ;
wire \ramaddr~11_combout ;
wire \ramaddr~12_combout ;
wire \ramaddr~13_combout ;
wire \ramaddr~14_combout ;
wire \ramaddr~15_combout ;
wire \ramaddr~16_combout ;
wire \ramaddr~17_combout ;
wire \ramaddr~18_combout ;
wire \ramaddr~19_combout ;
wire \ramaddr~20_combout ;
wire \ramaddr~21_combout ;
wire \ramaddr~22_combout ;
wire \ramaddr~23_combout ;
wire \ramaddr~24_combout ;
wire \ramaddr~25_combout ;
wire \ramaddr~26_combout ;
wire \ramaddr~27_combout ;
wire \ramaddr~28_combout ;
wire \ramaddr~29_combout ;
wire \ramaddr~30_combout ;
wire \ramaddr~31_combout ;
wire \ramaddr~32_combout ;
wire \ramaddr~33_combout ;
wire \ramaddr~34_combout ;
wire \ramaddr~35_combout ;
wire \ramaddr~36_combout ;
wire \ramaddr~37_combout ;
wire \ramaddr~38_combout ;
wire \ramaddr~39_combout ;
wire \ramaddr~40_combout ;
wire \ramaddr~41_combout ;
wire \ramaddr~42_combout ;
wire \ramaddr~43_combout ;
wire \ramaddr~44_combout ;
wire \ramaddr~45_combout ;
wire \ramaddr~46_combout ;
wire \ramaddr~47_combout ;
wire \ramaddr~48_combout ;
wire \ramaddr~49_combout ;
wire \ramaddr~50_combout ;
wire \ramaddr~51_combout ;
wire \ramaddr~52_combout ;
wire \ramaddr~53_combout ;
wire \ramaddr~54_combout ;
wire \ramaddr~55_combout ;
wire \ramaddr~56_combout ;
wire \ramaddr~57_combout ;
wire \ramaddr~58_combout ;
wire \ramaddr~59_combout ;
wire \ramaddr~60_combout ;
wire \ramaddr~61_combout ;
wire \ramaddr~62_combout ;
wire \ramaddr~63_combout ;
wire \RAM|ramif.ramload[0]~2_combout ;
wire \RAM|ramif.ramload[1]~3_combout ;
wire \RAM|ramif.ramload[1]~5_combout ;
wire \RAM|always1~0_combout ;
wire \RAM|always1~1_combout ;
wire \RAM|ramif.ramload[2]~6_combout ;
wire \RAM|ramif.ramload[3]~7_combout ;
wire \RAM|ramif.ramload[4]~8_combout ;
wire \RAM|ramif.ramload[5]~9_combout ;
wire \RAM|ramif.ramload[6]~10_combout ;
wire \RAM|ramif.ramload[7]~11_combout ;
wire \RAM|ramif.ramload[8]~12_combout ;
wire \RAM|ramif.ramload[9]~13_combout ;
wire \RAM|ramif.ramload[10]~14_combout ;
wire \RAM|ramif.ramload[11]~15_combout ;
wire \RAM|ramif.ramload[12]~16_combout ;
wire \RAM|ramif.ramload[13]~17_combout ;
wire \RAM|ramif.ramload[14]~18_combout ;
wire \RAM|ramif.ramload[15]~19_combout ;
wire \RAM|ramif.ramload[16]~20_combout ;
wire \RAM|ramif.ramload[17]~21_combout ;
wire \RAM|ramif.ramload[18]~22_combout ;
wire \RAM|ramif.ramload[19]~23_combout ;
wire \RAM|ramif.ramload[20]~24_combout ;
wire \RAM|ramif.ramload[21]~25_combout ;
wire \RAM|ramif.ramload[22]~26_combout ;
wire \RAM|ramif.ramload[23]~27_combout ;
wire \RAM|ramif.ramload[24]~28_combout ;
wire \RAM|ramif.ramload[25]~29_combout ;
wire \RAM|ramif.ramload[26]~30_combout ;
wire \RAM|ramif.ramload[27]~31_combout ;
wire \RAM|ramif.ramload[28]~32_combout ;
wire \RAM|ramif.ramload[29]~33_combout ;
wire \RAM|ramif.ramload[30]~34_combout ;
wire \RAM|ramif.ramload[31]~35_combout ;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ;
wire \CPUCLK~q ;
wire \ramWEN~0_combout ;
wire \ramstore~0_combout ;
wire \ramREN~0_combout ;
wire \RAM|ramstate~0_combout ;
wire \ramstore~1_combout ;
wire \ramstore~2_combout ;
wire \ramstore~3_combout ;
wire \ramstore~4_combout ;
wire \ramstore~5_combout ;
wire \ramstore~6_combout ;
wire \ramstore~7_combout ;
wire \ramstore~8_combout ;
wire \ramstore~9_combout ;
wire \ramstore~10_combout ;
wire \ramstore~11_combout ;
wire \ramstore~12_combout ;
wire \ramstore~13_combout ;
wire \ramstore~14_combout ;
wire \ramstore~15_combout ;
wire \ramstore~16_combout ;
wire \ramstore~17_combout ;
wire \ramstore~18_combout ;
wire \ramstore~19_combout ;
wire \ramstore~20_combout ;
wire \ramstore~21_combout ;
wire \ramstore~22_combout ;
wire \ramstore~23_combout ;
wire \ramstore~24_combout ;
wire \ramstore~25_combout ;
wire \ramstore~26_combout ;
wire \ramstore~27_combout ;
wire \ramstore~28_combout ;
wire \ramstore~29_combout ;
wire \ramstore~30_combout ;
wire \ramstore~31_combout ;
wire \Equal0~0_combout ;
wire \CPUCLK~0_combout ;
wire \count[3]~0_combout ;
wire \count[2]~1_combout ;
wire \count[1]~2_combout ;
wire \count~3_combout ;
wire \ramaddr~29_wirecell_combout ;
wire \altera_internal_jtag~TCKUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ;
wire \nRST~input_o ;
wire \syif.tbCTRL~input_o ;
wire \syif.addr[1]~input_o ;
wire \syif.addr[0]~input_o ;
wire \syif.addr[3]~input_o ;
wire \syif.addr[2]~input_o ;
wire \syif.addr[5]~input_o ;
wire \syif.addr[4]~input_o ;
wire \syif.addr[7]~input_o ;
wire \syif.addr[6]~input_o ;
wire \syif.addr[9]~input_o ;
wire \syif.addr[8]~input_o ;
wire \syif.addr[11]~input_o ;
wire \syif.addr[10]~input_o ;
wire \syif.addr[13]~input_o ;
wire \syif.addr[12]~input_o ;
wire \syif.addr[15]~input_o ;
wire \syif.addr[14]~input_o ;
wire \syif.addr[17]~input_o ;
wire \syif.addr[16]~input_o ;
wire \syif.addr[19]~input_o ;
wire \syif.addr[18]~input_o ;
wire \syif.addr[21]~input_o ;
wire \syif.addr[20]~input_o ;
wire \syif.addr[23]~input_o ;
wire \syif.addr[22]~input_o ;
wire \syif.addr[25]~input_o ;
wire \syif.addr[24]~input_o ;
wire \syif.addr[27]~input_o ;
wire \syif.addr[26]~input_o ;
wire \syif.addr[29]~input_o ;
wire \syif.addr[28]~input_o ;
wire \syif.addr[31]~input_o ;
wire \syif.addr[30]~input_o ;
wire \syif.WEN~input_o ;
wire \syif.REN~input_o ;
wire \CLK~input_o ;
wire \syif.store[0]~input_o ;
wire \syif.store[1]~input_o ;
wire \syif.store[2]~input_o ;
wire \syif.store[3]~input_o ;
wire \syif.store[4]~input_o ;
wire \syif.store[5]~input_o ;
wire \syif.store[6]~input_o ;
wire \syif.store[7]~input_o ;
wire \syif.store[8]~input_o ;
wire \syif.store[9]~input_o ;
wire \syif.store[10]~input_o ;
wire \syif.store[11]~input_o ;
wire \syif.store[12]~input_o ;
wire \syif.store[13]~input_o ;
wire \syif.store[14]~input_o ;
wire \syif.store[15]~input_o ;
wire \syif.store[16]~input_o ;
wire \syif.store[17]~input_o ;
wire \syif.store[18]~input_o ;
wire \syif.store[19]~input_o ;
wire \syif.store[20]~input_o ;
wire \syif.store[21]~input_o ;
wire \syif.store[22]~input_o ;
wire \syif.store[23]~input_o ;
wire \syif.store[24]~input_o ;
wire \syif.store[25]~input_o ;
wire \syif.store[26]~input_o ;
wire \syif.store[27]~input_o ;
wire \syif.store[28]~input_o ;
wire \syif.store[29]~input_o ;
wire \syif.store[30]~input_o ;
wire \syif.store[31]~input_o ;
wire \altera_internal_jtag~TCKUTAPclkctrl_outclk ;
wire \CPUCLK~clkctrl_outclk ;
wire \nRST~inputclkctrl_outclk ;
wire \CLK~inputclkctrl_outclk ;
wire \CPU|DP|dpif.halt~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TDIUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ;
wire \~QIC_CREATED_GND~I_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~8 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~10 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~14 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~16 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ;
wire \altera_internal_jtag~TDO ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg ;
wire [9:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg ;
wire [5:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt ;
wire [15:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR ;
wire [3:0] count;
wire [31:0] \CPU|DP|pc ;
wire [31:0] \CPU|DP|EXMEM|exmem_if.rdat2_o ;
wire [31:0] \CPU|DP|EXMEM|exmem_if.out_o ;
wire [3:0] \RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg ;


pipeline CPU(
	.ramiframload_0(\RAM|ramif.ramload[0]~0_combout ),
	.exmem_ifout_o_1(\CPU|DP|EXMEM|exmem_if.out_o [1]),
	.exmem_ifdWEN_o(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.exmem_ifdREN_o(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.pc_1(\CPU|DP|pc [1]),
	.exmem_ifout_o_0(\CPU|DP|EXMEM|exmem_if.out_o [0]),
	.pc_0(\CPU|DP|pc [0]),
	.exmem_ifout_o_3(\CPU|DP|EXMEM|exmem_if.out_o [3]),
	.pc_3(\CPU|DP|pc [3]),
	.exmem_ifout_o_2(\CPU|DP|EXMEM|exmem_if.out_o [2]),
	.pc_2(\CPU|DP|pc [2]),
	.exmem_ifout_o_5(\CPU|DP|EXMEM|exmem_if.out_o [5]),
	.pc_5(\CPU|DP|pc [5]),
	.pc_4(\CPU|DP|pc [4]),
	.exmem_ifout_o_4(\CPU|DP|EXMEM|exmem_if.out_o [4]),
	.exmem_ifout_o_7(\CPU|DP|EXMEM|exmem_if.out_o [7]),
	.pc_7(\CPU|DP|pc [7]),
	.exmem_ifout_o_6(\CPU|DP|EXMEM|exmem_if.out_o [6]),
	.pc_6(\CPU|DP|pc [6]),
	.exmem_ifout_o_9(\CPU|DP|EXMEM|exmem_if.out_o [9]),
	.pc_9(\CPU|DP|pc [9]),
	.pc_8(\CPU|DP|pc [8]),
	.exmem_ifout_o_8(\CPU|DP|EXMEM|exmem_if.out_o [8]),
	.exmem_ifout_o_11(\CPU|DP|EXMEM|exmem_if.out_o [11]),
	.pc_11(\CPU|DP|pc [11]),
	.exmem_ifout_o_10(\CPU|DP|EXMEM|exmem_if.out_o [10]),
	.pc_10(\CPU|DP|pc [10]),
	.pc_13(\CPU|DP|pc [13]),
	.exmem_ifout_o_13(\CPU|DP|EXMEM|exmem_if.out_o [13]),
	.pc_12(\CPU|DP|pc [12]),
	.exmem_ifout_o_12(\CPU|DP|EXMEM|exmem_if.out_o [12]),
	.exmem_ifout_o_15(\CPU|DP|EXMEM|exmem_if.out_o [15]),
	.pc_15(\CPU|DP|pc [15]),
	.pc_14(\CPU|DP|pc [14]),
	.exmem_ifout_o_14(\CPU|DP|EXMEM|exmem_if.out_o [14]),
	.pc_17(\CPU|DP|pc [17]),
	.exmem_ifout_o_17(\CPU|DP|EXMEM|exmem_if.out_o [17]),
	.exmem_ifout_o_16(\CPU|DP|EXMEM|exmem_if.out_o [16]),
	.pc_16(\CPU|DP|pc [16]),
	.exmem_ifout_o_19(\CPU|DP|EXMEM|exmem_if.out_o [19]),
	.pc_19(\CPU|DP|pc [19]),
	.exmem_ifout_o_18(\CPU|DP|EXMEM|exmem_if.out_o [18]),
	.pc_18(\CPU|DP|pc [18]),
	.pc_21(\CPU|DP|pc [21]),
	.exmem_ifout_o_21(\CPU|DP|EXMEM|exmem_if.out_o [21]),
	.pc_20(\CPU|DP|pc [20]),
	.exmem_ifout_o_20(\CPU|DP|EXMEM|exmem_if.out_o [20]),
	.exmem_ifout_o_23(\CPU|DP|EXMEM|exmem_if.out_o [23]),
	.pc_23(\CPU|DP|pc [23]),
	.exmem_ifout_o_22(\CPU|DP|EXMEM|exmem_if.out_o [22]),
	.pc_22(\CPU|DP|pc [22]),
	.pc_25(\CPU|DP|pc [25]),
	.exmem_ifout_o_25(\CPU|DP|EXMEM|exmem_if.out_o [25]),
	.pc_24(\CPU|DP|pc [24]),
	.exmem_ifout_o_24(\CPU|DP|EXMEM|exmem_if.out_o [24]),
	.exmem_ifout_o_27(\CPU|DP|EXMEM|exmem_if.out_o [27]),
	.pc_27(\CPU|DP|pc [27]),
	.exmem_ifout_o_26(\CPU|DP|EXMEM|exmem_if.out_o [26]),
	.pc_26(\CPU|DP|pc [26]),
	.pc_29(\CPU|DP|pc [29]),
	.exmem_ifout_o_29(\CPU|DP|EXMEM|exmem_if.out_o [29]),
	.exmem_ifout_o_28(\CPU|DP|EXMEM|exmem_if.out_o [28]),
	.pc_28(\CPU|DP|pc [28]),
	.exmem_ifout_o_31(\CPU|DP|EXMEM|exmem_if.out_o [31]),
	.pc_31(\CPU|DP|pc [31]),
	.exmem_ifout_o_30(\CPU|DP|EXMEM|exmem_if.out_o [30]),
	.pc_30(\CPU|DP|pc [30]),
	.ramiframload_01(\RAM|ramif.ramload[0]~2_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~3_combout ),
	.ramiframload_11(\RAM|ramif.ramload[1]~5_combout ),
	.always1(\RAM|always1~0_combout ),
	.always11(\RAM|always1~1_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~6_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~7_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~8_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~9_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~10_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~11_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~12_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~13_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~14_combout ),
	.ramiframload_111(\RAM|ramif.ramload[11]~15_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~16_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~17_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~18_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~19_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~20_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~21_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~22_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~23_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~24_combout ),
	.ramiframload_21(\RAM|ramif.ramload[21]~25_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~26_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~27_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~28_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~29_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~30_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~31_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~32_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~33_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~34_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~35_combout ),
	.exmem_ifrdat2_o_0(\CPU|DP|EXMEM|exmem_if.rdat2_o [0]),
	.ramstate(\RAM|ramstate~0_combout ),
	.exmem_ifrdat2_o_1(\CPU|DP|EXMEM|exmem_if.rdat2_o [1]),
	.exmem_ifrdat2_o_2(\CPU|DP|EXMEM|exmem_if.rdat2_o [2]),
	.exmem_ifrdat2_o_3(\CPU|DP|EXMEM|exmem_if.rdat2_o [3]),
	.exmem_ifrdat2_o_4(\CPU|DP|EXMEM|exmem_if.rdat2_o [4]),
	.exmem_ifrdat2_o_5(\CPU|DP|EXMEM|exmem_if.rdat2_o [5]),
	.exmem_ifrdat2_o_6(\CPU|DP|EXMEM|exmem_if.rdat2_o [6]),
	.exmem_ifrdat2_o_7(\CPU|DP|EXMEM|exmem_if.rdat2_o [7]),
	.exmem_ifrdat2_o_8(\CPU|DP|EXMEM|exmem_if.rdat2_o [8]),
	.exmem_ifrdat2_o_9(\CPU|DP|EXMEM|exmem_if.rdat2_o [9]),
	.exmem_ifrdat2_o_10(\CPU|DP|EXMEM|exmem_if.rdat2_o [10]),
	.exmem_ifrdat2_o_11(\CPU|DP|EXMEM|exmem_if.rdat2_o [11]),
	.exmem_ifrdat2_o_12(\CPU|DP|EXMEM|exmem_if.rdat2_o [12]),
	.exmem_ifrdat2_o_13(\CPU|DP|EXMEM|exmem_if.rdat2_o [13]),
	.exmem_ifrdat2_o_14(\CPU|DP|EXMEM|exmem_if.rdat2_o [14]),
	.exmem_ifrdat2_o_15(\CPU|DP|EXMEM|exmem_if.rdat2_o [15]),
	.exmem_ifrdat2_o_16(\CPU|DP|EXMEM|exmem_if.rdat2_o [16]),
	.exmem_ifrdat2_o_17(\CPU|DP|EXMEM|exmem_if.rdat2_o [17]),
	.exmem_ifrdat2_o_18(\CPU|DP|EXMEM|exmem_if.rdat2_o [18]),
	.exmem_ifrdat2_o_19(\CPU|DP|EXMEM|exmem_if.rdat2_o [19]),
	.exmem_ifrdat2_o_20(\CPU|DP|EXMEM|exmem_if.rdat2_o [20]),
	.exmem_ifrdat2_o_21(\CPU|DP|EXMEM|exmem_if.rdat2_o [21]),
	.exmem_ifrdat2_o_22(\CPU|DP|EXMEM|exmem_if.rdat2_o [22]),
	.exmem_ifrdat2_o_23(\CPU|DP|EXMEM|exmem_if.rdat2_o [23]),
	.exmem_ifrdat2_o_24(\CPU|DP|EXMEM|exmem_if.rdat2_o [24]),
	.exmem_ifrdat2_o_25(\CPU|DP|EXMEM|exmem_if.rdat2_o [25]),
	.exmem_ifrdat2_o_26(\CPU|DP|EXMEM|exmem_if.rdat2_o [26]),
	.exmem_ifrdat2_o_27(\CPU|DP|EXMEM|exmem_if.rdat2_o [27]),
	.exmem_ifrdat2_o_28(\CPU|DP|EXMEM|exmem_if.rdat2_o [28]),
	.exmem_ifrdat2_o_29(\CPU|DP|EXMEM|exmem_if.rdat2_o [29]),
	.exmem_ifrdat2_o_30(\CPU|DP|EXMEM|exmem_if.rdat2_o [30]),
	.exmem_ifrdat2_o_31(\CPU|DP|EXMEM|exmem_if.rdat2_o [31]),
	.CLK(\CPUCLK~clkctrl_outclk ),
	.nRST(\nRST~inputclkctrl_outclk ),
	.dpifhalt(\CPU|DP|dpif.halt~q ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

ram RAM(
	.is_in_use_reg(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.ramiframload_0(\RAM|ramif.ramload[0]~0_combout ),
	.ramaddr(\ramaddr~1_combout ),
	.ramaddr1(\ramaddr~3_combout ),
	.ramaddr2(\ramaddr~5_combout ),
	.ramaddr3(\ramaddr~7_combout ),
	.ramaddr4(\ramaddr~9_combout ),
	.ramaddr5(\ramaddr~11_combout ),
	.ramaddr6(\ramaddr~13_combout ),
	.ramaddr7(\ramaddr~15_combout ),
	.ramaddr8(\ramaddr~17_combout ),
	.ramaddr9(\ramaddr~19_combout ),
	.ramaddr10(\ramaddr~21_combout ),
	.ramaddr11(\ramaddr~23_combout ),
	.ramaddr12(\ramaddr~25_combout ),
	.ramaddr13(\ramaddr~27_combout ),
	.ramaddr14(\ramaddr~29_combout ),
	.ramaddr15(\ramaddr~31_combout ),
	.\ramif.ramaddr ({gnd,gnd,\ramaddr~57_combout ,gnd,\ramaddr~53_combout ,gnd,\ramaddr~49_combout ,gnd,\ramaddr~45_combout ,gnd,gnd,gnd,gnd,gnd,\ramaddr~33_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.ramaddr16(\ramaddr~35_combout ),
	.ramaddr17(\ramaddr~37_combout ),
	.ramaddr18(\ramaddr~39_combout ),
	.ramaddr19(\ramaddr~41_combout ),
	.ramaddr20(\ramaddr~43_combout ),
	.ramaddr21(\ramaddr~47_combout ),
	.ramaddr22(\ramaddr~51_combout ),
	.ramaddr23(\ramaddr~55_combout ),
	.ramaddr24(\ramaddr~59_combout ),
	.ramaddr25(\ramaddr~61_combout ),
	.ramaddr26(\ramaddr~63_combout ),
	.ramiframload_01(\RAM|ramif.ramload[0]~2_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~3_combout ),
	.ramiframload_11(\RAM|ramif.ramload[1]~5_combout ),
	.always1(\RAM|always1~0_combout ),
	.always11(\RAM|always1~1_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~6_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~7_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~8_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~9_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~10_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~11_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~12_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~13_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~14_combout ),
	.ramiframload_111(\RAM|ramif.ramload[11]~15_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~16_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~17_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~18_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~19_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~20_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~21_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~22_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~23_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~24_combout ),
	.ramiframload_21(\RAM|ramif.ramload[21]~25_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~26_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~27_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~28_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~29_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~30_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~31_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~32_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~33_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~34_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~35_combout ),
	.ir_loaded_address_reg_0(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.ir_loaded_address_reg_1(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.ir_loaded_address_reg_2(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.ir_loaded_address_reg_3(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.tdo(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.ramWEN(\ramWEN~0_combout ),
	.ramstore(\ramstore~0_combout ),
	.ramREN(\ramREN~0_combout ),
	.ramstate(\RAM|ramstate~0_combout ),
	.ramstore1(\ramstore~1_combout ),
	.ramstore2(\ramstore~2_combout ),
	.ramstore3(\ramstore~3_combout ),
	.ramstore4(\ramstore~4_combout ),
	.ramstore5(\ramstore~5_combout ),
	.ramstore6(\ramstore~6_combout ),
	.ramstore7(\ramstore~7_combout ),
	.ramstore8(\ramstore~8_combout ),
	.ramstore9(\ramstore~9_combout ),
	.ramstore10(\ramstore~10_combout ),
	.ramstore11(\ramstore~11_combout ),
	.ramstore12(\ramstore~12_combout ),
	.ramstore13(\ramstore~13_combout ),
	.ramstore14(\ramstore~14_combout ),
	.ramstore15(\ramstore~15_combout ),
	.ramstore16(\ramstore~16_combout ),
	.ramstore17(\ramstore~17_combout ),
	.ramstore18(\ramstore~18_combout ),
	.ramstore19(\ramstore~19_combout ),
	.ramstore20(\ramstore~20_combout ),
	.ramstore21(\ramstore~21_combout ),
	.ramstore22(\ramstore~22_combout ),
	.ramstore23(\ramstore~23_combout ),
	.ramstore24(\ramstore~24_combout ),
	.ramstore25(\ramstore~25_combout ),
	.ramstore26(\ramstore~26_combout ),
	.ramstore27(\ramstore~27_combout ),
	.ramstore28(\ramstore~28_combout ),
	.ramstore29(\ramstore~29_combout ),
	.ramstore30(\ramstore~30_combout ),
	.ramstore31(\ramstore~31_combout ),
	.ramaddr27(\ramaddr~29_wirecell_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.irf_reg_0_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.irf_reg_1_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.irf_reg_2_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.irf_reg_3_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.irf_reg_4_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.node_ena_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.clr_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.virtual_ir_scan_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.state_5(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.state_8(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.nRST(\nRST~input_o ),
	.syiftbCTRL(\syif.tbCTRL~input_o ),
	.syifWEN(\syif.WEN~input_o ),
	.syifREN(\syif.REN~input_o ),
	.altera_internal_jtag1(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.nRST1(\nRST~inputclkctrl_outclk ),
	.CLK(\CLK~inputclkctrl_outclk ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X54_Y33_N10
cycloneive_lcell_comb \ramaddr~0 (
// Equation(s):
// \ramaddr~0_combout  = (exmem_ifdWEN_o & (exmem_ifout_o_1)) # (!exmem_ifdWEN_o & ((exmem_ifdREN_o & (exmem_ifout_o_1)) # (!exmem_ifdREN_o & ((pc_1)))))

	.dataa(\CPU|DP|EXMEM|exmem_if.out_o [1]),
	.datab(\CPU|DP|pc [1]),
	.datac(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~0 .lut_mask = 16'hAAAC;
defparam \ramaddr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N24
cycloneive_lcell_comb \ramaddr~1 (
// Equation(s):
// \ramaddr~1_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[1]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~0_combout )))

	.dataa(\syif.addr[1]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~0_combout ),
	.cin(gnd),
	.combout(\ramaddr~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~1 .lut_mask = 16'hBB88;
defparam \ramaddr~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N30
cycloneive_lcell_comb \ramaddr~2 (
// Equation(s):
// \ramaddr~2_combout  = (exmem_ifdREN_o & (exmem_ifout_o_0)) # (!exmem_ifdREN_o & ((exmem_ifdWEN_o & (exmem_ifout_o_0)) # (!exmem_ifdWEN_o & ((pc_0)))))

	.dataa(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datab(\CPU|DP|EXMEM|exmem_if.out_o [0]),
	.datac(\CPU|DP|pc [0]),
	.datad(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~2 .lut_mask = 16'hCCD8;
defparam \ramaddr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N16
cycloneive_lcell_comb \ramaddr~3 (
// Equation(s):
// \ramaddr~3_combout  = (\syif.tbCTRL~input_o  & ((\syif.addr[0]~input_o ))) # (!\syif.tbCTRL~input_o  & (\ramaddr~2_combout ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramaddr~2_combout ),
	.datad(\syif.addr[0]~input_o ),
	.cin(gnd),
	.combout(\ramaddr~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~3 .lut_mask = 16'hFC30;
defparam \ramaddr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N22
cycloneive_lcell_comb \ramaddr~4 (
// Equation(s):
// \ramaddr~4_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[3]~input_o )) # (!\syif.tbCTRL~input_o  & (((exmem_ifdREN_o) # (exmem_ifdWEN_o))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[3]~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~4 .lut_mask = 16'hDDD8;
defparam \ramaddr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N24
cycloneive_lcell_comb \ramaddr~5 (
// Equation(s):
// \ramaddr~5_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~4_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~4_combout  & ((exmem_ifout_o_3))) # (!\ramaddr~4_combout  & (pc_3))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|pc [3]),
	.datac(\ramaddr~4_combout ),
	.datad(\CPU|DP|EXMEM|exmem_if.out_o [3]),
	.cin(gnd),
	.combout(\ramaddr~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~5 .lut_mask = 16'hF4A4;
defparam \ramaddr~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N28
cycloneive_lcell_comb \ramaddr~6 (
// Equation(s):
// \ramaddr~6_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[2]~input_o )) # (!\syif.tbCTRL~input_o  & (((exmem_ifdREN_o) # (exmem_ifdWEN_o))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[2]~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~6 .lut_mask = 16'hDDD8;
defparam \ramaddr~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N10
cycloneive_lcell_comb \ramaddr~7 (
// Equation(s):
// \ramaddr~7_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~6_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~6_combout  & (exmem_ifout_o_2)) # (!\ramaddr~6_combout  & ((pc_2)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|EXMEM|exmem_if.out_o [2]),
	.datac(\CPU|DP|pc [2]),
	.datad(\ramaddr~6_combout ),
	.cin(gnd),
	.combout(\ramaddr~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~7 .lut_mask = 16'hEE50;
defparam \ramaddr~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N10
cycloneive_lcell_comb \ramaddr~8 (
// Equation(s):
// \ramaddr~8_combout  = (exmem_ifdWEN_o & (((exmem_ifout_o_5)))) # (!exmem_ifdWEN_o & ((exmem_ifdREN_o & ((exmem_ifout_o_5))) # (!exmem_ifdREN_o & (pc_5))))

	.dataa(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datab(\CPU|DP|pc [5]),
	.datac(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.out_o [5]),
	.cin(gnd),
	.combout(\ramaddr~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~8 .lut_mask = 16'hFE04;
defparam \ramaddr~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N28
cycloneive_lcell_comb \ramaddr~9 (
// Equation(s):
// \ramaddr~9_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[5]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~8_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[5]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~8_combout ),
	.cin(gnd),
	.combout(\ramaddr~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~9 .lut_mask = 16'hDD88;
defparam \ramaddr~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N16
cycloneive_lcell_comb \ramaddr~10 (
// Equation(s):
// \ramaddr~10_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[4]~input_o )) # (!\syif.tbCTRL~input_o  & (((!exmem_ifdREN_o & !exmem_ifdWEN_o))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[4]~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~10 .lut_mask = 16'h888D;
defparam \ramaddr~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N18
cycloneive_lcell_comb \ramaddr~11 (
// Equation(s):
// \ramaddr~11_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~10_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~10_combout  & ((pc_4))) # (!\ramaddr~10_combout  & (exmem_ifout_o_4))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|EXMEM|exmem_if.out_o [4]),
	.datac(\CPU|DP|pc [4]),
	.datad(\ramaddr~10_combout ),
	.cin(gnd),
	.combout(\ramaddr~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~11 .lut_mask = 16'hFA44;
defparam \ramaddr~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N6
cycloneive_lcell_comb \ramaddr~12 (
// Equation(s):
// \ramaddr~12_combout  = (exmem_ifdWEN_o & (exmem_ifout_o_7)) # (!exmem_ifdWEN_o & ((exmem_ifdREN_o & (exmem_ifout_o_7)) # (!exmem_ifdREN_o & ((pc_7)))))

	.dataa(\CPU|DP|EXMEM|exmem_if.out_o [7]),
	.datab(\CPU|DP|pc [7]),
	.datac(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~12 .lut_mask = 16'hAAAC;
defparam \ramaddr~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N20
cycloneive_lcell_comb \ramaddr~13 (
// Equation(s):
// \ramaddr~13_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[7]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~12_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[7]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~12_combout ),
	.cin(gnd),
	.combout(\ramaddr~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~13 .lut_mask = 16'hDD88;
defparam \ramaddr~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N0
cycloneive_lcell_comb \ramaddr~14 (
// Equation(s):
// \ramaddr~14_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[6]~input_o )) # (!\syif.tbCTRL~input_o  & (((exmem_ifdWEN_o) # (exmem_ifdREN_o))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[6]~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~14 .lut_mask = 16'hDDD8;
defparam \ramaddr~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N18
cycloneive_lcell_comb \ramaddr~15 (
// Equation(s):
// \ramaddr~15_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~14_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~14_combout  & ((exmem_ifout_o_6))) # (!\ramaddr~14_combout  & (pc_6))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|pc [6]),
	.datac(\CPU|DP|EXMEM|exmem_if.out_o [6]),
	.datad(\ramaddr~14_combout ),
	.cin(gnd),
	.combout(\ramaddr~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~15 .lut_mask = 16'hFA44;
defparam \ramaddr~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N2
cycloneive_lcell_comb \ramaddr~16 (
// Equation(s):
// \ramaddr~16_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[9]~input_o )) # (!\syif.tbCTRL~input_o  & (((exmem_ifdWEN_o) # (exmem_ifdREN_o))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[9]~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~16 .lut_mask = 16'hDDD8;
defparam \ramaddr~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N8
cycloneive_lcell_comb \ramaddr~17 (
// Equation(s):
// \ramaddr~17_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~16_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~16_combout  & (exmem_ifout_o_9)) # (!\ramaddr~16_combout  & ((pc_9)))))

	.dataa(\CPU|DP|EXMEM|exmem_if.out_o [9]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|pc [9]),
	.datad(\ramaddr~16_combout ),
	.cin(gnd),
	.combout(\ramaddr~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~17 .lut_mask = 16'hEE30;
defparam \ramaddr~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N0
cycloneive_lcell_comb \ramaddr~18 (
// Equation(s):
// \ramaddr~18_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[8]~input_o )) # (!\syif.tbCTRL~input_o  & (((!exmem_ifdWEN_o & !exmem_ifdREN_o))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[8]~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~18 .lut_mask = 16'h888D;
defparam \ramaddr~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N18
cycloneive_lcell_comb \ramaddr~19 (
// Equation(s):
// \ramaddr~19_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~18_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~18_combout  & ((pc_8))) # (!\ramaddr~18_combout  & (exmem_ifout_o_8))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|EXMEM|exmem_if.out_o [8]),
	.datac(\CPU|DP|pc [8]),
	.datad(\ramaddr~18_combout ),
	.cin(gnd),
	.combout(\ramaddr~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~19 .lut_mask = 16'hFA44;
defparam \ramaddr~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N6
cycloneive_lcell_comb \ramaddr~20 (
// Equation(s):
// \ramaddr~20_combout  = (exmem_ifdREN_o & (((exmem_ifout_o_11)))) # (!exmem_ifdREN_o & ((exmem_ifdWEN_o & ((exmem_ifout_o_11))) # (!exmem_ifdWEN_o & (pc_11))))

	.dataa(\CPU|DP|pc [11]),
	.datab(\CPU|DP|EXMEM|exmem_if.out_o [11]),
	.datac(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~20 .lut_mask = 16'hCCCA;
defparam \ramaddr~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N20
cycloneive_lcell_comb \ramaddr~21 (
// Equation(s):
// \ramaddr~21_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[11]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~20_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[11]~input_o ),
	.datad(\ramaddr~20_combout ),
	.cin(gnd),
	.combout(\ramaddr~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~21 .lut_mask = 16'hF3C0;
defparam \ramaddr~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N16
cycloneive_lcell_comb \ramaddr~22 (
// Equation(s):
// \ramaddr~22_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[10]~input_o )) # (!\syif.tbCTRL~input_o  & (((exmem_ifdREN_o) # (exmem_ifdWEN_o))))

	.dataa(\syif.addr[10]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~22 .lut_mask = 16'hBBB8;
defparam \ramaddr~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N2
cycloneive_lcell_comb \ramaddr~23 (
// Equation(s):
// \ramaddr~23_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~22_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~22_combout  & ((exmem_ifout_o_10))) # (!\ramaddr~22_combout  & (pc_10))))

	.dataa(\CPU|DP|pc [10]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.out_o [10]),
	.datad(\ramaddr~22_combout ),
	.cin(gnd),
	.combout(\ramaddr~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~23 .lut_mask = 16'hFC22;
defparam \ramaddr~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N20
cycloneive_lcell_comb \ramaddr~24 (
// Equation(s):
// \ramaddr~24_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[13]~input_o )))) # (!\syif.tbCTRL~input_o  & (!exmem_ifdREN_o & (!exmem_ifdWEN_o)))

	.dataa(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datad(\syif.addr[13]~input_o ),
	.cin(gnd),
	.combout(\ramaddr~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~24 .lut_mask = 16'hCD01;
defparam \ramaddr~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N10
cycloneive_lcell_comb \ramaddr~25 (
// Equation(s):
// \ramaddr~25_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~24_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~24_combout  & ((pc_13))) # (!\ramaddr~24_combout  & (exmem_ifout_o_13))))

	.dataa(\CPU|DP|EXMEM|exmem_if.out_o [13]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|pc [13]),
	.datad(\ramaddr~24_combout ),
	.cin(gnd),
	.combout(\ramaddr~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~25 .lut_mask = 16'hFC22;
defparam \ramaddr~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N28
cycloneive_lcell_comb \ramaddr~26 (
// Equation(s):
// \ramaddr~26_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[12]~input_o )))) # (!\syif.tbCTRL~input_o  & (!exmem_ifdREN_o & ((!exmem_ifdWEN_o))))

	.dataa(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datab(\syif.addr[12]~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramaddr~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~26 .lut_mask = 16'hCC05;
defparam \ramaddr~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N18
cycloneive_lcell_comb \ramaddr~27 (
// Equation(s):
// \ramaddr~27_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~26_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~26_combout  & (pc_12)) # (!\ramaddr~26_combout  & ((exmem_ifout_o_12)))))

	.dataa(\CPU|DP|pc [12]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.out_o [12]),
	.datad(\ramaddr~26_combout ),
	.cin(gnd),
	.combout(\ramaddr~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~27 .lut_mask = 16'hEE30;
defparam \ramaddr~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N10
cycloneive_lcell_comb \ramaddr~28 (
// Equation(s):
// \ramaddr~28_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[15]~input_o )) # (!\syif.tbCTRL~input_o  & (((exmem_ifdWEN_o) # (exmem_ifdREN_o))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[15]~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~28 .lut_mask = 16'hDDD8;
defparam \ramaddr~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N20
cycloneive_lcell_comb \ramaddr~29 (
// Equation(s):
// \ramaddr~29_combout  = (\syif.tbCTRL~input_o  & (((!\ramaddr~28_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~28_combout  & (!exmem_ifout_o_15)) # (!\ramaddr~28_combout  & ((!pc_15)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|EXMEM|exmem_if.out_o [15]),
	.datac(\CPU|DP|pc [15]),
	.datad(\ramaddr~28_combout ),
	.cin(gnd),
	.combout(\ramaddr~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~29 .lut_mask = 16'h11AF;
defparam \ramaddr~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N14
cycloneive_lcell_comb \ramaddr~30 (
// Equation(s):
// \ramaddr~30_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[14]~input_o )) # (!\syif.tbCTRL~input_o  & (((!exmem_ifdWEN_o & !exmem_ifdREN_o))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[14]~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~30 .lut_mask = 16'h888D;
defparam \ramaddr~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N4
cycloneive_lcell_comb \ramaddr~31 (
// Equation(s):
// \ramaddr~31_combout  = (\syif.tbCTRL~input_o  & (\ramaddr~30_combout )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~30_combout  & (pc_14)) # (!\ramaddr~30_combout  & ((exmem_ifout_o_14)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\ramaddr~30_combout ),
	.datac(\CPU|DP|pc [14]),
	.datad(\CPU|DP|EXMEM|exmem_if.out_o [14]),
	.cin(gnd),
	.combout(\ramaddr~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~31 .lut_mask = 16'hD9C8;
defparam \ramaddr~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N6
cycloneive_lcell_comb \ramaddr~32 (
// Equation(s):
// \ramaddr~32_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[17]~input_o )))) # (!\syif.tbCTRL~input_o  & (!exmem_ifdREN_o & ((!exmem_ifdWEN_o))))

	.dataa(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datab(\syif.addr[17]~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramaddr~32_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~32 .lut_mask = 16'hCC05;
defparam \ramaddr~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N30
cycloneive_lcell_comb \ramaddr~33 (
// Equation(s):
// \ramaddr~33_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~32_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~32_combout  & ((pc_17))) # (!\ramaddr~32_combout  & (exmem_ifout_o_17))))

	.dataa(\CPU|DP|EXMEM|exmem_if.out_o [17]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|pc [17]),
	.datad(\ramaddr~32_combout ),
	.cin(gnd),
	.combout(\ramaddr~33_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~33 .lut_mask = 16'hFC22;
defparam \ramaddr~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N2
cycloneive_lcell_comb \ramaddr~34 (
// Equation(s):
// \ramaddr~34_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[16]~input_o )))) # (!\syif.tbCTRL~input_o  & ((exmem_ifdREN_o) # ((exmem_ifdWEN_o))))

	.dataa(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datad(\syif.addr[16]~input_o ),
	.cin(gnd),
	.combout(\ramaddr~34_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~34 .lut_mask = 16'hFE32;
defparam \ramaddr~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N16
cycloneive_lcell_comb \ramaddr~35 (
// Equation(s):
// \ramaddr~35_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~34_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~34_combout  & (exmem_ifout_o_16)) # (!\ramaddr~34_combout  & ((pc_16)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|EXMEM|exmem_if.out_o [16]),
	.datac(\CPU|DP|pc [16]),
	.datad(\ramaddr~34_combout ),
	.cin(gnd),
	.combout(\ramaddr~35_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~35 .lut_mask = 16'hEE50;
defparam \ramaddr~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N20
cycloneive_lcell_comb \ramaddr~36 (
// Equation(s):
// \ramaddr~36_combout  = (exmem_ifdWEN_o & (((exmem_ifout_o_19)))) # (!exmem_ifdWEN_o & ((exmem_ifdREN_o & ((exmem_ifout_o_19))) # (!exmem_ifdREN_o & (pc_19))))

	.dataa(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datab(\CPU|DP|pc [19]),
	.datac(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.out_o [19]),
	.cin(gnd),
	.combout(\ramaddr~36_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~36 .lut_mask = 16'hFE04;
defparam \ramaddr~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N22
cycloneive_lcell_comb \ramaddr~37 (
// Equation(s):
// \ramaddr~37_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[19]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~36_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[19]~input_o ),
	.datad(\ramaddr~36_combout ),
	.cin(gnd),
	.combout(\ramaddr~37_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~37 .lut_mask = 16'hF3C0;
defparam \ramaddr~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N12
cycloneive_lcell_comb \ramaddr~38 (
// Equation(s):
// \ramaddr~38_combout  = (exmem_ifdREN_o & (exmem_ifout_o_18)) # (!exmem_ifdREN_o & ((exmem_ifdWEN_o & (exmem_ifout_o_18)) # (!exmem_ifdWEN_o & ((pc_18)))))

	.dataa(\CPU|DP|EXMEM|exmem_if.out_o [18]),
	.datab(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datac(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datad(\CPU|DP|pc [18]),
	.cin(gnd),
	.combout(\ramaddr~38_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~38 .lut_mask = 16'hABA8;
defparam \ramaddr~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N2
cycloneive_lcell_comb \ramaddr~39 (
// Equation(s):
// \ramaddr~39_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[18]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~38_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[18]~input_o ),
	.datad(\ramaddr~38_combout ),
	.cin(gnd),
	.combout(\ramaddr~39_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~39 .lut_mask = 16'hF3C0;
defparam \ramaddr~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N12
cycloneive_lcell_comb \ramaddr~40 (
// Equation(s):
// \ramaddr~40_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[21]~input_o )) # (!\syif.tbCTRL~input_o  & (((!exmem_ifdREN_o & !exmem_ifdWEN_o))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[21]~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~40_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~40 .lut_mask = 16'h888D;
defparam \ramaddr~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N18
cycloneive_lcell_comb \ramaddr~41 (
// Equation(s):
// \ramaddr~41_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~40_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~40_combout  & ((pc_21))) # (!\ramaddr~40_combout  & (exmem_ifout_o_21))))

	.dataa(\CPU|DP|EXMEM|exmem_if.out_o [21]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|pc [21]),
	.datad(\ramaddr~40_combout ),
	.cin(gnd),
	.combout(\ramaddr~41_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~41 .lut_mask = 16'hFC22;
defparam \ramaddr~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N0
cycloneive_lcell_comb \ramaddr~42 (
// Equation(s):
// \ramaddr~42_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[20]~input_o )) # (!\syif.tbCTRL~input_o  & (((!exmem_ifdREN_o & !exmem_ifdWEN_o))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[20]~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~42_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~42 .lut_mask = 16'h888D;
defparam \ramaddr~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N2
cycloneive_lcell_comb \ramaddr~43 (
// Equation(s):
// \ramaddr~43_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~42_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~42_combout  & ((pc_20))) # (!\ramaddr~42_combout  & (exmem_ifout_o_20))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|EXMEM|exmem_if.out_o [20]),
	.datac(\CPU|DP|pc [20]),
	.datad(\ramaddr~42_combout ),
	.cin(gnd),
	.combout(\ramaddr~43_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~43 .lut_mask = 16'hFA44;
defparam \ramaddr~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N18
cycloneive_lcell_comb \ramaddr~44 (
// Equation(s):
// \ramaddr~44_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[23]~input_o )))) # (!\syif.tbCTRL~input_o  & ((exmem_ifdWEN_o) # ((exmem_ifdREN_o))))

	.dataa(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datab(\syif.addr[23]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~44_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~44 .lut_mask = 16'hCFCA;
defparam \ramaddr~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N10
cycloneive_lcell_comb \ramaddr~45 (
// Equation(s):
// \ramaddr~45_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~44_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~44_combout  & (exmem_ifout_o_23)) # (!\ramaddr~44_combout  & ((pc_23)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|EXMEM|exmem_if.out_o [23]),
	.datac(\CPU|DP|pc [23]),
	.datad(\ramaddr~44_combout ),
	.cin(gnd),
	.combout(\ramaddr~45_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~45 .lut_mask = 16'hEE50;
defparam \ramaddr~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N26
cycloneive_lcell_comb \ramaddr~46 (
// Equation(s):
// \ramaddr~46_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[22]~input_o )))) # (!\syif.tbCTRL~input_o  & ((exmem_ifdWEN_o) # ((exmem_ifdREN_o))))

	.dataa(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datab(\syif.addr[22]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~46_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~46 .lut_mask = 16'hCFCA;
defparam \ramaddr~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N0
cycloneive_lcell_comb \ramaddr~47 (
// Equation(s):
// \ramaddr~47_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~46_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~46_combout  & (exmem_ifout_o_22)) # (!\ramaddr~46_combout  & ((pc_22)))))

	.dataa(\CPU|DP|EXMEM|exmem_if.out_o [22]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramaddr~46_combout ),
	.datad(\CPU|DP|pc [22]),
	.cin(gnd),
	.combout(\ramaddr~47_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~47 .lut_mask = 16'hE3E0;
defparam \ramaddr~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N0
cycloneive_lcell_comb \ramaddr~48 (
// Equation(s):
// \ramaddr~48_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[25]~input_o )) # (!\syif.tbCTRL~input_o  & (((!exmem_ifdREN_o & !exmem_ifdWEN_o))))

	.dataa(\syif.addr[25]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~48_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~48 .lut_mask = 16'h888B;
defparam \ramaddr~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N6
cycloneive_lcell_comb \ramaddr~49 (
// Equation(s):
// \ramaddr~49_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~48_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~48_combout  & ((pc_25))) # (!\ramaddr~48_combout  & (exmem_ifout_o_25))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|EXMEM|exmem_if.out_o [25]),
	.datac(\CPU|DP|pc [25]),
	.datad(\ramaddr~48_combout ),
	.cin(gnd),
	.combout(\ramaddr~49_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~49 .lut_mask = 16'hFA44;
defparam \ramaddr~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N28
cycloneive_lcell_comb \ramaddr~50 (
// Equation(s):
// \ramaddr~50_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[24]~input_o )) # (!\syif.tbCTRL~input_o  & (((!exmem_ifdREN_o & !exmem_ifdWEN_o))))

	.dataa(\syif.addr[24]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~50_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~50 .lut_mask = 16'h888B;
defparam \ramaddr~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N10
cycloneive_lcell_comb \ramaddr~51 (
// Equation(s):
// \ramaddr~51_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~50_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~50_combout  & (pc_24)) # (!\ramaddr~50_combout  & ((exmem_ifout_o_24)))))

	.dataa(\CPU|DP|pc [24]),
	.datab(\CPU|DP|EXMEM|exmem_if.out_o [24]),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~50_combout ),
	.cin(gnd),
	.combout(\ramaddr~51_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~51 .lut_mask = 16'hFA0C;
defparam \ramaddr~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N18
cycloneive_lcell_comb \ramaddr~52 (
// Equation(s):
// \ramaddr~52_combout  = (exmem_ifdWEN_o & (((exmem_ifout_o_27)))) # (!exmem_ifdWEN_o & ((exmem_ifdREN_o & ((exmem_ifout_o_27))) # (!exmem_ifdREN_o & (pc_27))))

	.dataa(\CPU|DP|pc [27]),
	.datab(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datac(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.out_o [27]),
	.cin(gnd),
	.combout(\ramaddr~52_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~52 .lut_mask = 16'hFE02;
defparam \ramaddr~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N2
cycloneive_lcell_comb \ramaddr~53 (
// Equation(s):
// \ramaddr~53_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[27]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~52_combout )))

	.dataa(\syif.addr[27]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~52_combout ),
	.cin(gnd),
	.combout(\ramaddr~53_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~53 .lut_mask = 16'hBB88;
defparam \ramaddr~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N30
cycloneive_lcell_comb \ramaddr~54 (
// Equation(s):
// \ramaddr~54_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[26]~input_o )) # (!\syif.tbCTRL~input_o  & (((exmem_ifdREN_o) # (exmem_ifdWEN_o))))

	.dataa(\syif.addr[26]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~54_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~54 .lut_mask = 16'hBBB8;
defparam \ramaddr~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N20
cycloneive_lcell_comb \ramaddr~55 (
// Equation(s):
// \ramaddr~55_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~54_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~54_combout  & ((exmem_ifout_o_26))) # (!\ramaddr~54_combout  & (pc_26))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|pc [26]),
	.datac(\ramaddr~54_combout ),
	.datad(\CPU|DP|EXMEM|exmem_if.out_o [26]),
	.cin(gnd),
	.combout(\ramaddr~55_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~55 .lut_mask = 16'hF4A4;
defparam \ramaddr~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N30
cycloneive_lcell_comb \ramaddr~56 (
// Equation(s):
// \ramaddr~56_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[29]~input_o )))) # (!\syif.tbCTRL~input_o  & (!exmem_ifdWEN_o & ((!exmem_ifdREN_o))))

	.dataa(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datab(\syif.addr[29]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~56_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~56 .lut_mask = 16'hC0C5;
defparam \ramaddr~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N20
cycloneive_lcell_comb \ramaddr~57 (
// Equation(s):
// \ramaddr~57_combout  = (\ramaddr~56_combout  & ((\syif.tbCTRL~input_o ) # ((pc_29)))) # (!\ramaddr~56_combout  & (!\syif.tbCTRL~input_o  & ((exmem_ifout_o_29))))

	.dataa(\ramaddr~56_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|pc [29]),
	.datad(\CPU|DP|EXMEM|exmem_if.out_o [29]),
	.cin(gnd),
	.combout(\ramaddr~57_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~57 .lut_mask = 16'hB9A8;
defparam \ramaddr~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N24
cycloneive_lcell_comb \ramaddr~58 (
// Equation(s):
// \ramaddr~58_combout  = (exmem_ifdWEN_o & (((exmem_ifout_o_28)))) # (!exmem_ifdWEN_o & ((exmem_ifdREN_o & (exmem_ifout_o_28)) # (!exmem_ifdREN_o & ((pc_28)))))

	.dataa(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datab(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datac(\CPU|DP|EXMEM|exmem_if.out_o [28]),
	.datad(\CPU|DP|pc [28]),
	.cin(gnd),
	.combout(\ramaddr~58_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~58 .lut_mask = 16'hF1E0;
defparam \ramaddr~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N2
cycloneive_lcell_comb \ramaddr~59 (
// Equation(s):
// \ramaddr~59_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[28]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~58_combout )))

	.dataa(\syif.addr[28]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~58_combout ),
	.cin(gnd),
	.combout(\ramaddr~59_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~59 .lut_mask = 16'hBB88;
defparam \ramaddr~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N24
cycloneive_lcell_comb \ramaddr~60 (
// Equation(s):
// \ramaddr~60_combout  = (exmem_ifdWEN_o & (exmem_ifout_o_31)) # (!exmem_ifdWEN_o & ((exmem_ifdREN_o & (exmem_ifout_o_31)) # (!exmem_ifdREN_o & ((pc_31)))))

	.dataa(\CPU|DP|EXMEM|exmem_if.out_o [31]),
	.datab(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datac(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.datad(\CPU|DP|pc [31]),
	.cin(gnd),
	.combout(\ramaddr~60_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~60 .lut_mask = 16'hABA8;
defparam \ramaddr~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N18
cycloneive_lcell_comb \ramaddr~61 (
// Equation(s):
// \ramaddr~61_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[31]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~60_combout )))

	.dataa(\syif.addr[31]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~60_combout ),
	.cin(gnd),
	.combout(\ramaddr~61_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~61 .lut_mask = 16'hBB88;
defparam \ramaddr~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N8
cycloneive_lcell_comb \ramaddr~62 (
// Equation(s):
// \ramaddr~62_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[30]~input_o )) # (!\syif.tbCTRL~input_o  & (((exmem_ifdWEN_o) # (exmem_ifdREN_o))))

	.dataa(\syif.addr[30]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datad(\CPU|DP|EXMEM|exmem_if.dREN_o~q ),
	.cin(gnd),
	.combout(\ramaddr~62_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~62 .lut_mask = 16'hBBB8;
defparam \ramaddr~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N6
cycloneive_lcell_comb \ramaddr~63 (
// Equation(s):
// \ramaddr~63_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~62_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~62_combout  & (exmem_ifout_o_30)) # (!\ramaddr~62_combout  & ((pc_30)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|EXMEM|exmem_if.out_o [30]),
	.datac(\ramaddr~62_combout ),
	.datad(\CPU|DP|pc [30]),
	.cin(gnd),
	.combout(\ramaddr~63_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~63 .lut_mask = 16'hE5E0;
defparam \ramaddr~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y1_N25
dffeas CPUCLK(
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\CPUCLK~0_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\CPUCLK~q ),
	.prn(vcc));
// synopsys translate_off
defparam CPUCLK.is_wysiwyg = "true";
defparam CPUCLK.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N20
cycloneive_lcell_comb \ramWEN~0 (
// Equation(s):
// \ramWEN~0_combout  = (\syif.tbCTRL~input_o  & (!\syif.WEN~input_o )) # (!\syif.tbCTRL~input_o  & ((!exmem_ifdWEN_o)))

	.dataa(gnd),
	.datab(\syif.WEN~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramWEN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramWEN~0 .lut_mask = 16'h330F;
defparam \ramWEN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N2
cycloneive_lcell_comb \ramstore~0 (
// Equation(s):
// \ramstore~0_combout  = (\syif.tbCTRL~input_o  & (\syif.store[0]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_0)))

	.dataa(\syif.store[0]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [0]),
	.cin(gnd),
	.combout(\ramstore~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~0 .lut_mask = 16'hBB88;
defparam \ramstore~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N30
cycloneive_lcell_comb \ramREN~0 (
// Equation(s):
// \ramREN~0_combout  = (\syif.tbCTRL~input_o  & ((!\syif.REN~input_o ))) # (!\syif.tbCTRL~input_o  & (exmem_ifdWEN_o))

	.dataa(gnd),
	.datab(\CPU|DP|EXMEM|exmem_if.dWEN_o~q ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\syif.REN~input_o ),
	.cin(gnd),
	.combout(\ramREN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramREN~0 .lut_mask = 16'h0CFC;
defparam \ramREN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N16
cycloneive_lcell_comb \ramstore~1 (
// Equation(s):
// \ramstore~1_combout  = (\syif.tbCTRL~input_o  & (\syif.store[1]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_1)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[1]~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [1]),
	.cin(gnd),
	.combout(\ramstore~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~1 .lut_mask = 16'hF3C0;
defparam \ramstore~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N10
cycloneive_lcell_comb \ramstore~2 (
// Equation(s):
// \ramstore~2_combout  = (\syif.tbCTRL~input_o  & (\syif.store[2]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_2)))

	.dataa(\syif.store[2]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [2]),
	.cin(gnd),
	.combout(\ramstore~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~2 .lut_mask = 16'hBB88;
defparam \ramstore~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N6
cycloneive_lcell_comb \ramstore~3 (
// Equation(s):
// \ramstore~3_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[3]~input_o ))) # (!\syif.tbCTRL~input_o  & (exmem_ifrdat2_o_3))

	.dataa(\CPU|DP|EXMEM|exmem_if.rdat2_o [3]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\syif.store[3]~input_o ),
	.cin(gnd),
	.combout(\ramstore~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~3 .lut_mask = 16'hEE22;
defparam \ramstore~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N22
cycloneive_lcell_comb \ramstore~4 (
// Equation(s):
// \ramstore~4_combout  = (\syif.tbCTRL~input_o  & (\syif.store[4]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_4)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[4]~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [4]),
	.cin(gnd),
	.combout(\ramstore~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~4 .lut_mask = 16'hF5A0;
defparam \ramstore~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N8
cycloneive_lcell_comb \ramstore~5 (
// Equation(s):
// \ramstore~5_combout  = (\syif.tbCTRL~input_o  & (\syif.store[5]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_5)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[5]~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [5]),
	.cin(gnd),
	.combout(\ramstore~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~5 .lut_mask = 16'hF5A0;
defparam \ramstore~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N24
cycloneive_lcell_comb \ramstore~6 (
// Equation(s):
// \ramstore~6_combout  = (\syif.tbCTRL~input_o  & (\syif.store[6]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_6)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[6]~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [6]),
	.cin(gnd),
	.combout(\ramstore~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~6 .lut_mask = 16'hF5A0;
defparam \ramstore~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N24
cycloneive_lcell_comb \ramstore~7 (
// Equation(s):
// \ramstore~7_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[7]~input_o ))) # (!\syif.tbCTRL~input_o  & (exmem_ifrdat2_o_7))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|EXMEM|exmem_if.rdat2_o [7]),
	.datac(gnd),
	.datad(\syif.store[7]~input_o ),
	.cin(gnd),
	.combout(\ramstore~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~7 .lut_mask = 16'hEE44;
defparam \ramstore~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N8
cycloneive_lcell_comb \ramstore~8 (
// Equation(s):
// \ramstore~8_combout  = (\syif.tbCTRL~input_o  & (\syif.store[8]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_8)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[8]~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [8]),
	.cin(gnd),
	.combout(\ramstore~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~8 .lut_mask = 16'hF5A0;
defparam \ramstore~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N30
cycloneive_lcell_comb \ramstore~9 (
// Equation(s):
// \ramstore~9_combout  = (\syif.tbCTRL~input_o  & (\syif.store[9]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_9)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[9]~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [9]),
	.cin(gnd),
	.combout(\ramstore~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~9 .lut_mask = 16'hF5A0;
defparam \ramstore~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y16_N0
cycloneive_lcell_comb \ramstore~10 (
// Equation(s):
// \ramstore~10_combout  = (\syif.tbCTRL~input_o  & (\syif.store[10]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_10)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[10]~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [10]),
	.cin(gnd),
	.combout(\ramstore~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~10 .lut_mask = 16'hF3C0;
defparam \ramstore~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N14
cycloneive_lcell_comb \ramstore~11 (
// Equation(s):
// \ramstore~11_combout  = (\syif.tbCTRL~input_o  & (\syif.store[11]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_11)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[11]~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [11]),
	.cin(gnd),
	.combout(\ramstore~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~11 .lut_mask = 16'hF5A0;
defparam \ramstore~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N22
cycloneive_lcell_comb \ramstore~12 (
// Equation(s):
// \ramstore~12_combout  = (\syif.tbCTRL~input_o  & (\syif.store[12]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_12)))

	.dataa(\syif.store[12]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [12]),
	.cin(gnd),
	.combout(\ramstore~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~12 .lut_mask = 16'hBB88;
defparam \ramstore~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y24_N28
cycloneive_lcell_comb \ramstore~13 (
// Equation(s):
// \ramstore~13_combout  = (\syif.tbCTRL~input_o  & (\syif.store[13]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_13)))

	.dataa(\syif.store[13]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [13]),
	.cin(gnd),
	.combout(\ramstore~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~13 .lut_mask = 16'hAFA0;
defparam \ramstore~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N14
cycloneive_lcell_comb \ramstore~14 (
// Equation(s):
// \ramstore~14_combout  = (\syif.tbCTRL~input_o  & (\syif.store[14]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_14)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[14]~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [14]),
	.cin(gnd),
	.combout(\ramstore~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~14 .lut_mask = 16'hDD88;
defparam \ramstore~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N16
cycloneive_lcell_comb \ramstore~15 (
// Equation(s):
// \ramstore~15_combout  = (\syif.tbCTRL~input_o  & (\syif.store[15]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_15)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[15]~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [15]),
	.cin(gnd),
	.combout(\ramstore~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~15 .lut_mask = 16'hDD88;
defparam \ramstore~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N10
cycloneive_lcell_comb \ramstore~16 (
// Equation(s):
// \ramstore~16_combout  = (\syif.tbCTRL~input_o  & (\syif.store[16]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_16)))

	.dataa(\syif.store[16]~input_o ),
	.datab(\CPU|DP|EXMEM|exmem_if.rdat2_o [16]),
	.datac(gnd),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~16 .lut_mask = 16'hAACC;
defparam \ramstore~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N4
cycloneive_lcell_comb \ramstore~17 (
// Equation(s):
// \ramstore~17_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[17]~input_o ))) # (!\syif.tbCTRL~input_o  & (exmem_ifrdat2_o_17))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|EXMEM|exmem_if.rdat2_o [17]),
	.datac(\syif.store[17]~input_o ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramstore~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~17 .lut_mask = 16'hE4E4;
defparam \ramstore~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N6
cycloneive_lcell_comb \ramstore~18 (
// Equation(s):
// \ramstore~18_combout  = (\syif.tbCTRL~input_o  & (\syif.store[18]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_18)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[18]~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [18]),
	.cin(gnd),
	.combout(\ramstore~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~18 .lut_mask = 16'hF5A0;
defparam \ramstore~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y24_N26
cycloneive_lcell_comb \ramstore~19 (
// Equation(s):
// \ramstore~19_combout  = (\syif.tbCTRL~input_o  & (\syif.store[19]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_19)))

	.dataa(gnd),
	.datab(\syif.store[19]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [19]),
	.cin(gnd),
	.combout(\ramstore~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~19 .lut_mask = 16'hCFC0;
defparam \ramstore~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N2
cycloneive_lcell_comb \ramstore~20 (
// Equation(s):
// \ramstore~20_combout  = (\syif.tbCTRL~input_o  & (\syif.store[20]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_20)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[20]~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [20]),
	.cin(gnd),
	.combout(\ramstore~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~20 .lut_mask = 16'hF5A0;
defparam \ramstore~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N16
cycloneive_lcell_comb \ramstore~21 (
// Equation(s):
// \ramstore~21_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[21]~input_o ))) # (!\syif.tbCTRL~input_o  & (exmem_ifrdat2_o_21))

	.dataa(gnd),
	.datab(\CPU|DP|EXMEM|exmem_if.rdat2_o [21]),
	.datac(\syif.store[21]~input_o ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~21 .lut_mask = 16'hF0CC;
defparam \ramstore~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N24
cycloneive_lcell_comb \ramstore~22 (
// Equation(s):
// \ramstore~22_combout  = (\syif.tbCTRL~input_o  & (\syif.store[22]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_22)))

	.dataa(gnd),
	.datab(\syif.store[22]~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.rdat2_o [22]),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~22 .lut_mask = 16'hCCF0;
defparam \ramstore~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N14
cycloneive_lcell_comb \ramstore~23 (
// Equation(s):
// \ramstore~23_combout  = (\syif.tbCTRL~input_o  & (\syif.store[23]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_23)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[23]~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [23]),
	.cin(gnd),
	.combout(\ramstore~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~23 .lut_mask = 16'hF5A0;
defparam \ramstore~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N26
cycloneive_lcell_comb \ramstore~24 (
// Equation(s):
// \ramstore~24_combout  = (\syif.tbCTRL~input_o  & (\syif.store[24]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_24)))

	.dataa(\syif.store[24]~input_o ),
	.datab(gnd),
	.datac(\CPU|DP|EXMEM|exmem_if.rdat2_o [24]),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~24 .lut_mask = 16'hAAF0;
defparam \ramstore~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N8
cycloneive_lcell_comb \ramstore~25 (
// Equation(s):
// \ramstore~25_combout  = (\syif.tbCTRL~input_o  & (\syif.store[25]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_25)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[25]~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [25]),
	.cin(gnd),
	.combout(\ramstore~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~25 .lut_mask = 16'hF3C0;
defparam \ramstore~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N28
cycloneive_lcell_comb \ramstore~26 (
// Equation(s):
// \ramstore~26_combout  = (\syif.tbCTRL~input_o  & (\syif.store[26]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_26)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[26]~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [26]),
	.cin(gnd),
	.combout(\ramstore~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~26 .lut_mask = 16'hF3C0;
defparam \ramstore~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N22
cycloneive_lcell_comb \ramstore~27 (
// Equation(s):
// \ramstore~27_combout  = (\syif.tbCTRL~input_o  & (\syif.store[27]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_27)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[27]~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [27]),
	.cin(gnd),
	.combout(\ramstore~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~27 .lut_mask = 16'hF3C0;
defparam \ramstore~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N4
cycloneive_lcell_comb \ramstore~28 (
// Equation(s):
// \ramstore~28_combout  = (\syif.tbCTRL~input_o  & (\syif.store[28]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_28)))

	.dataa(\syif.store[28]~input_o ),
	.datab(gnd),
	.datac(\CPU|DP|EXMEM|exmem_if.rdat2_o [28]),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~28 .lut_mask = 16'hAAF0;
defparam \ramstore~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N12
cycloneive_lcell_comb \ramstore~29 (
// Equation(s):
// \ramstore~29_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[29]~input_o ))) # (!\syif.tbCTRL~input_o  & (exmem_ifrdat2_o_29))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.rdat2_o [29]),
	.datad(\syif.store[29]~input_o ),
	.cin(gnd),
	.combout(\ramstore~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~29 .lut_mask = 16'hFC30;
defparam \ramstore~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N18
cycloneive_lcell_comb \ramstore~30 (
// Equation(s):
// \ramstore~30_combout  = (\syif.tbCTRL~input_o  & (\syif.store[30]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_30)))

	.dataa(gnd),
	.datab(\syif.store[30]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|EXMEM|exmem_if.rdat2_o [30]),
	.cin(gnd),
	.combout(\ramstore~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~30 .lut_mask = 16'hCFC0;
defparam \ramstore~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N22
cycloneive_lcell_comb \ramstore~31 (
// Equation(s):
// \ramstore~31_combout  = (\syif.tbCTRL~input_o  & (\syif.store[31]~input_o )) # (!\syif.tbCTRL~input_o  & ((exmem_ifrdat2_o_31)))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[31]~input_o ),
	.datac(\CPU|DP|EXMEM|exmem_if.rdat2_o [31]),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramstore~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~31 .lut_mask = 16'hD8D8;
defparam \ramstore~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y1_N1
dffeas \count[3] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[3]~0_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[3]),
	.prn(vcc));
// synopsys translate_off
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y1_N23
dffeas \count[2] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[2]~1_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[2]),
	.prn(vcc));
// synopsys translate_off
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y1_N13
dffeas \count[1] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[1]~2_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[1]),
	.prn(vcc));
// synopsys translate_off
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y1_N3
dffeas \count[0] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[0]),
	.prn(vcc));
// synopsys translate_off
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y1_N24
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (!count[1] & (!count[0] & (!count[2] & !count[3])))

	.dataa(count[1]),
	.datab(count[0]),
	.datac(count[2]),
	.datad(count[3]),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h0001;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y1_N24
cycloneive_lcell_comb \CPUCLK~0 (
// Equation(s):
// \CPUCLK~0_combout  = \CPUCLK~q  $ (\Equal0~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\CPUCLK~q ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\CPUCLK~0_combout ),
	.cout());
// synopsys translate_off
defparam \CPUCLK~0 .lut_mask = 16'h0FF0;
defparam \CPUCLK~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y1_N0
cycloneive_lcell_comb \count[3]~0 (
// Equation(s):
// \count[3]~0_combout  = count[3] $ (((count[2] & (count[0] & count[1]))))

	.dataa(count[2]),
	.datab(count[0]),
	.datac(count[3]),
	.datad(count[1]),
	.cin(gnd),
	.combout(\count[3]~0_combout ),
	.cout());
// synopsys translate_off
defparam \count[3]~0 .lut_mask = 16'h78F0;
defparam \count[3]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y1_N22
cycloneive_lcell_comb \count[2]~1 (
// Equation(s):
// \count[2]~1_combout  = count[2] $ (((count[0] & count[1])))

	.dataa(gnd),
	.datab(count[0]),
	.datac(count[2]),
	.datad(count[1]),
	.cin(gnd),
	.combout(\count[2]~1_combout ),
	.cout());
// synopsys translate_off
defparam \count[2]~1 .lut_mask = 16'h3CF0;
defparam \count[2]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y1_N12
cycloneive_lcell_comb \count[1]~2 (
// Equation(s):
// \count[1]~2_combout  = count[1] $ (count[0])

	.dataa(gnd),
	.datab(gnd),
	.datac(count[1]),
	.datad(count[0]),
	.cin(gnd),
	.combout(\count[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \count[1]~2 .lut_mask = 16'h0FF0;
defparam \count[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y1_N2
cycloneive_lcell_comb \count~3 (
// Equation(s):
// \count~3_combout  = (!count[0] & ((count[2]) # ((count[3]) # (count[1]))))

	.dataa(count[2]),
	.datab(count[3]),
	.datac(count[0]),
	.datad(count[1]),
	.cin(gnd),
	.combout(\count~3_combout ),
	.cout());
// synopsys translate_off
defparam \count~3 .lut_mask = 16'h0F0E;
defparam \count~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N12
cycloneive_lcell_comb \ramaddr~29_wirecell (
// Equation(s):
// \ramaddr~29_wirecell_combout  = !\ramaddr~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\ramaddr~29_combout ),
	.cin(gnd),
	.combout(\ramaddr~29_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~29_wirecell .lut_mask = 16'h00FF;
defparam \ramaddr~29_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: JTAG_X1_Y37_N0
cycloneive_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

// Location: FF_X42_Y34_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y36_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y35_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y35_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y35_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y35_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y35_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y36_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~10 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~13_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~14 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~13 .lut_mask = 16'h5AAF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h33CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .lut_mask = 16'h3C3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .lut_mask = 16'hC30C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h5A5F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .lut_mask = 16'hC3C3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X46_Y34_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y34_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y34_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y34_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y34_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y34_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y34_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y34_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y34_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y34_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .lut_mask = 16'hE4CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .lut_mask = 16'h040C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .lut_mask = 16'hAA00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .lut_mask = 16'hF4A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .lut_mask = 16'hAA00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .lut_mask = 16'hCC50;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .lut_mask = 16'hFAFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .lut_mask = 16'hAAF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .lut_mask = 16'hBB88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .lut_mask = 16'hA001;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .lut_mask = 16'h0010;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .lut_mask = 16'hFFFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y35_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .lut_mask = 16'hC0CA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .lut_mask = 16'hFF01;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .lut_mask = 16'h0004;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y35_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .lut_mask = 16'hDCCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .lut_mask = 16'h1110;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .lut_mask = 16'h5540;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .lut_mask = 16'hF444;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .lut_mask = 16'hDCCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y36_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6 .lut_mask = 16'h14D4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y36_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7 .lut_mask = 16'h0A7A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y36_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 .lut_mask = 16'hDDA4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y36_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9 .lut_mask = 16'h5701;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y36_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .lut_mask = 16'hA13D;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y36_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .lut_mask = 16'h04C8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~5 .lut_mask = 16'h0080;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y36_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12 .lut_mask = 16'h945D;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y36_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 .lut_mask = 16'h7600;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N15
cycloneive_io_ibuf \nRST~input (
	.i(nRST),
	.ibar(gnd),
	.o(\nRST~input_o ));
// synopsys translate_off
defparam \nRST~input .bus_hold = "false";
defparam \nRST~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N8
cycloneive_io_ibuf \syif.tbCTRL~input (
	.i(\syif.tbCTRL ),
	.ibar(gnd),
	.o(\syif.tbCTRL~input_o ));
// synopsys translate_off
defparam \syif.tbCTRL~input .bus_hold = "false";
defparam \syif.tbCTRL~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N1
cycloneive_io_ibuf \syif.addr[1]~input (
	.i(\syif.addr [1]),
	.ibar(gnd),
	.o(\syif.addr[1]~input_o ));
// synopsys translate_off
defparam \syif.addr[1]~input .bus_hold = "false";
defparam \syif.addr[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N8
cycloneive_io_ibuf \syif.addr[0]~input (
	.i(\syif.addr [0]),
	.ibar(gnd),
	.o(\syif.addr[0]~input_o ));
// synopsys translate_off
defparam \syif.addr[0]~input .bus_hold = "false";
defparam \syif.addr[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N15
cycloneive_io_ibuf \syif.addr[3]~input (
	.i(\syif.addr [3]),
	.ibar(gnd),
	.o(\syif.addr[3]~input_o ));
// synopsys translate_off
defparam \syif.addr[3]~input .bus_hold = "false";
defparam \syif.addr[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X56_Y0_N1
cycloneive_io_ibuf \syif.addr[2]~input (
	.i(\syif.addr [2]),
	.ibar(gnd),
	.o(\syif.addr[2]~input_o ));
// synopsys translate_off
defparam \syif.addr[2]~input .bus_hold = "false";
defparam \syif.addr[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y0_N15
cycloneive_io_ibuf \syif.addr[5]~input (
	.i(\syif.addr [5]),
	.ibar(gnd),
	.o(\syif.addr[5]~input_o ));
// synopsys translate_off
defparam \syif.addr[5]~input .bus_hold = "false";
defparam \syif.addr[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N15
cycloneive_io_ibuf \syif.addr[4]~input (
	.i(\syif.addr [4]),
	.ibar(gnd),
	.o(\syif.addr[4]~input_o ));
// synopsys translate_off
defparam \syif.addr[4]~input .bus_hold = "false";
defparam \syif.addr[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N22
cycloneive_io_ibuf \syif.addr[7]~input (
	.i(\syif.addr [7]),
	.ibar(gnd),
	.o(\syif.addr[7]~input_o ));
// synopsys translate_off
defparam \syif.addr[7]~input .bus_hold = "false";
defparam \syif.addr[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y29_N22
cycloneive_io_ibuf \syif.addr[6]~input (
	.i(\syif.addr [6]),
	.ibar(gnd),
	.o(\syif.addr[6]~input_o ));
// synopsys translate_off
defparam \syif.addr[6]~input .bus_hold = "false";
defparam \syif.addr[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N8
cycloneive_io_ibuf \syif.addr[9]~input (
	.i(\syif.addr [9]),
	.ibar(gnd),
	.o(\syif.addr[9]~input_o ));
// synopsys translate_off
defparam \syif.addr[9]~input .bus_hold = "false";
defparam \syif.addr[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y73_N15
cycloneive_io_ibuf \syif.addr[8]~input (
	.i(\syif.addr [8]),
	.ibar(gnd),
	.o(\syif.addr[8]~input_o ));
// synopsys translate_off
defparam \syif.addr[8]~input .bus_hold = "false";
defparam \syif.addr[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y73_N1
cycloneive_io_ibuf \syif.addr[11]~input (
	.i(\syif.addr [11]),
	.ibar(gnd),
	.o(\syif.addr[11]~input_o ));
// synopsys translate_off
defparam \syif.addr[11]~input .bus_hold = "false";
defparam \syif.addr[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X35_Y0_N15
cycloneive_io_ibuf \syif.addr[10]~input (
	.i(\syif.addr [10]),
	.ibar(gnd),
	.o(\syif.addr[10]~input_o ));
// synopsys translate_off
defparam \syif.addr[10]~input .bus_hold = "false";
defparam \syif.addr[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y31_N8
cycloneive_io_ibuf \syif.addr[13]~input (
	.i(\syif.addr [13]),
	.ibar(gnd),
	.o(\syif.addr[13]~input_o ));
// synopsys translate_off
defparam \syif.addr[13]~input .bus_hold = "false";
defparam \syif.addr[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N15
cycloneive_io_ibuf \syif.addr[12]~input (
	.i(\syif.addr [12]),
	.ibar(gnd),
	.o(\syif.addr[12]~input_o ));
// synopsys translate_off
defparam \syif.addr[12]~input .bus_hold = "false";
defparam \syif.addr[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y73_N22
cycloneive_io_ibuf \syif.addr[15]~input (
	.i(\syif.addr [15]),
	.ibar(gnd),
	.o(\syif.addr[15]~input_o ));
// synopsys translate_off
defparam \syif.addr[15]~input .bus_hold = "false";
defparam \syif.addr[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y32_N15
cycloneive_io_ibuf \syif.addr[14]~input (
	.i(\syif.addr [14]),
	.ibar(gnd),
	.o(\syif.addr[14]~input_o ));
// synopsys translate_off
defparam \syif.addr[14]~input .bus_hold = "false";
defparam \syif.addr[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X35_Y0_N22
cycloneive_io_ibuf \syif.addr[17]~input (
	.i(\syif.addr [17]),
	.ibar(gnd),
	.o(\syif.addr[17]~input_o ));
// synopsys translate_off
defparam \syif.addr[17]~input .bus_hold = "false";
defparam \syif.addr[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y0_N22
cycloneive_io_ibuf \syif.addr[16]~input (
	.i(\syif.addr [16]),
	.ibar(gnd),
	.o(\syif.addr[16]~input_o ));
// synopsys translate_off
defparam \syif.addr[16]~input .bus_hold = "false";
defparam \syif.addr[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N8
cycloneive_io_ibuf \syif.addr[19]~input (
	.i(\syif.addr [19]),
	.ibar(gnd),
	.o(\syif.addr[19]~input_o ));
// synopsys translate_off
defparam \syif.addr[19]~input .bus_hold = "false";
defparam \syif.addr[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X47_Y73_N15
cycloneive_io_ibuf \syif.addr[18]~input (
	.i(\syif.addr [18]),
	.ibar(gnd),
	.o(\syif.addr[18]~input_o ));
// synopsys translate_off
defparam \syif.addr[18]~input .bus_hold = "false";
defparam \syif.addr[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N22
cycloneive_io_ibuf \syif.addr[21]~input (
	.i(\syif.addr [21]),
	.ibar(gnd),
	.o(\syif.addr[21]~input_o ));
// synopsys translate_off
defparam \syif.addr[21]~input .bus_hold = "false";
defparam \syif.addr[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X33_Y0_N8
cycloneive_io_ibuf \syif.addr[20]~input (
	.i(\syif.addr [20]),
	.ibar(gnd),
	.o(\syif.addr[20]~input_o ));
// synopsys translate_off
defparam \syif.addr[20]~input .bus_hold = "false";
defparam \syif.addr[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y73_N8
cycloneive_io_ibuf \syif.addr[23]~input (
	.i(\syif.addr [23]),
	.ibar(gnd),
	.o(\syif.addr[23]~input_o ));
// synopsys translate_off
defparam \syif.addr[23]~input .bus_hold = "false";
defparam \syif.addr[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y73_N8
cycloneive_io_ibuf \syif.addr[22]~input (
	.i(\syif.addr [22]),
	.ibar(gnd),
	.o(\syif.addr[22]~input_o ));
// synopsys translate_off
defparam \syif.addr[22]~input .bus_hold = "false";
defparam \syif.addr[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y73_N8
cycloneive_io_ibuf \syif.addr[25]~input (
	.i(\syif.addr [25]),
	.ibar(gnd),
	.o(\syif.addr[25]~input_o ));
// synopsys translate_off
defparam \syif.addr[25]~input .bus_hold = "false";
defparam \syif.addr[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y0_N22
cycloneive_io_ibuf \syif.addr[24]~input (
	.i(\syif.addr [24]),
	.ibar(gnd),
	.o(\syif.addr[24]~input_o ));
// synopsys translate_off
defparam \syif.addr[24]~input .bus_hold = "false";
defparam \syif.addr[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N8
cycloneive_io_ibuf \syif.addr[27]~input (
	.i(\syif.addr [27]),
	.ibar(gnd),
	.o(\syif.addr[27]~input_o ));
// synopsys translate_off
defparam \syif.addr[27]~input .bus_hold = "false";
defparam \syif.addr[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y0_N15
cycloneive_io_ibuf \syif.addr[26]~input (
	.i(\syif.addr [26]),
	.ibar(gnd),
	.o(\syif.addr[26]~input_o ));
// synopsys translate_off
defparam \syif.addr[26]~input .bus_hold = "false";
defparam \syif.addr[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N1
cycloneive_io_ibuf \syif.addr[29]~input (
	.i(\syif.addr [29]),
	.ibar(gnd),
	.o(\syif.addr[29]~input_o ));
// synopsys translate_off
defparam \syif.addr[29]~input .bus_hold = "false";
defparam \syif.addr[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N1
cycloneive_io_ibuf \syif.addr[28]~input (
	.i(\syif.addr [28]),
	.ibar(gnd),
	.o(\syif.addr[28]~input_o ));
// synopsys translate_off
defparam \syif.addr[28]~input .bus_hold = "false";
defparam \syif.addr[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N22
cycloneive_io_ibuf \syif.addr[31]~input (
	.i(\syif.addr [31]),
	.ibar(gnd),
	.o(\syif.addr[31]~input_o ));
// synopsys translate_off
defparam \syif.addr[31]~input .bus_hold = "false";
defparam \syif.addr[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X74_Y0_N15
cycloneive_io_ibuf \syif.addr[30]~input (
	.i(\syif.addr [30]),
	.ibar(gnd),
	.o(\syif.addr[30]~input_o ));
// synopsys translate_off
defparam \syif.addr[30]~input .bus_hold = "false";
defparam \syif.addr[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X56_Y0_N15
cycloneive_io_ibuf \syif.WEN~input (
	.i(\syif.WEN ),
	.ibar(gnd),
	.o(\syif.WEN~input_o ));
// synopsys translate_off
defparam \syif.WEN~input .bus_hold = "false";
defparam \syif.WEN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y28_N8
cycloneive_io_ibuf \syif.REN~input (
	.i(\syif.REN ),
	.ibar(gnd),
	.o(\syif.REN~input_o ));
// synopsys translate_off
defparam \syif.REN~input .bus_hold = "false";
defparam \syif.REN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N8
cycloneive_io_ibuf \CLK~input (
	.i(CLK),
	.ibar(gnd),
	.o(\CLK~input_o ));
// synopsys translate_off
defparam \CLK~input .bus_hold = "false";
defparam \CLK~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N1
cycloneive_io_ibuf \syif.store[0]~input (
	.i(\syif.store [0]),
	.ibar(gnd),
	.o(\syif.store[0]~input_o ));
// synopsys translate_off
defparam \syif.store[0]~input .bus_hold = "false";
defparam \syif.store[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y73_N1
cycloneive_io_ibuf \syif.store[1]~input (
	.i(\syif.store [1]),
	.ibar(gnd),
	.o(\syif.store[1]~input_o ));
// synopsys translate_off
defparam \syif.store[1]~input .bus_hold = "false";
defparam \syif.store[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y30_N8
cycloneive_io_ibuf \syif.store[2]~input (
	.i(\syif.store [2]),
	.ibar(gnd),
	.o(\syif.store[2]~input_o ));
// synopsys translate_off
defparam \syif.store[2]~input .bus_hold = "false";
defparam \syif.store[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y32_N22
cycloneive_io_ibuf \syif.store[3]~input (
	.i(\syif.store [3]),
	.ibar(gnd),
	.o(\syif.store[3]~input_o ));
// synopsys translate_off
defparam \syif.store[3]~input .bus_hold = "false";
defparam \syif.store[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N22
cycloneive_io_ibuf \syif.store[4]~input (
	.i(\syif.store [4]),
	.ibar(gnd),
	.o(\syif.store[4]~input_o ));
// synopsys translate_off
defparam \syif.store[4]~input .bus_hold = "false";
defparam \syif.store[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y0_N15
cycloneive_io_ibuf \syif.store[5]~input (
	.i(\syif.store [5]),
	.ibar(gnd),
	.o(\syif.store[5]~input_o ));
// synopsys translate_off
defparam \syif.store[5]~input .bus_hold = "false";
defparam \syif.store[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y73_N1
cycloneive_io_ibuf \syif.store[6]~input (
	.i(\syif.store [6]),
	.ibar(gnd),
	.o(\syif.store[6]~input_o ));
// synopsys translate_off
defparam \syif.store[6]~input .bus_hold = "false";
defparam \syif.store[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X38_Y0_N1
cycloneive_io_ibuf \syif.store[7]~input (
	.i(\syif.store [7]),
	.ibar(gnd),
	.o(\syif.store[7]~input_o ));
// synopsys translate_off
defparam \syif.store[7]~input .bus_hold = "false";
defparam \syif.store[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N22
cycloneive_io_ibuf \syif.store[8]~input (
	.i(\syif.store [8]),
	.ibar(gnd),
	.o(\syif.store[8]~input_o ));
// synopsys translate_off
defparam \syif.store[8]~input .bus_hold = "false";
defparam \syif.store[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y73_N1
cycloneive_io_ibuf \syif.store[9]~input (
	.i(\syif.store [9]),
	.ibar(gnd),
	.o(\syif.store[9]~input_o ));
// synopsys translate_off
defparam \syif.store[9]~input .bus_hold = "false";
defparam \syif.store[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N1
cycloneive_io_ibuf \syif.store[10]~input (
	.i(\syif.store [10]),
	.ibar(gnd),
	.o(\syif.store[10]~input_o ));
// synopsys translate_off
defparam \syif.store[10]~input .bus_hold = "false";
defparam \syif.store[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y0_N22
cycloneive_io_ibuf \syif.store[11]~input (
	.i(\syif.store [11]),
	.ibar(gnd),
	.o(\syif.store[11]~input_o ));
// synopsys translate_off
defparam \syif.store[11]~input .bus_hold = "false";
defparam \syif.store[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y73_N8
cycloneive_io_ibuf \syif.store[12]~input (
	.i(\syif.store [12]),
	.ibar(gnd),
	.o(\syif.store[12]~input_o ));
// synopsys translate_off
defparam \syif.store[12]~input .bus_hold = "false";
defparam \syif.store[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N8
cycloneive_io_ibuf \syif.store[13]~input (
	.i(\syif.store [13]),
	.ibar(gnd),
	.o(\syif.store[13]~input_o ));
// synopsys translate_off
defparam \syif.store[13]~input .bus_hold = "false";
defparam \syif.store[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X47_Y0_N8
cycloneive_io_ibuf \syif.store[14]~input (
	.i(\syif.store [14]),
	.ibar(gnd),
	.o(\syif.store[14]~input_o ));
// synopsys translate_off
defparam \syif.store[14]~input .bus_hold = "false";
defparam \syif.store[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y29_N15
cycloneive_io_ibuf \syif.store[15]~input (
	.i(\syif.store [15]),
	.ibar(gnd),
	.o(\syif.store[15]~input_o ));
// synopsys translate_off
defparam \syif.store[15]~input .bus_hold = "false";
defparam \syif.store[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N15
cycloneive_io_ibuf \syif.store[16]~input (
	.i(\syif.store [16]),
	.ibar(gnd),
	.o(\syif.store[16]~input_o ));
// synopsys translate_off
defparam \syif.store[16]~input .bus_hold = "false";
defparam \syif.store[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y35_N8
cycloneive_io_ibuf \syif.store[17]~input (
	.i(\syif.store [17]),
	.ibar(gnd),
	.o(\syif.store[17]~input_o ));
// synopsys translate_off
defparam \syif.store[17]~input .bus_hold = "false";
defparam \syif.store[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N8
cycloneive_io_ibuf \syif.store[18]~input (
	.i(\syif.store [18]),
	.ibar(gnd),
	.o(\syif.store[18]~input_o ));
// synopsys translate_off
defparam \syif.store[18]~input .bus_hold = "false";
defparam \syif.store[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N1
cycloneive_io_ibuf \syif.store[19]~input (
	.i(\syif.store [19]),
	.ibar(gnd),
	.o(\syif.store[19]~input_o ));
// synopsys translate_off
defparam \syif.store[19]~input .bus_hold = "false";
defparam \syif.store[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X38_Y73_N15
cycloneive_io_ibuf \syif.store[20]~input (
	.i(\syif.store [20]),
	.ibar(gnd),
	.o(\syif.store[20]~input_o ));
// synopsys translate_off
defparam \syif.store[20]~input .bus_hold = "false";
defparam \syif.store[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N8
cycloneive_io_ibuf \syif.store[21]~input (
	.i(\syif.store [21]),
	.ibar(gnd),
	.o(\syif.store[21]~input_o ));
// synopsys translate_off
defparam \syif.store[21]~input .bus_hold = "false";
defparam \syif.store[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y35_N15
cycloneive_io_ibuf \syif.store[22]~input (
	.i(\syif.store [22]),
	.ibar(gnd),
	.o(\syif.store[22]~input_o ));
// synopsys translate_off
defparam \syif.store[22]~input .bus_hold = "false";
defparam \syif.store[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y30_N1
cycloneive_io_ibuf \syif.store[23]~input (
	.i(\syif.store [23]),
	.ibar(gnd),
	.o(\syif.store[23]~input_o ));
// synopsys translate_off
defparam \syif.store[23]~input .bus_hold = "false";
defparam \syif.store[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N1
cycloneive_io_ibuf \syif.store[24]~input (
	.i(\syif.store [24]),
	.ibar(gnd),
	.o(\syif.store[24]~input_o ));
// synopsys translate_off
defparam \syif.store[24]~input .bus_hold = "false";
defparam \syif.store[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N1
cycloneive_io_ibuf \syif.store[25]~input (
	.i(\syif.store [25]),
	.ibar(gnd),
	.o(\syif.store[25]~input_o ));
// synopsys translate_off
defparam \syif.store[25]~input .bus_hold = "false";
defparam \syif.store[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X47_Y73_N1
cycloneive_io_ibuf \syif.store[26]~input (
	.i(\syif.store [26]),
	.ibar(gnd),
	.o(\syif.store[26]~input_o ));
// synopsys translate_off
defparam \syif.store[26]~input .bus_hold = "false";
defparam \syif.store[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X29_Y0_N15
cycloneive_io_ibuf \syif.store[27]~input (
	.i(\syif.store [27]),
	.ibar(gnd),
	.o(\syif.store[27]~input_o ));
// synopsys translate_off
defparam \syif.store[27]~input .bus_hold = "false";
defparam \syif.store[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y35_N1
cycloneive_io_ibuf \syif.store[28]~input (
	.i(\syif.store [28]),
	.ibar(gnd),
	.o(\syif.store[28]~input_o ));
// synopsys translate_off
defparam \syif.store[28]~input .bus_hold = "false";
defparam \syif.store[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y73_N8
cycloneive_io_ibuf \syif.store[29]~input (
	.i(\syif.store [29]),
	.ibar(gnd),
	.o(\syif.store[29]~input_o ));
// synopsys translate_off
defparam \syif.store[29]~input .bus_hold = "false";
defparam \syif.store[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N15
cycloneive_io_ibuf \syif.store[30]~input (
	.i(\syif.store [30]),
	.ibar(gnd),
	.o(\syif.store[30]~input_o ));
// synopsys translate_off
defparam \syif.store[30]~input .bus_hold = "false";
defparam \syif.store[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N22
cycloneive_io_ibuf \syif.store[31]~input (
	.i(\syif.store [31]),
	.ibar(gnd),
	.o(\syif.store[31]~input_o ));
// synopsys translate_off
defparam \syif.store[31]~input .bus_hold = "false";
defparam \syif.store[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: CLKCTRL_G4
cycloneive_clkctrl \altera_internal_jtag~TCKUTAPclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\altera_internal_jtag~TCKUTAP }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ));
// synopsys translate_off
defparam \altera_internal_jtag~TCKUTAPclkctrl .clock_type = "global clock";
defparam \altera_internal_jtag~TCKUTAPclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G19
cycloneive_clkctrl \CPUCLK~clkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CPUCLK~q }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CPUCLK~clkctrl_outclk ));
// synopsys translate_off
defparam \CPUCLK~clkctrl .clock_type = "global clock";
defparam \CPUCLK~clkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G1
cycloneive_clkctrl \nRST~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\nRST~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\nRST~inputclkctrl_outclk ));
// synopsys translate_off
defparam \nRST~inputclkctrl .clock_type = "global clock";
defparam \nRST~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G2
cycloneive_clkctrl \CLK~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CLK~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CLK~inputclkctrl_outclk ));
// synopsys translate_off
defparam \CLK~inputclkctrl .clock_type = "global clock";
defparam \CLK~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder .lut_mask = 16'hF0F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder .lut_mask = 16'hF0F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .lut_mask = 16'hF0F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOOBUF_X47_Y0_N2
cycloneive_io_obuf \syif.halt~output (
	.i(\CPU|DP|dpif.halt~q ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.halt ),
	.obar());
// synopsys translate_off
defparam \syif.halt~output .bus_hold = "false";
defparam \syif.halt~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N23
cycloneive_io_obuf \syif.load[0]~output (
	.i(\RAM|ramif.ramload[0]~2_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [0]),
	.obar());
// synopsys translate_off
defparam \syif.load[0]~output .bus_hold = "false";
defparam \syif.load[0]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N23
cycloneive_io_obuf \syif.load[1]~output (
	.i(\RAM|ramif.ramload[1]~5_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [1]),
	.obar());
// synopsys translate_off
defparam \syif.load[1]~output .bus_hold = "false";
defparam \syif.load[1]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N23
cycloneive_io_obuf \syif.load[2]~output (
	.i(\RAM|ramif.ramload[2]~6_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [2]),
	.obar());
// synopsys translate_off
defparam \syif.load[2]~output .bus_hold = "false";
defparam \syif.load[2]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y0_N16
cycloneive_io_obuf \syif.load[3]~output (
	.i(\RAM|ramif.ramload[3]~7_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [3]),
	.obar());
// synopsys translate_off
defparam \syif.load[3]~output .bus_hold = "false";
defparam \syif.load[3]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X38_Y0_N9
cycloneive_io_obuf \syif.load[4]~output (
	.i(\RAM|ramif.ramload[4]~8_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [4]),
	.obar());
// synopsys translate_off
defparam \syif.load[4]~output .bus_hold = "false";
defparam \syif.load[4]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N23
cycloneive_io_obuf \syif.load[5]~output (
	.i(\RAM|ramif.ramload[5]~9_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [5]),
	.obar());
// synopsys translate_off
defparam \syif.load[5]~output .bus_hold = "false";
defparam \syif.load[5]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N9
cycloneive_io_obuf \syif.load[6]~output (
	.i(\RAM|ramif.ramload[6]~10_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [6]),
	.obar());
// synopsys translate_off
defparam \syif.load[6]~output .bus_hold = "false";
defparam \syif.load[6]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X58_Y73_N16
cycloneive_io_obuf \syif.load[7]~output (
	.i(\RAM|ramif.ramload[7]~11_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [7]),
	.obar());
// synopsys translate_off
defparam \syif.load[7]~output .bus_hold = "false";
defparam \syif.load[7]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y33_N2
cycloneive_io_obuf \syif.load[8]~output (
	.i(\RAM|ramif.ramload[8]~12_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [8]),
	.obar());
// synopsys translate_off
defparam \syif.load[8]~output .bus_hold = "false";
defparam \syif.load[8]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y28_N23
cycloneive_io_obuf \syif.load[9]~output (
	.i(\RAM|ramif.ramload[9]~13_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [9]),
	.obar());
// synopsys translate_off
defparam \syif.load[9]~output .bus_hold = "false";
defparam \syif.load[9]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y73_N16
cycloneive_io_obuf \syif.load[10]~output (
	.i(\RAM|ramif.ramload[10]~14_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [10]),
	.obar());
// synopsys translate_off
defparam \syif.load[10]~output .bus_hold = "false";
defparam \syif.load[10]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y0_N23
cycloneive_io_obuf \syif.load[11]~output (
	.i(\RAM|ramif.ramload[11]~15_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [11]),
	.obar());
// synopsys translate_off
defparam \syif.load[11]~output .bus_hold = "false";
defparam \syif.load[11]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X67_Y0_N9
cycloneive_io_obuf \syif.load[12]~output (
	.i(\RAM|ramif.ramload[12]~16_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [12]),
	.obar());
// synopsys translate_off
defparam \syif.load[12]~output .bus_hold = "false";
defparam \syif.load[12]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y29_N9
cycloneive_io_obuf \syif.load[13]~output (
	.i(\RAM|ramif.ramload[13]~17_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [13]),
	.obar());
// synopsys translate_off
defparam \syif.load[13]~output .bus_hold = "false";
defparam \syif.load[13]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N16
cycloneive_io_obuf \syif.load[14]~output (
	.i(\RAM|ramif.ramload[14]~18_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [14]),
	.obar());
// synopsys translate_off
defparam \syif.load[14]~output .bus_hold = "false";
defparam \syif.load[14]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N9
cycloneive_io_obuf \syif.load[15]~output (
	.i(\RAM|ramif.ramload[15]~19_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [15]),
	.obar());
// synopsys translate_off
defparam \syif.load[15]~output .bus_hold = "false";
defparam \syif.load[15]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X58_Y73_N2
cycloneive_io_obuf \syif.load[16]~output (
	.i(\RAM|ramif.ramload[16]~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [16]),
	.obar());
// synopsys translate_off
defparam \syif.load[16]~output .bus_hold = "false";
defparam \syif.load[16]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X72_Y0_N9
cycloneive_io_obuf \syif.load[17]~output (
	.i(\RAM|ramif.ramload[17]~21_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [17]),
	.obar());
// synopsys translate_off
defparam \syif.load[17]~output .bus_hold = "false";
defparam \syif.load[17]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N2
cycloneive_io_obuf \syif.load[18]~output (
	.i(\RAM|ramif.ramload[18]~22_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [18]),
	.obar());
// synopsys translate_off
defparam \syif.load[18]~output .bus_hold = "false";
defparam \syif.load[18]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y73_N16
cycloneive_io_obuf \syif.load[19]~output (
	.i(\RAM|ramif.ramload[19]~23_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [19]),
	.obar());
// synopsys translate_off
defparam \syif.load[19]~output .bus_hold = "false";
defparam \syif.load[19]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X72_Y0_N2
cycloneive_io_obuf \syif.load[20]~output (
	.i(\RAM|ramif.ramload[20]~24_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [20]),
	.obar());
// synopsys translate_off
defparam \syif.load[20]~output .bus_hold = "false";
defparam \syif.load[20]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y73_N23
cycloneive_io_obuf \syif.load[21]~output (
	.i(\RAM|ramif.ramload[21]~25_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [21]),
	.obar());
// synopsys translate_off
defparam \syif.load[21]~output .bus_hold = "false";
defparam \syif.load[21]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y73_N23
cycloneive_io_obuf \syif.load[22]~output (
	.i(\RAM|ramif.ramload[22]~26_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [22]),
	.obar());
// synopsys translate_off
defparam \syif.load[22]~output .bus_hold = "false";
defparam \syif.load[22]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N16
cycloneive_io_obuf \syif.load[23]~output (
	.i(\RAM|ramif.ramload[23]~27_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [23]),
	.obar());
// synopsys translate_off
defparam \syif.load[23]~output .bus_hold = "false";
defparam \syif.load[23]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N16
cycloneive_io_obuf \syif.load[24]~output (
	.i(\RAM|ramif.ramload[24]~28_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [24]),
	.obar());
// synopsys translate_off
defparam \syif.load[24]~output .bus_hold = "false";
defparam \syif.load[24]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N9
cycloneive_io_obuf \syif.load[25]~output (
	.i(\RAM|ramif.ramload[25]~29_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [25]),
	.obar());
// synopsys translate_off
defparam \syif.load[25]~output .bus_hold = "false";
defparam \syif.load[25]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X67_Y0_N23
cycloneive_io_obuf \syif.load[26]~output (
	.i(\RAM|ramif.ramload[26]~30_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [26]),
	.obar());
// synopsys translate_off
defparam \syif.load[26]~output .bus_hold = "false";
defparam \syif.load[26]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y28_N16
cycloneive_io_obuf \syif.load[27]~output (
	.i(\RAM|ramif.ramload[27]~31_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [27]),
	.obar());
// synopsys translate_off
defparam \syif.load[27]~output .bus_hold = "false";
defparam \syif.load[27]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N9
cycloneive_io_obuf \syif.load[28]~output (
	.i(\RAM|ramif.ramload[28]~32_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [28]),
	.obar());
// synopsys translate_off
defparam \syif.load[28]~output .bus_hold = "false";
defparam \syif.load[28]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y73_N16
cycloneive_io_obuf \syif.load[29]~output (
	.i(\RAM|ramif.ramload[29]~33_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [29]),
	.obar());
// synopsys translate_off
defparam \syif.load[29]~output .bus_hold = "false";
defparam \syif.load[29]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N2
cycloneive_io_obuf \syif.load[30]~output (
	.i(\RAM|ramif.ramload[30]~34_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [30]),
	.obar());
// synopsys translate_off
defparam \syif.load[30]~output .bus_hold = "false";
defparam \syif.load[30]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X38_Y73_N2
cycloneive_io_obuf \syif.load[31]~output (
	.i(\RAM|ramif.ramload[31]~35_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [31]),
	.obar());
// synopsys translate_off
defparam \syif.load[31]~output .bus_hold = "false";
defparam \syif.load[31]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y37_N1
cycloneive_io_obuf \altera_reserved_tdo~output (
	.i(\altera_internal_jtag~TDO ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(altera_reserved_tdo),
	.obar());
// synopsys translate_off
defparam \altera_reserved_tdo~output .bus_hold = "false";
defparam \altera_reserved_tdo~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOIBUF_X0_Y38_N1
cycloneive_io_ibuf \altera_reserved_tms~input (
	.i(altera_reserved_tms),
	.ibar(gnd),
	.o(\altera_reserved_tms~input_o ));
// synopsys translate_off
defparam \altera_reserved_tms~input .bus_hold = "false";
defparam \altera_reserved_tms~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y39_N1
cycloneive_io_ibuf \altera_reserved_tck~input (
	.i(altera_reserved_tck),
	.ibar(gnd),
	.o(\altera_reserved_tck~input_o ));
// synopsys translate_off
defparam \altera_reserved_tck~input .bus_hold = "false";
defparam \altera_reserved_tck~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y40_N1
cycloneive_io_ibuf \altera_reserved_tdi~input (
	.i(altera_reserved_tdi),
	.ibar(gnd),
	.o(\altera_reserved_tdi~input_o ));
// synopsys translate_off
defparam \altera_reserved_tdi~input .bus_hold = "false";
defparam \altera_reserved_tdi~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .lut_mask = 16'hA0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .lut_mask = 16'hC8C8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .lut_mask = 16'h0C0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y35_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y35_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .lut_mask = 16'h3CF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y35_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .lut_mask = 16'h3373;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .lut_mask = 16'hCCC8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .lut_mask = 16'h5500;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y34_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .lut_mask = 16'hFEFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .lut_mask = 16'hCCF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N4
cycloneive_lcell_comb \~QIC_CREATED_GND~I (
// Equation(s):
// \~QIC_CREATED_GND~I_combout  = GND

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~QIC_CREATED_GND~I_combout ),
	.cout());
// synopsys translate_off
defparam \~QIC_CREATED_GND~I .lut_mask = 16'h0000;
defparam \~QIC_CREATED_GND~I .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .lut_mask = 16'h0808;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~3 .lut_mask = 16'h50D8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y34_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .lut_mask = 16'h3300;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.datac(gnd),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .lut_mask = 16'hEE44;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .lut_mask = 16'hF3C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .lut_mask = 16'hF0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .lut_mask = 16'hFFFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X42_Y35_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .lut_mask = 16'h0001;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .lut_mask = 16'h0F0F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .lut_mask = 16'h0010;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .lut_mask = 16'h0040;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hE0E0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .lut_mask = 16'hA0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y34_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .lut_mask = 16'hCCAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y34_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .lut_mask = 16'hFC30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y34_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .lut_mask = 16'hFC30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y34_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .lut_mask = 16'hF0CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y34_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~4 .lut_mask = 16'h22A4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~4_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~2 .lut_mask = 16'hF078;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y34_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .lut_mask = 16'hAA88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y34_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .lut_mask = 16'hC080;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y34_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~5_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~6 .lut_mask = 16'h22F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y34_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~6_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y34_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .lut_mask = 16'hCC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y34_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y34_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.asdata(\~QIC_CREATED_GND~I_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y35_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .lut_mask = 16'h2A2A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .lut_mask = 16'h4000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y35_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .lut_mask = 16'hFEAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y35_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .lut_mask = 16'hAEAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y35_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .lut_mask = 16'hFCFC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y33_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .lut_mask = 16'hDC98;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(gnd),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .lut_mask = 16'hEE30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .lut_mask = 16'hEE02;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .lut_mask = 16'hF8F8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y36_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~7 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~7_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~8 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~7 .lut_mask = 16'h33CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y36_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~11 .lut_mask = 16'hFFFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y36_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~11_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19 .lut_mask = 16'hF111;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12 .lut_mask = 16'hF888;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y36_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y36_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~8 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~10 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9 .lut_mask = 16'hC303;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X40_Y36_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y36_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~15 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~14 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~15_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~16 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~15 .lut_mask = 16'hC303;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X40_Y36_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y36_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~17 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~16 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~17 .lut_mask = 16'h5A5A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X40_Y36_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~19_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y36_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~4 .lut_mask = 16'h8000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y36_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .lut_mask = 16'h4000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .lut_mask = 16'h00C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y36_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y36_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y36_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y36_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .lut_mask = 16'h0020;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y36_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y36_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y36_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .lut_mask = 16'hCCAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y36_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y36_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~5_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .lut_mask = 16'hEE22;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .lut_mask = 16'h0FFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y35_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .lut_mask = 16'hFC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y35_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y35_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y35_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y35_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .lut_mask = 16'h535B;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y34_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo (
	.clk(!\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y34_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X85_Y47_N0
cycloneive_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y34_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y35_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module pipeline (
	ramiframload_0,
	exmem_ifout_o_1,
	exmem_ifdWEN_o,
	exmem_ifdREN_o,
	pc_1,
	exmem_ifout_o_0,
	pc_0,
	exmem_ifout_o_3,
	pc_3,
	exmem_ifout_o_2,
	pc_2,
	exmem_ifout_o_5,
	pc_5,
	pc_4,
	exmem_ifout_o_4,
	exmem_ifout_o_7,
	pc_7,
	exmem_ifout_o_6,
	pc_6,
	exmem_ifout_o_9,
	pc_9,
	pc_8,
	exmem_ifout_o_8,
	exmem_ifout_o_11,
	pc_11,
	exmem_ifout_o_10,
	pc_10,
	pc_13,
	exmem_ifout_o_13,
	pc_12,
	exmem_ifout_o_12,
	exmem_ifout_o_15,
	pc_15,
	pc_14,
	exmem_ifout_o_14,
	pc_17,
	exmem_ifout_o_17,
	exmem_ifout_o_16,
	pc_16,
	exmem_ifout_o_19,
	pc_19,
	exmem_ifout_o_18,
	pc_18,
	pc_21,
	exmem_ifout_o_21,
	pc_20,
	exmem_ifout_o_20,
	exmem_ifout_o_23,
	pc_23,
	exmem_ifout_o_22,
	pc_22,
	pc_25,
	exmem_ifout_o_25,
	pc_24,
	exmem_ifout_o_24,
	exmem_ifout_o_27,
	pc_27,
	exmem_ifout_o_26,
	pc_26,
	pc_29,
	exmem_ifout_o_29,
	exmem_ifout_o_28,
	pc_28,
	exmem_ifout_o_31,
	pc_31,
	exmem_ifout_o_30,
	pc_30,
	ramiframload_01,
	ramiframload_1,
	ramiframload_11,
	always1,
	always11,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_111,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	exmem_ifrdat2_o_0,
	ramstate,
	exmem_ifrdat2_o_1,
	exmem_ifrdat2_o_2,
	exmem_ifrdat2_o_3,
	exmem_ifrdat2_o_4,
	exmem_ifrdat2_o_5,
	exmem_ifrdat2_o_6,
	exmem_ifrdat2_o_7,
	exmem_ifrdat2_o_8,
	exmem_ifrdat2_o_9,
	exmem_ifrdat2_o_10,
	exmem_ifrdat2_o_11,
	exmem_ifrdat2_o_12,
	exmem_ifrdat2_o_13,
	exmem_ifrdat2_o_14,
	exmem_ifrdat2_o_15,
	exmem_ifrdat2_o_16,
	exmem_ifrdat2_o_17,
	exmem_ifrdat2_o_18,
	exmem_ifrdat2_o_19,
	exmem_ifrdat2_o_20,
	exmem_ifrdat2_o_21,
	exmem_ifrdat2_o_22,
	exmem_ifrdat2_o_23,
	exmem_ifrdat2_o_24,
	exmem_ifrdat2_o_25,
	exmem_ifrdat2_o_26,
	exmem_ifrdat2_o_27,
	exmem_ifrdat2_o_28,
	exmem_ifrdat2_o_29,
	exmem_ifrdat2_o_30,
	exmem_ifrdat2_o_31,
	CLK,
	nRST,
	dpifhalt,
	devpor,
	devclrn,
	devoe);
input 	ramiframload_0;
output 	exmem_ifout_o_1;
output 	exmem_ifdWEN_o;
output 	exmem_ifdREN_o;
output 	pc_1;
output 	exmem_ifout_o_0;
output 	pc_0;
output 	exmem_ifout_o_3;
output 	pc_3;
output 	exmem_ifout_o_2;
output 	pc_2;
output 	exmem_ifout_o_5;
output 	pc_5;
output 	pc_4;
output 	exmem_ifout_o_4;
output 	exmem_ifout_o_7;
output 	pc_7;
output 	exmem_ifout_o_6;
output 	pc_6;
output 	exmem_ifout_o_9;
output 	pc_9;
output 	pc_8;
output 	exmem_ifout_o_8;
output 	exmem_ifout_o_11;
output 	pc_11;
output 	exmem_ifout_o_10;
output 	pc_10;
output 	pc_13;
output 	exmem_ifout_o_13;
output 	pc_12;
output 	exmem_ifout_o_12;
output 	exmem_ifout_o_15;
output 	pc_15;
output 	pc_14;
output 	exmem_ifout_o_14;
output 	pc_17;
output 	exmem_ifout_o_17;
output 	exmem_ifout_o_16;
output 	pc_16;
output 	exmem_ifout_o_19;
output 	pc_19;
output 	exmem_ifout_o_18;
output 	pc_18;
output 	pc_21;
output 	exmem_ifout_o_21;
output 	pc_20;
output 	exmem_ifout_o_20;
output 	exmem_ifout_o_23;
output 	pc_23;
output 	exmem_ifout_o_22;
output 	pc_22;
output 	pc_25;
output 	exmem_ifout_o_25;
output 	pc_24;
output 	exmem_ifout_o_24;
output 	exmem_ifout_o_27;
output 	pc_27;
output 	exmem_ifout_o_26;
output 	pc_26;
output 	pc_29;
output 	exmem_ifout_o_29;
output 	exmem_ifout_o_28;
output 	pc_28;
output 	exmem_ifout_o_31;
output 	pc_31;
output 	exmem_ifout_o_30;
output 	pc_30;
input 	ramiframload_01;
input 	ramiframload_1;
input 	ramiframload_11;
input 	always1;
input 	always11;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_111;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
output 	exmem_ifrdat2_o_0;
input 	ramstate;
output 	exmem_ifrdat2_o_1;
output 	exmem_ifrdat2_o_2;
output 	exmem_ifrdat2_o_3;
output 	exmem_ifrdat2_o_4;
output 	exmem_ifrdat2_o_5;
output 	exmem_ifrdat2_o_6;
output 	exmem_ifrdat2_o_7;
output 	exmem_ifrdat2_o_8;
output 	exmem_ifrdat2_o_9;
output 	exmem_ifrdat2_o_10;
output 	exmem_ifrdat2_o_11;
output 	exmem_ifrdat2_o_12;
output 	exmem_ifrdat2_o_13;
output 	exmem_ifrdat2_o_14;
output 	exmem_ifrdat2_o_15;
output 	exmem_ifrdat2_o_16;
output 	exmem_ifrdat2_o_17;
output 	exmem_ifrdat2_o_18;
output 	exmem_ifrdat2_o_19;
output 	exmem_ifrdat2_o_20;
output 	exmem_ifrdat2_o_21;
output 	exmem_ifrdat2_o_22;
output 	exmem_ifrdat2_o_23;
output 	exmem_ifrdat2_o_24;
output 	exmem_ifrdat2_o_25;
output 	exmem_ifrdat2_o_26;
output 	exmem_ifrdat2_o_27;
output 	exmem_ifrdat2_o_28;
output 	exmem_ifrdat2_o_29;
output 	exmem_ifrdat2_o_30;
output 	exmem_ifrdat2_o_31;
input 	CLK;
input 	nRST;
output 	dpifhalt;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \CC|always1~0_combout ;
wire \CC|always1~1_combout ;


datapath DP(
	.ramiframload_0(ramiframload_0),
	.exmem_ifout_o_1(exmem_ifout_o_1),
	.exmem_ifdWEN_o(exmem_ifdWEN_o),
	.exmem_ifdREN_o(exmem_ifdREN_o),
	.pc_1(pc_1),
	.exmem_ifout_o_0(exmem_ifout_o_0),
	.pc_0(pc_0),
	.exmem_ifout_o_3(exmem_ifout_o_3),
	.pc_3(pc_3),
	.exmem_ifout_o_2(exmem_ifout_o_2),
	.pc_2(pc_2),
	.exmem_ifout_o_5(exmem_ifout_o_5),
	.pc_5(pc_5),
	.pc_4(pc_4),
	.exmem_ifout_o_4(exmem_ifout_o_4),
	.exmem_ifout_o_7(exmem_ifout_o_7),
	.pc_7(pc_7),
	.exmem_ifout_o_6(exmem_ifout_o_6),
	.pc_6(pc_6),
	.exmem_ifout_o_9(exmem_ifout_o_9),
	.pc_9(pc_9),
	.pc_8(pc_8),
	.exmem_ifout_o_8(exmem_ifout_o_8),
	.exmem_ifout_o_11(exmem_ifout_o_11),
	.pc_11(pc_11),
	.exmem_ifout_o_10(exmem_ifout_o_10),
	.pc_10(pc_10),
	.pc_13(pc_13),
	.exmem_ifout_o_13(exmem_ifout_o_13),
	.pc_12(pc_12),
	.exmem_ifout_o_12(exmem_ifout_o_12),
	.exmem_ifout_o_15(exmem_ifout_o_15),
	.pc_15(pc_15),
	.pc_14(pc_14),
	.exmem_ifout_o_14(exmem_ifout_o_14),
	.pc_17(pc_17),
	.exmem_ifout_o_17(exmem_ifout_o_17),
	.exmem_ifout_o_16(exmem_ifout_o_16),
	.pc_16(pc_16),
	.exmem_ifout_o_19(exmem_ifout_o_19),
	.pc_19(pc_19),
	.exmem_ifout_o_18(exmem_ifout_o_18),
	.pc_18(pc_18),
	.pc_21(pc_21),
	.exmem_ifout_o_21(exmem_ifout_o_21),
	.pc_20(pc_20),
	.exmem_ifout_o_20(exmem_ifout_o_20),
	.exmem_ifout_o_23(exmem_ifout_o_23),
	.pc_23(pc_23),
	.exmem_ifout_o_22(exmem_ifout_o_22),
	.pc_22(pc_22),
	.pc_25(pc_25),
	.exmem_ifout_o_25(exmem_ifout_o_25),
	.pc_24(pc_24),
	.exmem_ifout_o_24(exmem_ifout_o_24),
	.exmem_ifout_o_27(exmem_ifout_o_27),
	.pc_27(pc_27),
	.exmem_ifout_o_26(exmem_ifout_o_26),
	.pc_26(pc_26),
	.pc_29(pc_29),
	.exmem_ifout_o_29(exmem_ifout_o_29),
	.exmem_ifout_o_28(exmem_ifout_o_28),
	.pc_28(pc_28),
	.exmem_ifout_o_31(exmem_ifout_o_31),
	.pc_31(pc_31),
	.exmem_ifout_o_30(exmem_ifout_o_30),
	.pc_30(pc_30),
	.ramiframload_01(ramiframload_01),
	.ramiframload_1(ramiframload_1),
	.ramiframload_11(ramiframload_11),
	.always1(always1),
	.always11(always11),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_111(ramiframload_111),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.exmem_ifrdat2_o_0(exmem_ifrdat2_o_0),
	.always12(\CC|always1~0_combout ),
	.ramstate(ramstate),
	.always13(\CC|always1~1_combout ),
	.exmem_ifrdat2_o_1(exmem_ifrdat2_o_1),
	.exmem_ifrdat2_o_2(exmem_ifrdat2_o_2),
	.exmem_ifrdat2_o_3(exmem_ifrdat2_o_3),
	.exmem_ifrdat2_o_4(exmem_ifrdat2_o_4),
	.exmem_ifrdat2_o_5(exmem_ifrdat2_o_5),
	.exmem_ifrdat2_o_6(exmem_ifrdat2_o_6),
	.exmem_ifrdat2_o_7(exmem_ifrdat2_o_7),
	.exmem_ifrdat2_o_8(exmem_ifrdat2_o_8),
	.exmem_ifrdat2_o_9(exmem_ifrdat2_o_9),
	.exmem_ifrdat2_o_10(exmem_ifrdat2_o_10),
	.exmem_ifrdat2_o_11(exmem_ifrdat2_o_11),
	.exmem_ifrdat2_o_12(exmem_ifrdat2_o_12),
	.exmem_ifrdat2_o_13(exmem_ifrdat2_o_13),
	.exmem_ifrdat2_o_14(exmem_ifrdat2_o_14),
	.exmem_ifrdat2_o_15(exmem_ifrdat2_o_15),
	.exmem_ifrdat2_o_16(exmem_ifrdat2_o_16),
	.exmem_ifrdat2_o_17(exmem_ifrdat2_o_17),
	.exmem_ifrdat2_o_18(exmem_ifrdat2_o_18),
	.exmem_ifrdat2_o_19(exmem_ifrdat2_o_19),
	.exmem_ifrdat2_o_20(exmem_ifrdat2_o_20),
	.exmem_ifrdat2_o_21(exmem_ifrdat2_o_21),
	.exmem_ifrdat2_o_22(exmem_ifrdat2_o_22),
	.exmem_ifrdat2_o_23(exmem_ifrdat2_o_23),
	.exmem_ifrdat2_o_24(exmem_ifrdat2_o_24),
	.exmem_ifrdat2_o_25(exmem_ifrdat2_o_25),
	.exmem_ifrdat2_o_26(exmem_ifrdat2_o_26),
	.exmem_ifrdat2_o_27(exmem_ifrdat2_o_27),
	.exmem_ifrdat2_o_28(exmem_ifrdat2_o_28),
	.exmem_ifrdat2_o_29(exmem_ifrdat2_o_29),
	.exmem_ifrdat2_o_30(exmem_ifrdat2_o_30),
	.exmem_ifrdat2_o_31(exmem_ifrdat2_o_31),
	.CLK(CLK),
	.nRST(nRST),
	.dpifhalt(dpifhalt),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

memory_control CC(
	.exmem_ifdWEN_o(exmem_ifdWEN_o),
	.exmem_ifdREN_o(exmem_ifdREN_o),
	.always1(always1),
	.always11(always11),
	.always12(\CC|always1~0_combout ),
	.ramstate(ramstate),
	.always13(\CC|always1~1_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module datapath (
	ramiframload_0,
	exmem_ifout_o_1,
	exmem_ifdWEN_o,
	exmem_ifdREN_o,
	pc_1,
	exmem_ifout_o_0,
	pc_0,
	exmem_ifout_o_3,
	pc_3,
	exmem_ifout_o_2,
	pc_2,
	exmem_ifout_o_5,
	pc_5,
	pc_4,
	exmem_ifout_o_4,
	exmem_ifout_o_7,
	pc_7,
	exmem_ifout_o_6,
	pc_6,
	exmem_ifout_o_9,
	pc_9,
	pc_8,
	exmem_ifout_o_8,
	exmem_ifout_o_11,
	pc_11,
	exmem_ifout_o_10,
	pc_10,
	pc_13,
	exmem_ifout_o_13,
	pc_12,
	exmem_ifout_o_12,
	exmem_ifout_o_15,
	pc_15,
	pc_14,
	exmem_ifout_o_14,
	pc_17,
	exmem_ifout_o_17,
	exmem_ifout_o_16,
	pc_16,
	exmem_ifout_o_19,
	pc_19,
	exmem_ifout_o_18,
	pc_18,
	pc_21,
	exmem_ifout_o_21,
	pc_20,
	exmem_ifout_o_20,
	exmem_ifout_o_23,
	pc_23,
	exmem_ifout_o_22,
	pc_22,
	pc_25,
	exmem_ifout_o_25,
	pc_24,
	exmem_ifout_o_24,
	exmem_ifout_o_27,
	pc_27,
	exmem_ifout_o_26,
	pc_26,
	pc_29,
	exmem_ifout_o_29,
	exmem_ifout_o_28,
	pc_28,
	exmem_ifout_o_31,
	pc_31,
	exmem_ifout_o_30,
	pc_30,
	ramiframload_01,
	ramiframload_1,
	ramiframload_11,
	always1,
	always11,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_111,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	exmem_ifrdat2_o_0,
	always12,
	ramstate,
	always13,
	exmem_ifrdat2_o_1,
	exmem_ifrdat2_o_2,
	exmem_ifrdat2_o_3,
	exmem_ifrdat2_o_4,
	exmem_ifrdat2_o_5,
	exmem_ifrdat2_o_6,
	exmem_ifrdat2_o_7,
	exmem_ifrdat2_o_8,
	exmem_ifrdat2_o_9,
	exmem_ifrdat2_o_10,
	exmem_ifrdat2_o_11,
	exmem_ifrdat2_o_12,
	exmem_ifrdat2_o_13,
	exmem_ifrdat2_o_14,
	exmem_ifrdat2_o_15,
	exmem_ifrdat2_o_16,
	exmem_ifrdat2_o_17,
	exmem_ifrdat2_o_18,
	exmem_ifrdat2_o_19,
	exmem_ifrdat2_o_20,
	exmem_ifrdat2_o_21,
	exmem_ifrdat2_o_22,
	exmem_ifrdat2_o_23,
	exmem_ifrdat2_o_24,
	exmem_ifrdat2_o_25,
	exmem_ifrdat2_o_26,
	exmem_ifrdat2_o_27,
	exmem_ifrdat2_o_28,
	exmem_ifrdat2_o_29,
	exmem_ifrdat2_o_30,
	exmem_ifrdat2_o_31,
	CLK,
	nRST,
	dpifhalt,
	devpor,
	devclrn,
	devoe);
input 	ramiframload_0;
output 	exmem_ifout_o_1;
output 	exmem_ifdWEN_o;
output 	exmem_ifdREN_o;
output 	pc_1;
output 	exmem_ifout_o_0;
output 	pc_0;
output 	exmem_ifout_o_3;
output 	pc_3;
output 	exmem_ifout_o_2;
output 	pc_2;
output 	exmem_ifout_o_5;
output 	pc_5;
output 	pc_4;
output 	exmem_ifout_o_4;
output 	exmem_ifout_o_7;
output 	pc_7;
output 	exmem_ifout_o_6;
output 	pc_6;
output 	exmem_ifout_o_9;
output 	pc_9;
output 	pc_8;
output 	exmem_ifout_o_8;
output 	exmem_ifout_o_11;
output 	pc_11;
output 	exmem_ifout_o_10;
output 	pc_10;
output 	pc_13;
output 	exmem_ifout_o_13;
output 	pc_12;
output 	exmem_ifout_o_12;
output 	exmem_ifout_o_15;
output 	pc_15;
output 	pc_14;
output 	exmem_ifout_o_14;
output 	pc_17;
output 	exmem_ifout_o_17;
output 	exmem_ifout_o_16;
output 	pc_16;
output 	exmem_ifout_o_19;
output 	pc_19;
output 	exmem_ifout_o_18;
output 	pc_18;
output 	pc_21;
output 	exmem_ifout_o_21;
output 	pc_20;
output 	exmem_ifout_o_20;
output 	exmem_ifout_o_23;
output 	pc_23;
output 	exmem_ifout_o_22;
output 	pc_22;
output 	pc_25;
output 	exmem_ifout_o_25;
output 	pc_24;
output 	exmem_ifout_o_24;
output 	exmem_ifout_o_27;
output 	pc_27;
output 	exmem_ifout_o_26;
output 	pc_26;
output 	pc_29;
output 	exmem_ifout_o_29;
output 	exmem_ifout_o_28;
output 	pc_28;
output 	exmem_ifout_o_31;
output 	pc_31;
output 	exmem_ifout_o_30;
output 	pc_30;
input 	ramiframload_01;
input 	ramiframload_1;
input 	ramiframload_11;
input 	always1;
input 	always11;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_111;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
output 	exmem_ifrdat2_o_0;
input 	always12;
input 	ramstate;
input 	always13;
output 	exmem_ifrdat2_o_1;
output 	exmem_ifrdat2_o_2;
output 	exmem_ifrdat2_o_3;
output 	exmem_ifrdat2_o_4;
output 	exmem_ifrdat2_o_5;
output 	exmem_ifrdat2_o_6;
output 	exmem_ifrdat2_o_7;
output 	exmem_ifrdat2_o_8;
output 	exmem_ifrdat2_o_9;
output 	exmem_ifrdat2_o_10;
output 	exmem_ifrdat2_o_11;
output 	exmem_ifrdat2_o_12;
output 	exmem_ifrdat2_o_13;
output 	exmem_ifrdat2_o_14;
output 	exmem_ifrdat2_o_15;
output 	exmem_ifrdat2_o_16;
output 	exmem_ifrdat2_o_17;
output 	exmem_ifrdat2_o_18;
output 	exmem_ifrdat2_o_19;
output 	exmem_ifrdat2_o_20;
output 	exmem_ifrdat2_o_21;
output 	exmem_ifrdat2_o_22;
output 	exmem_ifrdat2_o_23;
output 	exmem_ifrdat2_o_24;
output 	exmem_ifrdat2_o_25;
output 	exmem_ifrdat2_o_26;
output 	exmem_ifrdat2_o_27;
output 	exmem_ifrdat2_o_28;
output 	exmem_ifrdat2_o_29;
output 	exmem_ifrdat2_o_30;
output 	exmem_ifrdat2_o_31;
input 	CLK;
input 	nRST;
output 	dpifhalt;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \nextpc[16]~28_combout ;
wire \nextpc[18]~32_combout ;
wire \nextpc[24]~44_combout ;
wire \nextpc[26]~48_combout ;
wire \nextpc[28]~52_combout ;
wire \EXMEM|exmem_if.halt_o~q ;
wire \rwMEM~0_combout ;
wire \rwMEM~1_combout ;
wire \rwMEM~2_combout ;
wire \rwMEM~3_combout ;
wire \EXMEM|exmem_if.regWEN_o~q ;
wire \rwMEM~4_combout ;
wire \FU|always0~3_combout ;
wire \rwWB~0_combout ;
wire \rwWB~1_combout ;
wire \rwWB~2_combout ;
wire \rwWB~3_combout ;
wire \MEMWB|memwb_if.regWEN_o~q ;
wire \rwWB~4_combout ;
wire \FU|always0~7_combout ;
wire \port_b~0_combout ;
wire \MEMWB|memwb_if.memToReg_o~q ;
wire \MEMWB|memwb_if.jal_o~q ;
wire \wdat~0_combout ;
wire \MEMWB|memwb_if.lui_o~q ;
wire \wdat~1_combout ;
wire \EXMEM|exmem_if.jal_o~q ;
wire \EXMEM|exmem_if.lui_o~q ;
wire \mem_data~0_combout ;
wire \EXMEM|exmem_if.memToReg_o~q ;
wire \mem_data~1_combout ;
wire \mem_data~2_combout ;
wire \mem_data~3_combout ;
wire \mem_data~4_combout ;
wire \FU|fuif.rtReplace[1]~4_combout ;
wire \port_b~1_combout ;
wire \port_b~2_combout ;
wire \port_b~3_combout ;
wire \FU|always0~11_combout ;
wire \FU|always0~15_combout ;
wire \rdat1[1]~0_combout ;
wire \rdat1[1]~1_combout ;
wire \port_b~4_combout ;
wire \port_b~5_combout ;
wire \port_b~6_combout ;
wire \mem_data~5_combout ;
wire \mem_data~6_combout ;
wire \wdat~2_combout ;
wire \wdat~3_combout ;
wire \FU|fuif.rtReplace[0]~5_combout ;
wire \port_b~7_combout ;
wire \rdat1[0]~2_combout ;
wire \rdat1[0]~3_combout ;
wire \wdat~4_combout ;
wire \wdat~5_combout ;
wire \rdat1[2]~4_combout ;
wire \mem_data~7_combout ;
wire \mem_data~8_combout ;
wire \rdat1[2]~5_combout ;
wire \wdat~6_combout ;
wire \wdat~7_combout ;
wire \rdat1[4]~6_combout ;
wire \mem_data~9_combout ;
wire \mem_data~10_combout ;
wire \rdat1[4]~7_combout ;
wire \wdat~8_combout ;
wire \wdat~9_combout ;
wire \rdat1[3]~8_combout ;
wire \mem_data~11_combout ;
wire \mem_data~12_combout ;
wire \rdat1[3]~9_combout ;
wire \port_b~8_combout ;
wire \port_b~9_combout ;
wire \FU|fuif.rtReplace[2]~6_combout ;
wire \port_b~10_combout ;
wire \wdat~10_combout ;
wire \wdat~11_combout ;
wire \rdat1[8]~10_combout ;
wire \mem_data~13_combout ;
wire \mem_data~14_combout ;
wire \rdat1[8]~11_combout ;
wire \wdat~12_combout ;
wire \wdat~13_combout ;
wire \rdat1[7]~12_combout ;
wire \mem_data~15_combout ;
wire \mem_data~16_combout ;
wire \rdat1[7]~13_combout ;
wire \wdat~14_combout ;
wire \wdat~15_combout ;
wire \rdat1[6]~14_combout ;
wire \mem_data~17_combout ;
wire \mem_data~18_combout ;
wire \rdat1[6]~15_combout ;
wire \wdat~16_combout ;
wire \wdat~17_combout ;
wire \rdat1[5]~16_combout ;
wire \mem_data~19_combout ;
wire \mem_data~20_combout ;
wire \rdat1[5]~17_combout ;
wire \port_b~11_combout ;
wire \port_b~12_combout ;
wire \port_b~13_combout ;
wire \FU|fuif.rtReplace[3]~7_combout ;
wire \port_b~14_combout ;
wire \wdat~18_combout ;
wire \wdat~19_combout ;
wire \wdat~20_combout ;
wire \wdat~21_combout ;
wire \rdat1[16]~18_combout ;
wire \mem_data~21_combout ;
wire \mem_data~22_combout ;
wire \mem_data~23_combout ;
wire \mem_data~24_combout ;
wire \rdat1[16]~19_combout ;
wire \wdat~22_combout ;
wire \wdat~23_combout ;
wire \rdat1[15]~20_combout ;
wire \mem_data~25_combout ;
wire \mem_data~26_combout ;
wire \rdat1[15]~21_combout ;
wire \wdat~24_combout ;
wire \wdat~25_combout ;
wire \rdat1[14]~22_combout ;
wire \mem_data~27_combout ;
wire \mem_data~28_combout ;
wire \rdat1[14]~23_combout ;
wire \wdat~26_combout ;
wire \wdat~27_combout ;
wire \rdat1[13]~24_combout ;
wire \mem_data~29_combout ;
wire \mem_data~30_combout ;
wire \rdat1[13]~25_combout ;
wire \wdat~28_combout ;
wire \wdat~29_combout ;
wire \rdat1[12]~26_combout ;
wire \mem_data~31_combout ;
wire \mem_data~32_combout ;
wire \rdat1[12]~27_combout ;
wire \wdat~30_combout ;
wire \wdat~31_combout ;
wire \rdat1[11]~28_combout ;
wire \mem_data~33_combout ;
wire \mem_data~34_combout ;
wire \rdat1[11]~29_combout ;
wire \wdat~32_combout ;
wire \wdat~33_combout ;
wire \rdat1[10]~30_combout ;
wire \mem_data~35_combout ;
wire \mem_data~36_combout ;
wire \rdat1[10]~31_combout ;
wire \wdat~34_combout ;
wire \wdat~35_combout ;
wire \rdat1[9]~32_combout ;
wire \mem_data~37_combout ;
wire \mem_data~38_combout ;
wire \rdat1[9]~33_combout ;
wire \port_b~15_combout ;
wire \port_b~16_combout ;
wire \FU|fuif.rtReplace[4]~8_combout ;
wire \port_b~17_combout ;
wire \wdat~36_combout ;
wire \wdat~37_combout ;
wire \rdat1[31]~34_combout ;
wire \mem_data~39_combout ;
wire \mem_data~40_combout ;
wire \rdat1[31]~35_combout ;
wire \wdat~38_combout ;
wire \wdat~39_combout ;
wire \rdat1[29]~36_combout ;
wire \mem_data~41_combout ;
wire \mem_data~42_combout ;
wire \rdat1[29]~37_combout ;
wire \wdat~40_combout ;
wire \wdat~41_combout ;
wire \rdat1[30]~38_combout ;
wire \mem_data~43_combout ;
wire \mem_data~44_combout ;
wire \rdat1[30]~39_combout ;
wire \wdat~42_combout ;
wire \wdat~43_combout ;
wire \rdat1[28]~40_combout ;
wire \mem_data~45_combout ;
wire \mem_data~46_combout ;
wire \rdat1[28]~41_combout ;
wire \wdat~44_combout ;
wire \wdat~45_combout ;
wire \rdat1[26]~42_combout ;
wire \mem_data~47_combout ;
wire \mem_data~48_combout ;
wire \rdat1[26]~43_combout ;
wire \wdat~46_combout ;
wire \wdat~47_combout ;
wire \rdat1[27]~44_combout ;
wire \mem_data~49_combout ;
wire \mem_data~50_combout ;
wire \rdat1[27]~45_combout ;
wire \wdat~48_combout ;
wire \wdat~49_combout ;
wire \rdat1[25]~46_combout ;
wire \mem_data~51_combout ;
wire \mem_data~52_combout ;
wire \rdat1[25]~47_combout ;
wire \wdat~50_combout ;
wire \wdat~51_combout ;
wire \rdat1[24]~48_combout ;
wire \mem_data~53_combout ;
wire \mem_data~54_combout ;
wire \rdat1[24]~49_combout ;
wire \wdat~52_combout ;
wire \wdat~53_combout ;
wire \rdat1[22]~50_combout ;
wire \mem_data~55_combout ;
wire \mem_data~56_combout ;
wire \rdat1[22]~51_combout ;
wire \wdat~54_combout ;
wire \wdat~55_combout ;
wire \rdat1[23]~52_combout ;
wire \mem_data~57_combout ;
wire \mem_data~58_combout ;
wire \rdat1[23]~53_combout ;
wire \wdat~56_combout ;
wire \wdat~57_combout ;
wire \rdat1[21]~54_combout ;
wire \mem_data~59_combout ;
wire \mem_data~60_combout ;
wire \rdat1[21]~55_combout ;
wire \wdat~58_combout ;
wire \wdat~59_combout ;
wire \rdat1[20]~56_combout ;
wire \mem_data~61_combout ;
wire \mem_data~62_combout ;
wire \rdat1[20]~57_combout ;
wire \wdat~60_combout ;
wire \wdat~61_combout ;
wire \rdat1[18]~58_combout ;
wire \mem_data~63_combout ;
wire \mem_data~64_combout ;
wire \rdat1[18]~59_combout ;
wire \wdat~62_combout ;
wire \wdat~63_combout ;
wire \rdat1[19]~60_combout ;
wire \mem_data~65_combout ;
wire \mem_data~66_combout ;
wire \rdat1[19]~61_combout ;
wire \wdat~64_combout ;
wire \wdat~65_combout ;
wire \rdat1[17]~62_combout ;
wire \mem_data~67_combout ;
wire \mem_data~68_combout ;
wire \rdat1[17]~63_combout ;
wire \port_b~18_combout ;
wire \port_b~19_combout ;
wire \FU|fuif.rtReplace[31]~9_combout ;
wire \port_b~20_combout ;
wire \port_b~21_combout ;
wire \FU|fuif.rtReplace[16]~10_combout ;
wire \port_b~22_combout ;
wire \port_b~23_combout ;
wire \FU|fuif.rtReplace[17]~11_combout ;
wire \port_b~24_combout ;
wire \port_b~25_combout ;
wire \FU|fuif.rtReplace[18]~12_combout ;
wire \port_b~26_combout ;
wire \port_b~27_combout ;
wire \FU|fuif.rtReplace[19]~13_combout ;
wire \port_b~28_combout ;
wire \port_b~29_combout ;
wire \FU|fuif.rtReplace[20]~14_combout ;
wire \port_b~30_combout ;
wire \port_b~31_combout ;
wire \FU|fuif.rtReplace[21]~15_combout ;
wire \port_b~32_combout ;
wire \port_b~33_combout ;
wire \FU|fuif.rtReplace[22]~16_combout ;
wire \port_b~34_combout ;
wire \port_b~35_combout ;
wire \FU|fuif.rtReplace[23]~17_combout ;
wire \port_b~36_combout ;
wire \port_b~37_combout ;
wire \FU|fuif.rtReplace[24]~18_combout ;
wire \port_b~38_combout ;
wire \port_b~39_combout ;
wire \FU|fuif.rtReplace[25]~19_combout ;
wire \port_b~40_combout ;
wire \port_b~41_combout ;
wire \FU|fuif.rtReplace[26]~20_combout ;
wire \port_b~42_combout ;
wire \port_b~43_combout ;
wire \FU|fuif.rtReplace[5]~21_combout ;
wire \port_b~44_combout ;
wire \port_b~45_combout ;
wire \FU|fuif.rtReplace[6]~22_combout ;
wire \port_b~46_combout ;
wire \port_b~47_combout ;
wire \FU|fuif.rtReplace[7]~23_combout ;
wire \port_b~48_combout ;
wire \port_b~49_combout ;
wire \FU|fuif.rtReplace[8]~24_combout ;
wire \port_b~50_combout ;
wire \port_b~51_combout ;
wire \FU|fuif.rtReplace[27]~25_combout ;
wire \port_b~52_combout ;
wire \port_b~53_combout ;
wire \FU|fuif.rtReplace[28]~26_combout ;
wire \port_b~54_combout ;
wire \port_b~55_combout ;
wire \FU|fuif.rtReplace[29]~27_combout ;
wire \port_b~56_combout ;
wire \port_b~57_combout ;
wire \FU|fuif.rtReplace[30]~28_combout ;
wire \port_b~58_combout ;
wire \port_b~59_combout ;
wire \FU|fuif.rtReplace[9]~29_combout ;
wire \port_b~60_combout ;
wire \port_b~61_combout ;
wire \FU|fuif.rtReplace[14]~30_combout ;
wire \port_b~62_combout ;
wire \FU|fuif.rtReplace[15]~31_combout ;
wire \port_b~63_combout ;
wire \port_b~64_combout ;
wire \FU|fuif.rtReplace[10]~32_combout ;
wire \port_b~65_combout ;
wire \port_b~66_combout ;
wire \FU|fuif.rtReplace[11]~33_combout ;
wire \port_b~67_combout ;
wire \port_b~68_combout ;
wire \FU|fuif.rtReplace[12]~34_combout ;
wire \port_b~69_combout ;
wire \FU|fuif.rtReplace[13]~35_combout ;
wire \port_b~70_combout ;
wire \ALU|myif.out[1]~15_combout ;
wire \EXMEM|exmem_if.imm_o[0]~0_combout ;
wire \IDEX|idex_if.dWEN_o~q ;
wire \IDEX|idex_if.dREN_o~q ;
wire \HU|huif.freeze~2_combout ;
wire \IDEX|idex_if.bne_o~q ;
wire \ALU|myif.out[6]~26_combout ;
wire \ALU|myif.out[4]~33_combout ;
wire \port_b~71_combout ;
wire \port_b~72_combout ;
wire \ALU|myif.out[24]~40_combout ;
wire \ALU|myif.out[26]~47_combout ;
wire \ALU|myif.out[25]~54_combout ;
wire \ALU|myif.out[27]~61_combout ;
wire \ALU|myif.out[5]~68_combout ;
wire \ALU|myif.out[7]~81_combout ;
wire \ALU|myif.out[13]~92_combout ;
wire \ALU|myif.out[9]~98_combout ;
wire \ALU|myif.out[8]~104_combout ;
wire \ALU|myif.out[14]~110_combout ;
wire \ALU|myif.out[12]~116_combout ;
wire \ALU|myif.out[15]~122_combout ;
wire \ALU|myif.out[10]~128_combout ;
wire \ALU|myif.out[11]~134_combout ;
wire \ALU|myif.out[23]~152_combout ;
wire \ALU|myif.out[16]~158_combout ;
wire \ALU|myif.out[17]~174_combout ;
wire \ALU|myif.out[18]~180_combout ;
wire \ALU|myif.out[19]~196_combout ;
wire \ALU|myif.out[30]~204_combout ;
wire \ALU|myif.out[21]~220_combout ;
wire \ALU|myif.negative~8_combout ;
wire \ALU|myif.out[22]~226_combout ;
wire \ALU|myif.out[20]~232_combout ;
wire \ALU|myif.out[0]~239_combout ;
wire \ALU|Equal10~10_combout ;
wire \ALU|myif.out[28]~252_combout ;
wire \ALU|myif.out[29]~264_combout ;
wire \ALU|myif.out[2]~274_combout ;
wire \ALU|myif.out[3]~283_combout ;
wire \ALU|myif.out[3]~285_combout ;
wire \ALU|myif.out[2]~289_combout ;
wire \ALU|Equal10~12_combout ;
wire \HU|flush~0_combout ;
wire \IDEX|idex_if.PCSel_o~q ;
wire \HU|huif.flush~0_combout ;
wire \IDEX|idex_if.halt_o~q ;
wire \FU|fuif.rdat2_ow~0_combout ;
wire \CU|always0~0_combout ;
wire \IDEX|idex_if.regWEN_o~q ;
wire \CU|cuif.regWEN~0_combout ;
wire \CU|Equal0~0_combout ;
wire \CU|Equal3~0_combout ;
wire \CU|Equal2~0_combout ;
wire \IDEX|idex_if.jal_o~q ;
wire \IDEX|idex_if.lui_o~q ;
wire \IDEX|idex_if.memToReg_o~q ;
wire \RF|Mux62~9_combout ;
wire \RF|Mux62~19_combout ;
wire \RF|Mux30~9_combout ;
wire \RF|Mux30~19_combout ;
wire \RF|Mux63~9_combout ;
wire \RF|Mux63~19_combout ;
wire \RF|Mux31~9_combout ;
wire \RF|Mux31~19_combout ;
wire \CU|Equal10~0_combout ;
wire \RF|Mux29~9_combout ;
wire \RF|Mux29~19_combout ;
wire \RF|Mux27~9_combout ;
wire \RF|Mux27~19_combout ;
wire \RF|Mux28~9_combout ;
wire \RF|Mux28~19_combout ;
wire \RF|Mux61~9_combout ;
wire \RF|Mux61~19_combout ;
wire \RF|Mux23~9_combout ;
wire \RF|Mux23~19_combout ;
wire \RF|Mux24~9_combout ;
wire \RF|Mux24~19_combout ;
wire \RF|Mux25~9_combout ;
wire \RF|Mux25~19_combout ;
wire \RF|Mux26~9_combout ;
wire \RF|Mux26~19_combout ;
wire \RF|Mux60~9_combout ;
wire \RF|Mux60~19_combout ;
wire \RF|Mux15~9_combout ;
wire \RF|Mux15~19_combout ;
wire \RF|Mux16~9_combout ;
wire \RF|Mux16~19_combout ;
wire \RF|Mux17~9_combout ;
wire \RF|Mux17~19_combout ;
wire \RF|Mux18~9_combout ;
wire \RF|Mux18~19_combout ;
wire \RF|Mux19~9_combout ;
wire \RF|Mux19~19_combout ;
wire \RF|Mux20~9_combout ;
wire \RF|Mux20~19_combout ;
wire \RF|Mux21~9_combout ;
wire \RF|Mux21~19_combout ;
wire \RF|Mux22~9_combout ;
wire \RF|Mux22~19_combout ;
wire \RF|Mux59~9_combout ;
wire \RF|Mux59~19_combout ;
wire \RF|Mux0~9_combout ;
wire \RF|Mux0~19_combout ;
wire \RF|Mux2~9_combout ;
wire \RF|Mux2~19_combout ;
wire \RF|Mux1~9_combout ;
wire \RF|Mux1~19_combout ;
wire \RF|Mux3~9_combout ;
wire \RF|Mux3~19_combout ;
wire \RF|Mux5~9_combout ;
wire \RF|Mux5~19_combout ;
wire \RF|Mux4~9_combout ;
wire \RF|Mux4~19_combout ;
wire \RF|Mux6~9_combout ;
wire \RF|Mux6~19_combout ;
wire \RF|Mux7~9_combout ;
wire \RF|Mux7~19_combout ;
wire \RF|Mux9~9_combout ;
wire \RF|Mux9~19_combout ;
wire \RF|Mux8~9_combout ;
wire \RF|Mux8~19_combout ;
wire \RF|Mux10~9_combout ;
wire \RF|Mux10~19_combout ;
wire \RF|Mux11~9_combout ;
wire \RF|Mux11~19_combout ;
wire \RF|Mux13~9_combout ;
wire \RF|Mux13~19_combout ;
wire \RF|Mux12~9_combout ;
wire \RF|Mux12~19_combout ;
wire \RF|Mux14~9_combout ;
wire \RF|Mux14~19_combout ;
wire \RF|Mux32~9_combout ;
wire \RF|Mux32~19_combout ;
wire \RF|Mux47~9_combout ;
wire \RF|Mux47~19_combout ;
wire \RF|Mux46~9_combout ;
wire \RF|Mux46~19_combout ;
wire \RF|Mux45~9_combout ;
wire \RF|Mux45~19_combout ;
wire \RF|Mux44~9_combout ;
wire \RF|Mux44~19_combout ;
wire \RF|Mux43~9_combout ;
wire \RF|Mux43~19_combout ;
wire \RF|Mux42~9_combout ;
wire \RF|Mux42~19_combout ;
wire \RF|Mux41~9_combout ;
wire \RF|Mux41~19_combout ;
wire \RF|Mux40~9_combout ;
wire \RF|Mux40~19_combout ;
wire \RF|Mux39~9_combout ;
wire \RF|Mux39~19_combout ;
wire \RF|Mux38~9_combout ;
wire \RF|Mux38~19_combout ;
wire \RF|Mux37~9_combout ;
wire \RF|Mux37~19_combout ;
wire \RF|Mux58~9_combout ;
wire \RF|Mux58~19_combout ;
wire \RF|Mux57~9_combout ;
wire \RF|Mux57~19_combout ;
wire \RF|Mux56~9_combout ;
wire \RF|Mux56~19_combout ;
wire \RF|Mux55~9_combout ;
wire \RF|Mux55~19_combout ;
wire \RF|Mux36~9_combout ;
wire \RF|Mux36~19_combout ;
wire \RF|Mux35~9_combout ;
wire \RF|Mux35~19_combout ;
wire \RF|Mux34~9_combout ;
wire \RF|Mux34~19_combout ;
wire \RF|Mux33~9_combout ;
wire \RF|Mux33~19_combout ;
wire \RF|Mux54~9_combout ;
wire \RF|Mux54~19_combout ;
wire \RF|Mux49~9_combout ;
wire \RF|Mux49~19_combout ;
wire \RF|Mux48~9_combout ;
wire \RF|Mux48~19_combout ;
wire \RF|Mux53~9_combout ;
wire \RF|Mux53~19_combout ;
wire \RF|Mux52~9_combout ;
wire \RF|Mux52~19_combout ;
wire \RF|Mux51~9_combout ;
wire \RF|Mux51~19_combout ;
wire \RF|Mux50~9_combout ;
wire \RF|Mux50~19_combout ;
wire \CU|Equal14~0_combout ;
wire \CU|Equal2~1_combout ;
wire \CU|Equal0~1_combout ;
wire \CU|Equal5~0_combout ;
wire \CU|cuif.regWEN~5_combout ;
wire \CU|Equal1~0_combout ;
wire \ALU|myif.out[3]~291_combout ;
wire \new_pc~0_combout ;
wire \pc[1]~feeder_combout ;
wire \always0~0_combout ;
wire \pc[1]~0_combout ;
wire \new_pc~1_combout ;
wire \pc[31]~1_combout ;
wire \Add1~1 ;
wire \Add1~2_combout ;
wire \nextpc[2]~1 ;
wire \nextpc[3]~2_combout ;
wire \pc[31]~2_combout ;
wire \new_pc[3]~2_combout ;
wire \new_pc[3]~3_combout ;
wire \Add1~0_combout ;
wire \nextpc[2]~0_combout ;
wire \new_pc[2]~4_combout ;
wire \new_pc[2]~5_combout ;
wire \nextpc[3]~3 ;
wire \nextpc[4]~5 ;
wire \nextpc[5]~6_combout ;
wire \Add1~3 ;
wire \Add1~5 ;
wire \Add1~6_combout ;
wire \new_pc[5]~6_combout ;
wire \new_pc[5]~7_combout ;
wire \Add1~4_combout ;
wire \nextpc[4]~4_combout ;
wire \new_pc[4]~8_combout ;
wire \new_pc[4]~9_combout ;
wire \Add1~7 ;
wire \Add1~9 ;
wire \Add1~10_combout ;
wire \nextpc[5]~7 ;
wire \nextpc[6]~9 ;
wire \nextpc[7]~10_combout ;
wire \new_pc[7]~10_combout ;
wire \new_pc[7]~11_combout ;
wire \Add1~8_combout ;
wire \nextpc[6]~8_combout ;
wire \new_pc[6]~12_combout ;
wire \new_pc[6]~13_combout ;
wire \nextpc[7]~11 ;
wire \nextpc[8]~13 ;
wire \nextpc[9]~14_combout ;
wire \Add1~11 ;
wire \Add1~13 ;
wire \Add1~14_combout ;
wire \new_pc[9]~14_combout ;
wire \new_pc[9]~15_combout ;
wire \nextpc[8]~12_combout ;
wire \new_pc[8]~16_combout ;
wire \Add1~12_combout ;
wire \new_pc[8]~17_combout ;
wire \nextpc[9]~15 ;
wire \nextpc[10]~17 ;
wire \nextpc[11]~18_combout ;
wire \Add1~15 ;
wire \Add1~17 ;
wire \Add1~18_combout ;
wire \new_pc[11]~18_combout ;
wire \new_pc[11]~19_combout ;
wire \Add1~16_combout ;
wire \nextpc[10]~16_combout ;
wire \new_pc[10]~20_combout ;
wire \new_pc[10]~21_combout ;
wire \Add1~19 ;
wire \Add1~21 ;
wire \Add1~22_combout ;
wire \nextpc[11]~19 ;
wire \nextpc[12]~21 ;
wire \nextpc[13]~22_combout ;
wire \new_pc[13]~22_combout ;
wire \new_pc[13]~23_combout ;
wire \Add1~20_combout ;
wire \nextpc[12]~20_combout ;
wire \new_pc[12]~24_combout ;
wire \new_pc[12]~25_combout ;
wire \nextpc[13]~23 ;
wire \nextpc[14]~25 ;
wire \nextpc[15]~26_combout ;
wire \Add1~23 ;
wire \Add1~25 ;
wire \Add1~26_combout ;
wire \new_pc[15]~26_combout ;
wire \new_pc[15]~27_combout ;
wire \Add1~24_combout ;
wire \nextpc[14]~24_combout ;
wire \new_pc[14]~28_combout ;
wire \new_pc[14]~29_combout ;
wire \Add1~27 ;
wire \Add1~29 ;
wire \Add1~30_combout ;
wire \nextpc[15]~27 ;
wire \nextpc[16]~29 ;
wire \nextpc[17]~30_combout ;
wire \new_pc[17]~30_combout ;
wire \new_pc[17]~31_combout ;
wire \Add1~28_combout ;
wire \new_pc[16]~32_combout ;
wire \new_pc[16]~33_combout ;
wire \Add1~31 ;
wire \Add1~33 ;
wire \Add1~34_combout ;
wire \nextpc[17]~31 ;
wire \nextpc[18]~33 ;
wire \nextpc[19]~34_combout ;
wire \new_pc[19]~34_combout ;
wire \new_pc[19]~35_combout ;
wire \Add1~32_combout ;
wire \new_pc[18]~36_combout ;
wire \new_pc[18]~37_combout ;
wire \Add1~35 ;
wire \Add1~37 ;
wire \Add1~38_combout ;
wire \nextpc[19]~35 ;
wire \nextpc[20]~37 ;
wire \nextpc[21]~38_combout ;
wire \new_pc[21]~38_combout ;
wire \new_pc[21]~39_combout ;
wire \Add1~36_combout ;
wire \nextpc[20]~36_combout ;
wire \new_pc[20]~40_combout ;
wire \new_pc[20]~41_combout ;
wire \Add1~39 ;
wire \Add1~41 ;
wire \Add1~42_combout ;
wire \nextpc[21]~39 ;
wire \nextpc[22]~41 ;
wire \nextpc[23]~42_combout ;
wire \new_pc[23]~42_combout ;
wire \new_pc[23]~43_combout ;
wire \Add1~40_combout ;
wire \nextpc[22]~40_combout ;
wire \new_pc[22]~44_combout ;
wire \new_pc[22]~45_combout ;
wire \nextpc[23]~43 ;
wire \nextpc[24]~45 ;
wire \nextpc[25]~46_combout ;
wire \Add1~43 ;
wire \Add1~45 ;
wire \Add1~46_combout ;
wire \new_pc[25]~46_combout ;
wire \new_pc[25]~47_combout ;
wire \Add1~44_combout ;
wire \new_pc[24]~48_combout ;
wire \new_pc[24]~49_combout ;
wire \nextpc[25]~47 ;
wire \nextpc[26]~49 ;
wire \nextpc[27]~50_combout ;
wire \Add1~47 ;
wire \Add1~49 ;
wire \Add1~50_combout ;
wire \new_pc[27]~50_combout ;
wire \new_pc[27]~51_combout ;
wire \Add1~48_combout ;
wire \new_pc[26]~52_combout ;
wire \new_pc[26]~53_combout ;
wire \Add1~51 ;
wire \Add1~53 ;
wire \Add1~54_combout ;
wire \nextpc[27]~51 ;
wire \nextpc[28]~53 ;
wire \nextpc[29]~54_combout ;
wire \new_pc[29]~54_combout ;
wire \new_pc[29]~55_combout ;
wire \Add1~52_combout ;
wire \new_pc[28]~56_combout ;
wire \new_pc[28]~57_combout ;
wire \nextpc[29]~55 ;
wire \nextpc[30]~57 ;
wire \nextpc[31]~58_combout ;
wire \Add1~55 ;
wire \Add1~57 ;
wire \Add1~58_combout ;
wire \new_pc[31]~58_combout ;
wire \new_pc[31]~59_combout ;
wire \nextpc[30]~56_combout ;
wire \Add1~56_combout ;
wire \new_pc[30]~60_combout ;
wire \new_pc[30]~61_combout ;
wire \dpif.halt~_Duplicate_1_q ;
wire \dpif.halt~0_combout ;
wire [31:0] \IFID|ifid_if.next_pc_o ;
wire [31:0] \IFID|ifid_if.instr_o ;
wire [31:0] \IDEX|idex_if.shamt_o ;
wire [4:0] \IDEX|idex_if.rt_o ;
wire [4:0] \IDEX|idex_if.rs_o ;
wire [31:0] \IDEX|idex_if.rdat2_o ;
wire [31:0] \IDEX|idex_if.rdat1_o ;
wire [4:0] \IDEX|idex_if.rd_o ;
wire [31:0] \IDEX|idex_if.next_pc_o ;
wire [1:0] \IDEX|idex_if.jumpSel_o ;
wire [31:0] \IDEX|idex_if.instr_o ;
wire [15:0] \IDEX|idex_if.imm_o ;
wire [25:0] \IDEX|idex_if.imm_26_o ;
wire [3:0] \IDEX|idex_if.aluop_o ;
wire [1:0] \IDEX|idex_if.RegDest_o ;
wire [1:0] \IDEX|idex_if.ALUSel_o ;
wire [4:0] \EXMEM|exmem_if.rt_o ;
wire [4:0] \EXMEM|exmem_if.rd_o ;
wire [31:0] \EXMEM|exmem_if.next_pc_o ;
wire [15:0] \EXMEM|exmem_if.imm_o ;
wire [1:0] \EXMEM|exmem_if.RegDest_o ;
wire [4:0] \MEMWB|memwb_if.rt_o ;
wire [4:0] \MEMWB|memwb_if.rd_o ;
wire [31:0] \MEMWB|memwb_if.out_o ;
wire [31:0] \MEMWB|memwb_if.next_pc_o ;
wire [15:0] \MEMWB|memwb_if.imm_o ;
wire [31:0] \MEMWB|memwb_if.dmemload_o ;
wire [1:0] \MEMWB|memwb_if.RegDest_o ;


hazard_unit HU(
	.exmem_ifdWEN_o(exmem_ifdWEN_o),
	.exmem_ifdREN_o(exmem_ifdREN_o),
	.rwMEM(\rwMEM~0_combout ),
	.rwMEM1(\rwMEM~1_combout ),
	.rwMEM2(\rwMEM~2_combout ),
	.rwMEM3(\rwMEM~3_combout ),
	.exmem_ifregWEN_o(\EXMEM|exmem_if.regWEN_o~q ),
	.rwMEM4(\rwMEM~4_combout ),
	.myifout_1(\ALU|myif.out[1]~15_combout ),
	.idex_ifjumpSel_o_1(\IDEX|idex_if.jumpSel_o [1]),
	.idex_ifjumpSel_o_0(\IDEX|idex_if.jumpSel_o [0]),
	.idex_ifinstr_o_31(\IDEX|idex_if.instr_o [31]),
	.idex_ifinstr_o_30(\IDEX|idex_if.instr_o [30]),
	.idex_ifinstr_o_27(\IDEX|idex_if.instr_o [27]),
	.idex_ifinstr_o_26(\IDEX|idex_if.instr_o [26]),
	.idex_ifinstr_o_28(\IDEX|idex_if.instr_o [28]),
	.ifid_ifinstr_o_17(\IFID|ifid_if.instr_o [17]),
	.ifid_ifinstr_o_16(\IFID|ifid_if.instr_o [16]),
	.ifid_ifinstr_o_19(\IFID|ifid_if.instr_o [19]),
	.ifid_ifinstr_o_18(\IFID|ifid_if.instr_o [18]),
	.ifid_ifinstr_o_20(\IFID|ifid_if.instr_o [20]),
	.ifid_ifinstr_o_22(\IFID|ifid_if.instr_o [22]),
	.ifid_ifinstr_o_21(\IFID|ifid_if.instr_o [21]),
	.ifid_ifinstr_o_24(\IFID|ifid_if.instr_o [24]),
	.ifid_ifinstr_o_23(\IFID|ifid_if.instr_o [23]),
	.ifid_ifinstr_o_25(\IFID|ifid_if.instr_o [25]),
	.huiffreeze(\HU|huif.freeze~2_combout ),
	.idex_ifbne_o(\IDEX|idex_if.bne_o~q ),
	.Equal10(\ALU|Equal10~10_combout ),
	.Equal101(\ALU|Equal10~12_combout ),
	.flush(\HU|flush~0_combout ),
	.idex_ifPCSel_o(\IDEX|idex_if.PCSel_o~q ),
	.huifflush(\HU|huif.flush~0_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

mem_wb MEMWB(
	.exmem_ifout_o_1(exmem_ifout_o_1),
	.exmem_ifout_o_0(exmem_ifout_o_0),
	.exmem_ifout_o_3(exmem_ifout_o_3),
	.exmem_ifout_o_2(exmem_ifout_o_2),
	.exmem_ifout_o_5(exmem_ifout_o_5),
	.exmem_ifout_o_4(exmem_ifout_o_4),
	.exmem_ifout_o_7(exmem_ifout_o_7),
	.exmem_ifout_o_6(exmem_ifout_o_6),
	.exmem_ifout_o_9(exmem_ifout_o_9),
	.exmem_ifout_o_8(exmem_ifout_o_8),
	.exmem_ifout_o_11(exmem_ifout_o_11),
	.exmem_ifout_o_10(exmem_ifout_o_10),
	.exmem_ifout_o_13(exmem_ifout_o_13),
	.exmem_ifout_o_12(exmem_ifout_o_12),
	.exmem_ifout_o_15(exmem_ifout_o_15),
	.exmem_ifout_o_14(exmem_ifout_o_14),
	.exmem_ifout_o_17(exmem_ifout_o_17),
	.exmem_ifout_o_16(exmem_ifout_o_16),
	.exmem_ifout_o_19(exmem_ifout_o_19),
	.exmem_ifout_o_18(exmem_ifout_o_18),
	.exmem_ifout_o_21(exmem_ifout_o_21),
	.exmem_ifout_o_20(exmem_ifout_o_20),
	.exmem_ifout_o_23(exmem_ifout_o_23),
	.exmem_ifout_o_22(exmem_ifout_o_22),
	.exmem_ifout_o_25(exmem_ifout_o_25),
	.exmem_ifout_o_24(exmem_ifout_o_24),
	.exmem_ifout_o_27(exmem_ifout_o_27),
	.exmem_ifout_o_26(exmem_ifout_o_26),
	.exmem_ifout_o_29(exmem_ifout_o_29),
	.exmem_ifout_o_28(exmem_ifout_o_28),
	.exmem_ifout_o_31(exmem_ifout_o_31),
	.exmem_ifout_o_30(exmem_ifout_o_30),
	.ramiframload_0(ramiframload_01),
	.ramiframload_1(ramiframload_11),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_111),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.exmem_ifRegDest_o_1(\EXMEM|exmem_if.RegDest_o [1]),
	.exmem_ifrt_o_1(\EXMEM|exmem_if.rt_o [1]),
	.exmem_ifrd_o_1(\EXMEM|exmem_if.rd_o [1]),
	.exmem_ifRegDest_o_0(\EXMEM|exmem_if.RegDest_o [0]),
	.exmem_ifrt_o_0(\EXMEM|exmem_if.rt_o [0]),
	.exmem_ifrd_o_0(\EXMEM|exmem_if.rd_o [0]),
	.exmem_ifrt_o_3(\EXMEM|exmem_if.rt_o [3]),
	.exmem_ifrd_o_3(\EXMEM|exmem_if.rd_o [3]),
	.exmem_ifrt_o_2(\EXMEM|exmem_if.rt_o [2]),
	.exmem_ifrd_o_2(\EXMEM|exmem_if.rd_o [2]),
	.exmem_ifregWEN_o(\EXMEM|exmem_if.regWEN_o~q ),
	.exmem_ifrt_o_4(\EXMEM|exmem_if.rt_o [4]),
	.exmem_ifrd_o_4(\EXMEM|exmem_if.rd_o [4]),
	.memwb_ifRegDest_o_1(\MEMWB|memwb_if.RegDest_o [1]),
	.memwb_ifrt_o_1(\MEMWB|memwb_if.rt_o [1]),
	.memwb_ifrd_o_1(\MEMWB|memwb_if.rd_o [1]),
	.memwb_ifRegDest_o_0(\MEMWB|memwb_if.RegDest_o [0]),
	.memwb_ifrt_o_0(\MEMWB|memwb_if.rt_o [0]),
	.memwb_ifrd_o_0(\MEMWB|memwb_if.rd_o [0]),
	.memwb_ifrt_o_3(\MEMWB|memwb_if.rt_o [3]),
	.memwb_ifrd_o_3(\MEMWB|memwb_if.rd_o [3]),
	.memwb_ifrt_o_2(\MEMWB|memwb_if.rt_o [2]),
	.memwb_ifrd_o_2(\MEMWB|memwb_if.rd_o [2]),
	.memwb_ifregWEN_o(\MEMWB|memwb_if.regWEN_o~q ),
	.memwb_ifrt_o_4(\MEMWB|memwb_if.rt_o [4]),
	.memwb_ifrd_o_4(\MEMWB|memwb_if.rd_o [4]),
	.memwb_ifdmemload_o_1(\MEMWB|memwb_if.dmemload_o [1]),
	.memwb_ifout_o_1(\MEMWB|memwb_if.out_o [1]),
	.memwb_ifmemToReg_o(\MEMWB|memwb_if.memToReg_o~q ),
	.memwb_ifjal_o(\MEMWB|memwb_if.jal_o~q ),
	.memwb_ifnext_pc_o_1(\MEMWB|memwb_if.next_pc_o [1]),
	.memwb_iflui_o(\MEMWB|memwb_if.lui_o~q ),
	.exmem_ifjal_o(\EXMEM|exmem_if.jal_o~q ),
	.exmem_iflui_o(\EXMEM|exmem_if.lui_o~q ),
	.exmem_ifnext_pc_o_1(\EXMEM|exmem_if.next_pc_o [1]),
	.exmem_ifmemToReg_o(\EXMEM|exmem_if.memToReg_o~q ),
	.exmem_ifnext_pc_o_0(\EXMEM|exmem_if.next_pc_o [0]),
	.memwb_ifdmemload_o_0(\MEMWB|memwb_if.dmemload_o [0]),
	.memwb_ifout_o_0(\MEMWB|memwb_if.out_o [0]),
	.memwb_ifnext_pc_o_0(\MEMWB|memwb_if.next_pc_o [0]),
	.memwb_ifdmemload_o_2(\MEMWB|memwb_if.dmemload_o [2]),
	.memwb_ifout_o_2(\MEMWB|memwb_if.out_o [2]),
	.memwb_ifnext_pc_o_2(\MEMWB|memwb_if.next_pc_o [2]),
	.exmem_ifnext_pc_o_2(\EXMEM|exmem_if.next_pc_o [2]),
	.memwb_ifdmemload_o_4(\MEMWB|memwb_if.dmemload_o [4]),
	.memwb_ifout_o_4(\MEMWB|memwb_if.out_o [4]),
	.memwb_ifnext_pc_o_4(\MEMWB|memwb_if.next_pc_o [4]),
	.exmem_ifnext_pc_o_4(\EXMEM|exmem_if.next_pc_o [4]),
	.memwb_ifdmemload_o_3(\MEMWB|memwb_if.dmemload_o [3]),
	.memwb_ifout_o_3(\MEMWB|memwb_if.out_o [3]),
	.memwb_ifnext_pc_o_3(\MEMWB|memwb_if.next_pc_o [3]),
	.exmem_ifnext_pc_o_3(\EXMEM|exmem_if.next_pc_o [3]),
	.memwb_ifdmemload_o_8(\MEMWB|memwb_if.dmemload_o [8]),
	.memwb_ifout_o_8(\MEMWB|memwb_if.out_o [8]),
	.memwb_ifnext_pc_o_8(\MEMWB|memwb_if.next_pc_o [8]),
	.exmem_ifnext_pc_o_8(\EXMEM|exmem_if.next_pc_o [8]),
	.memwb_ifdmemload_o_7(\MEMWB|memwb_if.dmemload_o [7]),
	.memwb_ifout_o_7(\MEMWB|memwb_if.out_o [7]),
	.memwb_ifnext_pc_o_7(\MEMWB|memwb_if.next_pc_o [7]),
	.exmem_ifnext_pc_o_7(\EXMEM|exmem_if.next_pc_o [7]),
	.memwb_ifdmemload_o_6(\MEMWB|memwb_if.dmemload_o [6]),
	.memwb_ifout_o_6(\MEMWB|memwb_if.out_o [6]),
	.memwb_ifnext_pc_o_6(\MEMWB|memwb_if.next_pc_o [6]),
	.exmem_ifnext_pc_o_6(\EXMEM|exmem_if.next_pc_o [6]),
	.memwb_ifdmemload_o_5(\MEMWB|memwb_if.dmemload_o [5]),
	.memwb_ifout_o_5(\MEMWB|memwb_if.out_o [5]),
	.memwb_ifnext_pc_o_5(\MEMWB|memwb_if.next_pc_o [5]),
	.exmem_ifnext_pc_o_5(\EXMEM|exmem_if.next_pc_o [5]),
	.memwb_ifdmemload_o_16(\MEMWB|memwb_if.dmemload_o [16]),
	.memwb_ifnext_pc_o_16(\MEMWB|memwb_if.next_pc_o [16]),
	.memwb_ifout_o_16(\MEMWB|memwb_if.out_o [16]),
	.memwb_ifimm_o_0(\MEMWB|memwb_if.imm_o [0]),
	.exmem_ifimm_o_0(\EXMEM|exmem_if.imm_o [0]),
	.exmem_ifnext_pc_o_16(\EXMEM|exmem_if.next_pc_o [16]),
	.memwb_ifdmemload_o_15(\MEMWB|memwb_if.dmemload_o [15]),
	.memwb_ifout_o_15(\MEMWB|memwb_if.out_o [15]),
	.memwb_ifnext_pc_o_15(\MEMWB|memwb_if.next_pc_o [15]),
	.exmem_ifnext_pc_o_15(\EXMEM|exmem_if.next_pc_o [15]),
	.memwb_ifdmemload_o_14(\MEMWB|memwb_if.dmemload_o [14]),
	.memwb_ifout_o_14(\MEMWB|memwb_if.out_o [14]),
	.memwb_ifnext_pc_o_14(\MEMWB|memwb_if.next_pc_o [14]),
	.exmem_ifnext_pc_o_14(\EXMEM|exmem_if.next_pc_o [14]),
	.memwb_ifdmemload_o_13(\MEMWB|memwb_if.dmemload_o [13]),
	.memwb_ifout_o_13(\MEMWB|memwb_if.out_o [13]),
	.memwb_ifnext_pc_o_13(\MEMWB|memwb_if.next_pc_o [13]),
	.exmem_ifnext_pc_o_13(\EXMEM|exmem_if.next_pc_o [13]),
	.memwb_ifdmemload_o_12(\MEMWB|memwb_if.dmemload_o [12]),
	.memwb_ifout_o_12(\MEMWB|memwb_if.out_o [12]),
	.memwb_ifnext_pc_o_12(\MEMWB|memwb_if.next_pc_o [12]),
	.exmem_ifnext_pc_o_12(\EXMEM|exmem_if.next_pc_o [12]),
	.memwb_ifdmemload_o_11(\MEMWB|memwb_if.dmemload_o [11]),
	.memwb_ifout_o_11(\MEMWB|memwb_if.out_o [11]),
	.memwb_ifnext_pc_o_11(\MEMWB|memwb_if.next_pc_o [11]),
	.exmem_ifnext_pc_o_11(\EXMEM|exmem_if.next_pc_o [11]),
	.memwb_ifdmemload_o_10(\MEMWB|memwb_if.dmemload_o [10]),
	.memwb_ifout_o_10(\MEMWB|memwb_if.out_o [10]),
	.memwb_ifnext_pc_o_10(\MEMWB|memwb_if.next_pc_o [10]),
	.exmem_ifnext_pc_o_10(\EXMEM|exmem_if.next_pc_o [10]),
	.memwb_ifdmemload_o_9(\MEMWB|memwb_if.dmemload_o [9]),
	.memwb_ifout_o_9(\MEMWB|memwb_if.out_o [9]),
	.memwb_ifnext_pc_o_9(\MEMWB|memwb_if.next_pc_o [9]),
	.exmem_ifnext_pc_o_9(\EXMEM|exmem_if.next_pc_o [9]),
	.memwb_ifnext_pc_o_31(\MEMWB|memwb_if.next_pc_o [31]),
	.memwb_ifdmemload_o_31(\MEMWB|memwb_if.dmemload_o [31]),
	.memwb_ifout_o_31(\MEMWB|memwb_if.out_o [31]),
	.memwb_ifimm_o_15(\MEMWB|memwb_if.imm_o [15]),
	.exmem_ifnext_pc_o_31(\EXMEM|exmem_if.next_pc_o [31]),
	.exmem_ifimm_o_15(\EXMEM|exmem_if.imm_o [15]),
	.memwb_ifnext_pc_o_29(\MEMWB|memwb_if.next_pc_o [29]),
	.memwb_ifdmemload_o_29(\MEMWB|memwb_if.dmemload_o [29]),
	.memwb_ifout_o_29(\MEMWB|memwb_if.out_o [29]),
	.memwb_ifimm_o_13(\MEMWB|memwb_if.imm_o [13]),
	.exmem_ifnext_pc_o_29(\EXMEM|exmem_if.next_pc_o [29]),
	.exmem_ifimm_o_13(\EXMEM|exmem_if.imm_o [13]),
	.memwb_ifdmemload_o_30(\MEMWB|memwb_if.dmemload_o [30]),
	.memwb_ifnext_pc_o_30(\MEMWB|memwb_if.next_pc_o [30]),
	.memwb_ifout_o_30(\MEMWB|memwb_if.out_o [30]),
	.memwb_ifimm_o_14(\MEMWB|memwb_if.imm_o [14]),
	.exmem_ifimm_o_14(\EXMEM|exmem_if.imm_o [14]),
	.exmem_ifnext_pc_o_30(\EXMEM|exmem_if.next_pc_o [30]),
	.memwb_ifdmemload_o_28(\MEMWB|memwb_if.dmemload_o [28]),
	.memwb_ifnext_pc_o_28(\MEMWB|memwb_if.next_pc_o [28]),
	.memwb_ifout_o_28(\MEMWB|memwb_if.out_o [28]),
	.memwb_ifimm_o_12(\MEMWB|memwb_if.imm_o [12]),
	.exmem_ifimm_o_12(\EXMEM|exmem_if.imm_o [12]),
	.exmem_ifnext_pc_o_28(\EXMEM|exmem_if.next_pc_o [28]),
	.memwb_ifdmemload_o_26(\MEMWB|memwb_if.dmemload_o [26]),
	.memwb_ifnext_pc_o_26(\MEMWB|memwb_if.next_pc_o [26]),
	.memwb_ifout_o_26(\MEMWB|memwb_if.out_o [26]),
	.memwb_ifimm_o_10(\MEMWB|memwb_if.imm_o [10]),
	.exmem_ifimm_o_10(\EXMEM|exmem_if.imm_o [10]),
	.exmem_ifnext_pc_o_26(\EXMEM|exmem_if.next_pc_o [26]),
	.memwb_ifnext_pc_o_27(\MEMWB|memwb_if.next_pc_o [27]),
	.memwb_ifdmemload_o_27(\MEMWB|memwb_if.dmemload_o [27]),
	.memwb_ifout_o_27(\MEMWB|memwb_if.out_o [27]),
	.memwb_ifimm_o_11(\MEMWB|memwb_if.imm_o [11]),
	.exmem_ifnext_pc_o_27(\EXMEM|exmem_if.next_pc_o [27]),
	.exmem_ifimm_o_11(\EXMEM|exmem_if.imm_o [11]),
	.memwb_ifnext_pc_o_25(\MEMWB|memwb_if.next_pc_o [25]),
	.memwb_ifdmemload_o_25(\MEMWB|memwb_if.dmemload_o [25]),
	.memwb_ifout_o_25(\MEMWB|memwb_if.out_o [25]),
	.memwb_ifimm_o_9(\MEMWB|memwb_if.imm_o [9]),
	.exmem_ifnext_pc_o_25(\EXMEM|exmem_if.next_pc_o [25]),
	.exmem_ifimm_o_9(\EXMEM|exmem_if.imm_o [9]),
	.memwb_ifdmemload_o_24(\MEMWB|memwb_if.dmemload_o [24]),
	.memwb_ifnext_pc_o_24(\MEMWB|memwb_if.next_pc_o [24]),
	.memwb_ifout_o_24(\MEMWB|memwb_if.out_o [24]),
	.memwb_ifimm_o_8(\MEMWB|memwb_if.imm_o [8]),
	.exmem_ifimm_o_8(\EXMEM|exmem_if.imm_o [8]),
	.exmem_ifnext_pc_o_24(\EXMEM|exmem_if.next_pc_o [24]),
	.memwb_ifdmemload_o_22(\MEMWB|memwb_if.dmemload_o [22]),
	.memwb_ifnext_pc_o_22(\MEMWB|memwb_if.next_pc_o [22]),
	.memwb_ifout_o_22(\MEMWB|memwb_if.out_o [22]),
	.memwb_ifimm_o_6(\MEMWB|memwb_if.imm_o [6]),
	.exmem_ifimm_o_6(\EXMEM|exmem_if.imm_o [6]),
	.exmem_ifnext_pc_o_22(\EXMEM|exmem_if.next_pc_o [22]),
	.memwb_ifnext_pc_o_23(\MEMWB|memwb_if.next_pc_o [23]),
	.memwb_ifdmemload_o_23(\MEMWB|memwb_if.dmemload_o [23]),
	.memwb_ifout_o_23(\MEMWB|memwb_if.out_o [23]),
	.memwb_ifimm_o_7(\MEMWB|memwb_if.imm_o [7]),
	.exmem_ifnext_pc_o_23(\EXMEM|exmem_if.next_pc_o [23]),
	.exmem_ifimm_o_7(\EXMEM|exmem_if.imm_o [7]),
	.memwb_ifnext_pc_o_21(\MEMWB|memwb_if.next_pc_o [21]),
	.memwb_ifdmemload_o_21(\MEMWB|memwb_if.dmemload_o [21]),
	.memwb_ifout_o_21(\MEMWB|memwb_if.out_o [21]),
	.memwb_ifimm_o_5(\MEMWB|memwb_if.imm_o [5]),
	.exmem_ifnext_pc_o_21(\EXMEM|exmem_if.next_pc_o [21]),
	.exmem_ifimm_o_5(\EXMEM|exmem_if.imm_o [5]),
	.memwb_ifdmemload_o_20(\MEMWB|memwb_if.dmemload_o [20]),
	.memwb_ifnext_pc_o_20(\MEMWB|memwb_if.next_pc_o [20]),
	.memwb_ifout_o_20(\MEMWB|memwb_if.out_o [20]),
	.memwb_ifimm_o_4(\MEMWB|memwb_if.imm_o [4]),
	.exmem_ifimm_o_4(\EXMEM|exmem_if.imm_o [4]),
	.exmem_ifnext_pc_o_20(\EXMEM|exmem_if.next_pc_o [20]),
	.memwb_ifdmemload_o_18(\MEMWB|memwb_if.dmemload_o [18]),
	.memwb_ifnext_pc_o_18(\MEMWB|memwb_if.next_pc_o [18]),
	.memwb_ifout_o_18(\MEMWB|memwb_if.out_o [18]),
	.memwb_ifimm_o_2(\MEMWB|memwb_if.imm_o [2]),
	.exmem_ifimm_o_2(\EXMEM|exmem_if.imm_o [2]),
	.exmem_ifnext_pc_o_18(\EXMEM|exmem_if.next_pc_o [18]),
	.memwb_ifnext_pc_o_19(\MEMWB|memwb_if.next_pc_o [19]),
	.memwb_ifdmemload_o_19(\MEMWB|memwb_if.dmemload_o [19]),
	.memwb_ifout_o_19(\MEMWB|memwb_if.out_o [19]),
	.memwb_ifimm_o_3(\MEMWB|memwb_if.imm_o [3]),
	.exmem_ifnext_pc_o_19(\EXMEM|exmem_if.next_pc_o [19]),
	.exmem_ifimm_o_3(\EXMEM|exmem_if.imm_o [3]),
	.memwb_ifnext_pc_o_17(\MEMWB|memwb_if.next_pc_o [17]),
	.memwb_ifdmemload_o_17(\MEMWB|memwb_if.dmemload_o [17]),
	.memwb_ifout_o_17(\MEMWB|memwb_if.out_o [17]),
	.memwb_ifimm_o_1(\MEMWB|memwb_if.imm_o [1]),
	.exmem_ifnext_pc_o_17(\EXMEM|exmem_if.next_pc_o [17]),
	.exmem_ifimm_o_1(\EXMEM|exmem_if.imm_o [1]),
	.exmem_ifimm_o_01(\EXMEM|exmem_if.imm_o[0]~0_combout ),
	.CPUCLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

ex_mem EXMEM(
	.exmem_ifout_o_1(exmem_ifout_o_1),
	.exmem_ifdWEN_o(exmem_ifdWEN_o),
	.exmem_ifdREN_o(exmem_ifdREN_o),
	.exmem_ifout_o_0(exmem_ifout_o_0),
	.exmem_ifout_o_3(exmem_ifout_o_3),
	.exmem_ifout_o_2(exmem_ifout_o_2),
	.exmem_ifout_o_5(exmem_ifout_o_5),
	.exmem_ifout_o_4(exmem_ifout_o_4),
	.exmem_ifout_o_7(exmem_ifout_o_7),
	.exmem_ifout_o_6(exmem_ifout_o_6),
	.exmem_ifout_o_9(exmem_ifout_o_9),
	.exmem_ifout_o_8(exmem_ifout_o_8),
	.exmem_ifout_o_11(exmem_ifout_o_11),
	.exmem_ifout_o_10(exmem_ifout_o_10),
	.exmem_ifout_o_13(exmem_ifout_o_13),
	.exmem_ifout_o_12(exmem_ifout_o_12),
	.exmem_ifout_o_15(exmem_ifout_o_15),
	.exmem_ifout_o_14(exmem_ifout_o_14),
	.exmem_ifout_o_17(exmem_ifout_o_17),
	.exmem_ifout_o_16(exmem_ifout_o_16),
	.exmem_ifout_o_19(exmem_ifout_o_19),
	.exmem_ifout_o_18(exmem_ifout_o_18),
	.exmem_ifout_o_21(exmem_ifout_o_21),
	.exmem_ifout_o_20(exmem_ifout_o_20),
	.exmem_ifout_o_23(exmem_ifout_o_23),
	.exmem_ifout_o_22(exmem_ifout_o_22),
	.exmem_ifout_o_25(exmem_ifout_o_25),
	.exmem_ifout_o_24(exmem_ifout_o_24),
	.exmem_ifout_o_27(exmem_ifout_o_27),
	.exmem_ifout_o_26(exmem_ifout_o_26),
	.exmem_ifout_o_29(exmem_ifout_o_29),
	.exmem_ifout_o_28(exmem_ifout_o_28),
	.exmem_ifout_o_31(exmem_ifout_o_31),
	.exmem_ifout_o_30(exmem_ifout_o_30),
	.always1(always1),
	.always11(always11),
	.exmem_ifhalt_o(\EXMEM|exmem_if.halt_o~q ),
	.exmem_ifrdat2_o_0(exmem_ifrdat2_o_0),
	.always12(always12),
	.idex_ifrt_o_0(\IDEX|idex_if.rt_o [0]),
	.idex_ifrt_o_1(\IDEX|idex_if.rt_o [1]),
	.exmem_ifRegDest_o_1(\EXMEM|exmem_if.RegDest_o [1]),
	.exmem_ifrt_o_1(\EXMEM|exmem_if.rt_o [1]),
	.exmem_ifrd_o_1(\EXMEM|exmem_if.rd_o [1]),
	.exmem_ifRegDest_o_0(\EXMEM|exmem_if.RegDest_o [0]),
	.exmem_ifrt_o_0(\EXMEM|exmem_if.rt_o [0]),
	.exmem_ifrd_o_0(\EXMEM|exmem_if.rd_o [0]),
	.idex_ifrt_o_2(\IDEX|idex_if.rt_o [2]),
	.idex_ifrt_o_3(\IDEX|idex_if.rt_o [3]),
	.exmem_ifrt_o_3(\EXMEM|exmem_if.rt_o [3]),
	.exmem_ifrd_o_3(\EXMEM|exmem_if.rd_o [3]),
	.exmem_ifrt_o_2(\EXMEM|exmem_if.rt_o [2]),
	.exmem_ifrd_o_2(\EXMEM|exmem_if.rd_o [2]),
	.exmem_ifregWEN_o(\EXMEM|exmem_if.regWEN_o~q ),
	.idex_ifrt_o_4(\IDEX|idex_if.rt_o [4]),
	.exmem_ifrt_o_4(\EXMEM|exmem_if.rt_o [4]),
	.exmem_ifrd_o_4(\EXMEM|exmem_if.rd_o [4]),
	.exmem_ifjal_o(\EXMEM|exmem_if.jal_o~q ),
	.exmem_iflui_o(\EXMEM|exmem_if.lui_o~q ),
	.exmem_ifnext_pc_o_1(\EXMEM|exmem_if.next_pc_o [1]),
	.exmem_ifmemToReg_o(\EXMEM|exmem_if.memToReg_o~q ),
	.fuifrtReplace_1(\FU|fuif.rtReplace[1]~4_combout ),
	.idex_ifimm_o_1(\IDEX|idex_if.imm_o [1]),
	.idex_ifrdat2_o_1(\IDEX|idex_if.rdat2_o [1]),
	.idex_ifimm_o_0(\IDEX|idex_if.imm_o [0]),
	.idex_ifrdat2_o_0(\IDEX|idex_if.rdat2_o [0]),
	.exmem_ifnext_pc_o_0(\EXMEM|exmem_if.next_pc_o [0]),
	.fuifrtReplace_0(\FU|fuif.rtReplace[0]~5_combout ),
	.exmem_ifnext_pc_o_2(\EXMEM|exmem_if.next_pc_o [2]),
	.exmem_ifnext_pc_o_4(\EXMEM|exmem_if.next_pc_o [4]),
	.exmem_ifnext_pc_o_3(\EXMEM|exmem_if.next_pc_o [3]),
	.idex_ifimm_o_2(\IDEX|idex_if.imm_o [2]),
	.idex_ifrdat2_o_2(\IDEX|idex_if.rdat2_o [2]),
	.fuifrtReplace_2(\FU|fuif.rtReplace[2]~6_combout ),
	.exmem_ifnext_pc_o_8(\EXMEM|exmem_if.next_pc_o [8]),
	.exmem_ifnext_pc_o_7(\EXMEM|exmem_if.next_pc_o [7]),
	.exmem_ifnext_pc_o_6(\EXMEM|exmem_if.next_pc_o [6]),
	.exmem_ifnext_pc_o_5(\EXMEM|exmem_if.next_pc_o [5]),
	.idex_ifrdat2_o_3(\IDEX|idex_if.rdat2_o [3]),
	.idex_ifimm_o_3(\IDEX|idex_if.imm_o [3]),
	.fuifrtReplace_3(\FU|fuif.rtReplace[3]~7_combout ),
	.exmem_ifimm_o_0(\EXMEM|exmem_if.imm_o [0]),
	.exmem_ifnext_pc_o_16(\EXMEM|exmem_if.next_pc_o [16]),
	.exmem_ifnext_pc_o_15(\EXMEM|exmem_if.next_pc_o [15]),
	.exmem_ifnext_pc_o_14(\EXMEM|exmem_if.next_pc_o [14]),
	.exmem_ifnext_pc_o_13(\EXMEM|exmem_if.next_pc_o [13]),
	.exmem_ifnext_pc_o_12(\EXMEM|exmem_if.next_pc_o [12]),
	.exmem_ifnext_pc_o_11(\EXMEM|exmem_if.next_pc_o [11]),
	.exmem_ifnext_pc_o_10(\EXMEM|exmem_if.next_pc_o [10]),
	.exmem_ifnext_pc_o_9(\EXMEM|exmem_if.next_pc_o [9]),
	.idex_ifrdat2_o_4(\IDEX|idex_if.rdat2_o [4]),
	.idex_ifimm_o_4(\IDEX|idex_if.imm_o [4]),
	.fuifrtReplace_4(\FU|fuif.rtReplace[4]~8_combout ),
	.exmem_ifnext_pc_o_31(\EXMEM|exmem_if.next_pc_o [31]),
	.exmem_ifimm_o_15(\EXMEM|exmem_if.imm_o [15]),
	.exmem_ifnext_pc_o_29(\EXMEM|exmem_if.next_pc_o [29]),
	.exmem_ifimm_o_13(\EXMEM|exmem_if.imm_o [13]),
	.exmem_ifimm_o_14(\EXMEM|exmem_if.imm_o [14]),
	.exmem_ifnext_pc_o_30(\EXMEM|exmem_if.next_pc_o [30]),
	.exmem_ifimm_o_12(\EXMEM|exmem_if.imm_o [12]),
	.exmem_ifnext_pc_o_28(\EXMEM|exmem_if.next_pc_o [28]),
	.exmem_ifimm_o_10(\EXMEM|exmem_if.imm_o [10]),
	.exmem_ifnext_pc_o_26(\EXMEM|exmem_if.next_pc_o [26]),
	.exmem_ifnext_pc_o_27(\EXMEM|exmem_if.next_pc_o [27]),
	.exmem_ifimm_o_11(\EXMEM|exmem_if.imm_o [11]),
	.exmem_ifnext_pc_o_25(\EXMEM|exmem_if.next_pc_o [25]),
	.exmem_ifimm_o_9(\EXMEM|exmem_if.imm_o [9]),
	.exmem_ifimm_o_8(\EXMEM|exmem_if.imm_o [8]),
	.exmem_ifnext_pc_o_24(\EXMEM|exmem_if.next_pc_o [24]),
	.exmem_ifimm_o_6(\EXMEM|exmem_if.imm_o [6]),
	.exmem_ifnext_pc_o_22(\EXMEM|exmem_if.next_pc_o [22]),
	.exmem_ifnext_pc_o_23(\EXMEM|exmem_if.next_pc_o [23]),
	.exmem_ifimm_o_7(\EXMEM|exmem_if.imm_o [7]),
	.exmem_ifnext_pc_o_21(\EXMEM|exmem_if.next_pc_o [21]),
	.exmem_ifimm_o_5(\EXMEM|exmem_if.imm_o [5]),
	.exmem_ifimm_o_4(\EXMEM|exmem_if.imm_o [4]),
	.exmem_ifnext_pc_o_20(\EXMEM|exmem_if.next_pc_o [20]),
	.exmem_ifimm_o_2(\EXMEM|exmem_if.imm_o [2]),
	.exmem_ifnext_pc_o_18(\EXMEM|exmem_if.next_pc_o [18]),
	.exmem_ifnext_pc_o_19(\EXMEM|exmem_if.next_pc_o [19]),
	.exmem_ifimm_o_3(\EXMEM|exmem_if.imm_o [3]),
	.exmem_ifnext_pc_o_17(\EXMEM|exmem_if.next_pc_o [17]),
	.exmem_ifimm_o_1(\EXMEM|exmem_if.imm_o [1]),
	.idex_ifimm_o_15(\IDEX|idex_if.imm_o [15]),
	.idex_ifrdat2_o_31(\IDEX|idex_if.rdat2_o [31]),
	.fuifrtReplace_31(\FU|fuif.rtReplace[31]~9_combout ),
	.idex_ifrdat2_o_16(\IDEX|idex_if.rdat2_o [16]),
	.fuifrtReplace_16(\FU|fuif.rtReplace[16]~10_combout ),
	.idex_ifrdat2_o_17(\IDEX|idex_if.rdat2_o [17]),
	.fuifrtReplace_17(\FU|fuif.rtReplace[17]~11_combout ),
	.idex_ifrdat2_o_18(\IDEX|idex_if.rdat2_o [18]),
	.fuifrtReplace_18(\FU|fuif.rtReplace[18]~12_combout ),
	.idex_ifrdat2_o_19(\IDEX|idex_if.rdat2_o [19]),
	.fuifrtReplace_19(\FU|fuif.rtReplace[19]~13_combout ),
	.idex_ifrdat2_o_20(\IDEX|idex_if.rdat2_o [20]),
	.fuifrtReplace_20(\FU|fuif.rtReplace[20]~14_combout ),
	.idex_ifrdat2_o_21(\IDEX|idex_if.rdat2_o [21]),
	.fuifrtReplace_21(\FU|fuif.rtReplace[21]~15_combout ),
	.idex_ifrdat2_o_22(\IDEX|idex_if.rdat2_o [22]),
	.fuifrtReplace_22(\FU|fuif.rtReplace[22]~16_combout ),
	.idex_ifrdat2_o_23(\IDEX|idex_if.rdat2_o [23]),
	.fuifrtReplace_23(\FU|fuif.rtReplace[23]~17_combout ),
	.idex_ifrdat2_o_24(\IDEX|idex_if.rdat2_o [24]),
	.fuifrtReplace_24(\FU|fuif.rtReplace[24]~18_combout ),
	.idex_ifrdat2_o_25(\IDEX|idex_if.rdat2_o [25]),
	.fuifrtReplace_25(\FU|fuif.rtReplace[25]~19_combout ),
	.idex_ifrdat2_o_26(\IDEX|idex_if.rdat2_o [26]),
	.fuifrtReplace_26(\FU|fuif.rtReplace[26]~20_combout ),
	.idex_ifrdat2_o_5(\IDEX|idex_if.rdat2_o [5]),
	.idex_ifimm_o_5(\IDEX|idex_if.imm_o [5]),
	.fuifrtReplace_5(\FU|fuif.rtReplace[5]~21_combout ),
	.idex_ifrdat2_o_6(\IDEX|idex_if.rdat2_o [6]),
	.idex_ifimm_o_6(\IDEX|idex_if.imm_o [6]),
	.fuifrtReplace_6(\FU|fuif.rtReplace[6]~22_combout ),
	.idex_ifrdat2_o_7(\IDEX|idex_if.rdat2_o [7]),
	.idex_ifimm_o_7(\IDEX|idex_if.imm_o [7]),
	.fuifrtReplace_7(\FU|fuif.rtReplace[7]~23_combout ),
	.idex_ifrdat2_o_8(\IDEX|idex_if.rdat2_o [8]),
	.idex_ifimm_o_8(\IDEX|idex_if.imm_o [8]),
	.fuifrtReplace_8(\FU|fuif.rtReplace[8]~24_combout ),
	.idex_ifrdat2_o_27(\IDEX|idex_if.rdat2_o [27]),
	.fuifrtReplace_27(\FU|fuif.rtReplace[27]~25_combout ),
	.idex_ifrdat2_o_28(\IDEX|idex_if.rdat2_o [28]),
	.fuifrtReplace_28(\FU|fuif.rtReplace[28]~26_combout ),
	.idex_ifrdat2_o_29(\IDEX|idex_if.rdat2_o [29]),
	.fuifrtReplace_29(\FU|fuif.rtReplace[29]~27_combout ),
	.idex_ifrdat2_o_30(\IDEX|idex_if.rdat2_o [30]),
	.fuifrtReplace_30(\FU|fuif.rtReplace[30]~28_combout ),
	.idex_ifrdat2_o_9(\IDEX|idex_if.rdat2_o [9]),
	.idex_ifimm_o_9(\IDEX|idex_if.imm_o [9]),
	.fuifrtReplace_9(\FU|fuif.rtReplace[9]~29_combout ),
	.idex_ifrdat2_o_14(\IDEX|idex_if.rdat2_o [14]),
	.idex_ifimm_o_14(\IDEX|idex_if.imm_o [14]),
	.fuifrtReplace_14(\FU|fuif.rtReplace[14]~30_combout ),
	.idex_ifrdat2_o_15(\IDEX|idex_if.rdat2_o [15]),
	.fuifrtReplace_15(\FU|fuif.rtReplace[15]~31_combout ),
	.idex_ifrdat2_o_10(\IDEX|idex_if.rdat2_o [10]),
	.idex_ifimm_o_10(\IDEX|idex_if.imm_o [10]),
	.fuifrtReplace_10(\FU|fuif.rtReplace[10]~32_combout ),
	.idex_ifrdat2_o_11(\IDEX|idex_if.rdat2_o [11]),
	.idex_ifimm_o_11(\IDEX|idex_if.imm_o [11]),
	.fuifrtReplace_11(\FU|fuif.rtReplace[11]~33_combout ),
	.idex_ifrdat2_o_12(\IDEX|idex_if.rdat2_o [12]),
	.idex_ifimm_o_12(\IDEX|idex_if.imm_o [12]),
	.fuifrtReplace_12(\FU|fuif.rtReplace[12]~34_combout ),
	.idex_ifrdat2_o_13(\IDEX|idex_if.rdat2_o [13]),
	.idex_ifimm_o_13(\IDEX|idex_if.imm_o [13]),
	.fuifrtReplace_13(\FU|fuif.rtReplace[13]~35_combout ),
	.idex_ifaluop_o_3(\IDEX|idex_if.aluop_o [3]),
	.myifout_1(\ALU|myif.out[1]~15_combout ),
	.ramstate(ramstate),
	.exmem_ifimm_o_01(\EXMEM|exmem_if.imm_o[0]~0_combout ),
	.idex_ifdWEN_o(\IDEX|idex_if.dWEN_o~q ),
	.idex_ifdREN_o(\IDEX|idex_if.dREN_o~q ),
	.idex_ifnext_pc_o_1(\IDEX|idex_if.next_pc_o [1]),
	.myifout_6(\ALU|myif.out[6]~26_combout ),
	.myifout_4(\ALU|myif.out[4]~33_combout ),
	.myifout_24(\ALU|myif.out[24]~40_combout ),
	.myifout_26(\ALU|myif.out[26]~47_combout ),
	.myifout_25(\ALU|myif.out[25]~54_combout ),
	.myifout_27(\ALU|myif.out[27]~61_combout ),
	.myifout_5(\ALU|myif.out[5]~68_combout ),
	.myifout_7(\ALU|myif.out[7]~81_combout ),
	.myifout_13(\ALU|myif.out[13]~92_combout ),
	.myifout_9(\ALU|myif.out[9]~98_combout ),
	.myifout_8(\ALU|myif.out[8]~104_combout ),
	.myifout_14(\ALU|myif.out[14]~110_combout ),
	.myifout_12(\ALU|myif.out[12]~116_combout ),
	.myifout_15(\ALU|myif.out[15]~122_combout ),
	.myifout_10(\ALU|myif.out[10]~128_combout ),
	.myifout_11(\ALU|myif.out[11]~134_combout ),
	.myifout_23(\ALU|myif.out[23]~152_combout ),
	.myifout_16(\ALU|myif.out[16]~158_combout ),
	.myifout_17(\ALU|myif.out[17]~174_combout ),
	.myifout_18(\ALU|myif.out[18]~180_combout ),
	.myifout_19(\ALU|myif.out[19]~196_combout ),
	.myifout_30(\ALU|myif.out[30]~204_combout ),
	.myifout_21(\ALU|myif.out[21]~220_combout ),
	.myifnegative(\ALU|myif.negative~8_combout ),
	.myifout_22(\ALU|myif.out[22]~226_combout ),
	.myifout_20(\ALU|myif.out[20]~232_combout ),
	.myifout_0(\ALU|myif.out[0]~239_combout ),
	.myifout_28(\ALU|myif.out[28]~252_combout ),
	.myifout_29(\ALU|myif.out[29]~264_combout ),
	.myifout_2(\ALU|myif.out[2]~274_combout ),
	.myifout_3(\ALU|myif.out[3]~283_combout ),
	.myifout_31(\ALU|myif.out[3]~285_combout ),
	.myifout_210(\ALU|myif.out[2]~289_combout ),
	.idex_ifnext_pc_o_0(\IDEX|idex_if.next_pc_o [0]),
	.idex_ifnext_pc_o_3(\IDEX|idex_if.next_pc_o [3]),
	.idex_ifnext_pc_o_2(\IDEX|idex_if.next_pc_o [2]),
	.idex_ifnext_pc_o_5(\IDEX|idex_if.next_pc_o [5]),
	.idex_ifnext_pc_o_4(\IDEX|idex_if.next_pc_o [4]),
	.idex_ifnext_pc_o_7(\IDEX|idex_if.next_pc_o [7]),
	.idex_ifnext_pc_o_6(\IDEX|idex_if.next_pc_o [6]),
	.idex_ifnext_pc_o_9(\IDEX|idex_if.next_pc_o [9]),
	.idex_ifnext_pc_o_8(\IDEX|idex_if.next_pc_o [8]),
	.idex_ifnext_pc_o_11(\IDEX|idex_if.next_pc_o [11]),
	.idex_ifnext_pc_o_10(\IDEX|idex_if.next_pc_o [10]),
	.idex_ifnext_pc_o_13(\IDEX|idex_if.next_pc_o [13]),
	.idex_ifnext_pc_o_12(\IDEX|idex_if.next_pc_o [12]),
	.idex_ifnext_pc_o_15(\IDEX|idex_if.next_pc_o [15]),
	.idex_ifnext_pc_o_14(\IDEX|idex_if.next_pc_o [14]),
	.idex_ifnext_pc_o_17(\IDEX|idex_if.next_pc_o [17]),
	.idex_ifnext_pc_o_16(\IDEX|idex_if.next_pc_o [16]),
	.idex_ifnext_pc_o_19(\IDEX|idex_if.next_pc_o [19]),
	.idex_ifnext_pc_o_18(\IDEX|idex_if.next_pc_o [18]),
	.idex_ifnext_pc_o_21(\IDEX|idex_if.next_pc_o [21]),
	.idex_ifnext_pc_o_20(\IDEX|idex_if.next_pc_o [20]),
	.idex_ifnext_pc_o_23(\IDEX|idex_if.next_pc_o [23]),
	.idex_ifnext_pc_o_22(\IDEX|idex_if.next_pc_o [22]),
	.idex_ifnext_pc_o_25(\IDEX|idex_if.next_pc_o [25]),
	.idex_ifnext_pc_o_24(\IDEX|idex_if.next_pc_o [24]),
	.idex_ifnext_pc_o_27(\IDEX|idex_if.next_pc_o [27]),
	.idex_ifnext_pc_o_26(\IDEX|idex_if.next_pc_o [26]),
	.idex_ifnext_pc_o_29(\IDEX|idex_if.next_pc_o [29]),
	.idex_ifnext_pc_o_28(\IDEX|idex_if.next_pc_o [28]),
	.idex_ifnext_pc_o_31(\IDEX|idex_if.next_pc_o [31]),
	.idex_ifnext_pc_o_30(\IDEX|idex_if.next_pc_o [30]),
	.exmem_ifrdat2_o_1(exmem_ifrdat2_o_1),
	.exmem_ifrdat2_o_2(exmem_ifrdat2_o_2),
	.exmem_ifrdat2_o_3(exmem_ifrdat2_o_3),
	.exmem_ifrdat2_o_4(exmem_ifrdat2_o_4),
	.exmem_ifrdat2_o_5(exmem_ifrdat2_o_5),
	.exmem_ifrdat2_o_6(exmem_ifrdat2_o_6),
	.exmem_ifrdat2_o_7(exmem_ifrdat2_o_7),
	.exmem_ifrdat2_o_8(exmem_ifrdat2_o_8),
	.exmem_ifrdat2_o_9(exmem_ifrdat2_o_9),
	.exmem_ifrdat2_o_10(exmem_ifrdat2_o_10),
	.exmem_ifrdat2_o_11(exmem_ifrdat2_o_11),
	.exmem_ifrdat2_o_12(exmem_ifrdat2_o_12),
	.exmem_ifrdat2_o_13(exmem_ifrdat2_o_13),
	.exmem_ifrdat2_o_14(exmem_ifrdat2_o_14),
	.exmem_ifrdat2_o_15(exmem_ifrdat2_o_15),
	.exmem_ifrdat2_o_16(exmem_ifrdat2_o_16),
	.exmem_ifrdat2_o_17(exmem_ifrdat2_o_17),
	.exmem_ifrdat2_o_18(exmem_ifrdat2_o_18),
	.exmem_ifrdat2_o_19(exmem_ifrdat2_o_19),
	.exmem_ifrdat2_o_20(exmem_ifrdat2_o_20),
	.exmem_ifrdat2_o_21(exmem_ifrdat2_o_21),
	.exmem_ifrdat2_o_22(exmem_ifrdat2_o_22),
	.exmem_ifrdat2_o_23(exmem_ifrdat2_o_23),
	.exmem_ifrdat2_o_24(exmem_ifrdat2_o_24),
	.exmem_ifrdat2_o_25(exmem_ifrdat2_o_25),
	.exmem_ifrdat2_o_26(exmem_ifrdat2_o_26),
	.exmem_ifrdat2_o_27(exmem_ifrdat2_o_27),
	.exmem_ifrdat2_o_28(exmem_ifrdat2_o_28),
	.exmem_ifrdat2_o_29(exmem_ifrdat2_o_29),
	.exmem_ifrdat2_o_30(exmem_ifrdat2_o_30),
	.exmem_ifrdat2_o_31(exmem_ifrdat2_o_31),
	.idex_ifhalt_o(\IDEX|idex_if.halt_o~q ),
	.fuifrdat2_ow(\FU|fuif.rdat2_ow~0_combout ),
	.idex_ifRegDest_o_1(\IDEX|idex_if.RegDest_o [1]),
	.idex_ifrd_o_1(\IDEX|idex_if.rd_o [1]),
	.idex_ifRegDest_o_0(\IDEX|idex_if.RegDest_o [0]),
	.idex_ifrd_o_0(\IDEX|idex_if.rd_o [0]),
	.idex_ifrd_o_3(\IDEX|idex_if.rd_o [3]),
	.idex_ifrd_o_2(\IDEX|idex_if.rd_o [2]),
	.idex_ifregWEN_o(\IDEX|idex_if.regWEN_o~q ),
	.idex_ifrd_o_4(\IDEX|idex_if.rd_o [4]),
	.idex_ifjal_o(\IDEX|idex_if.jal_o~q ),
	.idex_iflui_o(\IDEX|idex_if.lui_o~q ),
	.idex_ifmemToReg_o(\IDEX|idex_if.memToReg_o~q ),
	.myifout_32(\ALU|myif.out[3]~291_combout ),
	.CPUCLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

id_ex IDEX(
	.idex_ifaluop_o_1(\IDEX|idex_if.aluop_o [1]),
	.idex_ifrt_o_0(\IDEX|idex_if.rt_o [0]),
	.idex_ifrt_o_1(\IDEX|idex_if.rt_o [1]),
	.idex_ifrt_o_2(\IDEX|idex_if.rt_o [2]),
	.idex_ifrt_o_3(\IDEX|idex_if.rt_o [3]),
	.idex_ifrt_o_4(\IDEX|idex_if.rt_o [4]),
	.idex_ifALUSel_o_1(\IDEX|idex_if.ALUSel_o [1]),
	.idex_ifALUSel_o_0(\IDEX|idex_if.ALUSel_o [0]),
	.idex_ifimm_o_1(\IDEX|idex_if.imm_o [1]),
	.idex_ifshamt_o_1(\IDEX|idex_if.shamt_o [1]),
	.idex_ifrdat2_o_1(\IDEX|idex_if.rdat2_o [1]),
	.idex_ifrdat1_o_1(\IDEX|idex_if.rdat1_o [1]),
	.idex_ifrs_o_1(\IDEX|idex_if.rs_o [1]),
	.idex_ifrs_o_0(\IDEX|idex_if.rs_o [0]),
	.idex_ifrs_o_3(\IDEX|idex_if.rs_o [3]),
	.idex_ifrs_o_2(\IDEX|idex_if.rs_o [2]),
	.idex_ifrs_o_4(\IDEX|idex_if.rs_o [4]),
	.idex_ifimm_o_0(\IDEX|idex_if.imm_o [0]),
	.idex_ifshamt_o_0(\IDEX|idex_if.shamt_o [0]),
	.idex_ifrdat2_o_0(\IDEX|idex_if.rdat2_o [0]),
	.idex_ifrdat1_o_0(\IDEX|idex_if.rdat1_o [0]),
	.idex_ifaluop_o_2(\IDEX|idex_if.aluop_o [2]),
	.idex_ifrdat1_o_2(\IDEX|idex_if.rdat1_o [2]),
	.idex_ifrdat1_o_4(\IDEX|idex_if.rdat1_o [4]),
	.idex_ifrdat1_o_3(\IDEX|idex_if.rdat1_o [3]),
	.idex_ifimm_o_2(\IDEX|idex_if.imm_o [2]),
	.idex_ifshamt_o_2(\IDEX|idex_if.shamt_o [2]),
	.idex_ifrdat2_o_2(\IDEX|idex_if.rdat2_o [2]),
	.idex_ifrdat1_o_8(\IDEX|idex_if.rdat1_o [8]),
	.idex_ifrdat1_o_7(\IDEX|idex_if.rdat1_o [7]),
	.idex_ifrdat1_o_6(\IDEX|idex_if.rdat1_o [6]),
	.idex_ifrdat1_o_5(\IDEX|idex_if.rdat1_o [5]),
	.idex_ifrdat2_o_3(\IDEX|idex_if.rdat2_o [3]),
	.idex_ifimm_o_3(\IDEX|idex_if.imm_o [3]),
	.idex_ifshamt_o_3(\IDEX|idex_if.shamt_o [3]),
	.idex_ifrdat1_o_16(\IDEX|idex_if.rdat1_o [16]),
	.idex_ifrdat1_o_15(\IDEX|idex_if.rdat1_o [15]),
	.idex_ifrdat1_o_14(\IDEX|idex_if.rdat1_o [14]),
	.idex_ifrdat1_o_13(\IDEX|idex_if.rdat1_o [13]),
	.idex_ifrdat1_o_12(\IDEX|idex_if.rdat1_o [12]),
	.idex_ifrdat1_o_11(\IDEX|idex_if.rdat1_o [11]),
	.idex_ifrdat1_o_10(\IDEX|idex_if.rdat1_o [10]),
	.idex_ifrdat1_o_9(\IDEX|idex_if.rdat1_o [9]),
	.idex_ifrdat2_o_4(\IDEX|idex_if.rdat2_o [4]),
	.idex_ifimm_o_4(\IDEX|idex_if.imm_o [4]),
	.idex_ifshamt_o_4(\IDEX|idex_if.shamt_o [4]),
	.idex_ifrdat1_o_31(\IDEX|idex_if.rdat1_o [31]),
	.idex_ifrdat1_o_29(\IDEX|idex_if.rdat1_o [29]),
	.idex_ifrdat1_o_30(\IDEX|idex_if.rdat1_o [30]),
	.idex_ifrdat1_o_28(\IDEX|idex_if.rdat1_o [28]),
	.idex_ifrdat1_o_26(\IDEX|idex_if.rdat1_o [26]),
	.idex_ifrdat1_o_27(\IDEX|idex_if.rdat1_o [27]),
	.idex_ifrdat1_o_25(\IDEX|idex_if.rdat1_o [25]),
	.idex_ifrdat1_o_24(\IDEX|idex_if.rdat1_o [24]),
	.idex_ifrdat1_o_22(\IDEX|idex_if.rdat1_o [22]),
	.idex_ifrdat1_o_23(\IDEX|idex_if.rdat1_o [23]),
	.idex_ifrdat1_o_21(\IDEX|idex_if.rdat1_o [21]),
	.idex_ifrdat1_o_20(\IDEX|idex_if.rdat1_o [20]),
	.idex_ifrdat1_o_18(\IDEX|idex_if.rdat1_o [18]),
	.idex_ifrdat1_o_19(\IDEX|idex_if.rdat1_o [19]),
	.idex_ifrdat1_o_17(\IDEX|idex_if.rdat1_o [17]),
	.idex_ifimm_o_15(\IDEX|idex_if.imm_o [15]),
	.idex_ifrdat2_o_31(\IDEX|idex_if.rdat2_o [31]),
	.idex_ifrdat2_o_16(\IDEX|idex_if.rdat2_o [16]),
	.idex_ifrdat2_o_17(\IDEX|idex_if.rdat2_o [17]),
	.idex_ifrdat2_o_18(\IDEX|idex_if.rdat2_o [18]),
	.idex_ifrdat2_o_19(\IDEX|idex_if.rdat2_o [19]),
	.idex_ifrdat2_o_20(\IDEX|idex_if.rdat2_o [20]),
	.idex_ifrdat2_o_21(\IDEX|idex_if.rdat2_o [21]),
	.idex_ifrdat2_o_22(\IDEX|idex_if.rdat2_o [22]),
	.idex_ifrdat2_o_23(\IDEX|idex_if.rdat2_o [23]),
	.idex_ifrdat2_o_24(\IDEX|idex_if.rdat2_o [24]),
	.idex_ifrdat2_o_25(\IDEX|idex_if.rdat2_o [25]),
	.idex_ifrdat2_o_26(\IDEX|idex_if.rdat2_o [26]),
	.idex_ifrdat2_o_5(\IDEX|idex_if.rdat2_o [5]),
	.idex_ifimm_o_5(\IDEX|idex_if.imm_o [5]),
	.idex_ifrdat2_o_6(\IDEX|idex_if.rdat2_o [6]),
	.idex_ifimm_o_6(\IDEX|idex_if.imm_o [6]),
	.idex_ifrdat2_o_7(\IDEX|idex_if.rdat2_o [7]),
	.idex_ifimm_o_7(\IDEX|idex_if.imm_o [7]),
	.idex_ifrdat2_o_8(\IDEX|idex_if.rdat2_o [8]),
	.idex_ifimm_o_8(\IDEX|idex_if.imm_o [8]),
	.idex_ifrdat2_o_27(\IDEX|idex_if.rdat2_o [27]),
	.idex_ifrdat2_o_28(\IDEX|idex_if.rdat2_o [28]),
	.idex_ifrdat2_o_29(\IDEX|idex_if.rdat2_o [29]),
	.idex_ifrdat2_o_30(\IDEX|idex_if.rdat2_o [30]),
	.idex_ifrdat2_o_9(\IDEX|idex_if.rdat2_o [9]),
	.idex_ifimm_o_9(\IDEX|idex_if.imm_o [9]),
	.idex_ifrdat2_o_14(\IDEX|idex_if.rdat2_o [14]),
	.idex_ifimm_o_14(\IDEX|idex_if.imm_o [14]),
	.idex_ifrdat2_o_15(\IDEX|idex_if.rdat2_o [15]),
	.idex_ifrdat2_o_10(\IDEX|idex_if.rdat2_o [10]),
	.idex_ifimm_o_10(\IDEX|idex_if.imm_o [10]),
	.idex_ifrdat2_o_11(\IDEX|idex_if.rdat2_o [11]),
	.idex_ifimm_o_11(\IDEX|idex_if.imm_o [11]),
	.idex_ifrdat2_o_12(\IDEX|idex_if.rdat2_o [12]),
	.idex_ifimm_o_12(\IDEX|idex_if.imm_o [12]),
	.idex_ifrdat2_o_13(\IDEX|idex_if.rdat2_o [13]),
	.idex_ifimm_o_13(\IDEX|idex_if.imm_o [13]),
	.idex_ifaluop_o_0(\IDEX|idex_if.aluop_o [0]),
	.idex_ifaluop_o_3(\IDEX|idex_if.aluop_o [3]),
	.idex_ifdWEN_o(\IDEX|idex_if.dWEN_o~q ),
	.idex_ifdREN_o(\IDEX|idex_if.dREN_o~q ),
	.idex_ifnext_pc_o_1(\IDEX|idex_if.next_pc_o [1]),
	.idex_ifjumpSel_o_1(\IDEX|idex_if.jumpSel_o [1]),
	.idex_ifjumpSel_o_0(\IDEX|idex_if.jumpSel_o [0]),
	.always1(always13),
	.idex_ifinstr_o_31(\IDEX|idex_if.instr_o [31]),
	.idex_ifinstr_o_30(\IDEX|idex_if.instr_o [30]),
	.idex_ifinstr_o_27(\IDEX|idex_if.instr_o [27]),
	.idex_ifinstr_o_26(\IDEX|idex_if.instr_o [26]),
	.idex_ifinstr_o_28(\IDEX|idex_if.instr_o [28]),
	.ifid_ifinstr_o_17(\IFID|ifid_if.instr_o [17]),
	.ifid_ifinstr_o_16(\IFID|ifid_if.instr_o [16]),
	.ifid_ifinstr_o_19(\IFID|ifid_if.instr_o [19]),
	.ifid_ifinstr_o_18(\IFID|ifid_if.instr_o [18]),
	.ifid_ifinstr_o_20(\IFID|ifid_if.instr_o [20]),
	.ifid_ifinstr_o_22(\IFID|ifid_if.instr_o [22]),
	.ifid_ifinstr_o_21(\IFID|ifid_if.instr_o [21]),
	.ifid_ifinstr_o_24(\IFID|ifid_if.instr_o [24]),
	.ifid_ifinstr_o_23(\IFID|ifid_if.instr_o [23]),
	.ifid_ifinstr_o_25(\IFID|ifid_if.instr_o [25]),
	.huiffreeze(\HU|huif.freeze~2_combout ),
	.idex_ifbne_o(\IDEX|idex_if.bne_o~q ),
	.idex_ifPCSel_o(\IDEX|idex_if.PCSel_o~q ),
	.huifflush(\HU|huif.flush~0_combout ),
	.idex_ifnext_pc_o_0(\IDEX|idex_if.next_pc_o [0]),
	.idex_ifnext_pc_o_3(\IDEX|idex_if.next_pc_o [3]),
	.idex_ifnext_pc_o_2(\IDEX|idex_if.next_pc_o [2]),
	.idex_ifimm_26_o_1(\IDEX|idex_if.imm_26_o [1]),
	.idex_ifimm_26_o_0(\IDEX|idex_if.imm_26_o [0]),
	.idex_ifnext_pc_o_5(\IDEX|idex_if.next_pc_o [5]),
	.idex_ifnext_pc_o_4(\IDEX|idex_if.next_pc_o [4]),
	.idex_ifimm_26_o_3(\IDEX|idex_if.imm_26_o [3]),
	.idex_ifimm_26_o_2(\IDEX|idex_if.imm_26_o [2]),
	.idex_ifnext_pc_o_7(\IDEX|idex_if.next_pc_o [7]),
	.idex_ifnext_pc_o_6(\IDEX|idex_if.next_pc_o [6]),
	.idex_ifimm_26_o_5(\IDEX|idex_if.imm_26_o [5]),
	.idex_ifimm_26_o_4(\IDEX|idex_if.imm_26_o [4]),
	.idex_ifnext_pc_o_9(\IDEX|idex_if.next_pc_o [9]),
	.idex_ifnext_pc_o_8(\IDEX|idex_if.next_pc_o [8]),
	.idex_ifimm_26_o_7(\IDEX|idex_if.imm_26_o [7]),
	.idex_ifimm_26_o_6(\IDEX|idex_if.imm_26_o [6]),
	.idex_ifnext_pc_o_11(\IDEX|idex_if.next_pc_o [11]),
	.idex_ifnext_pc_o_10(\IDEX|idex_if.next_pc_o [10]),
	.idex_ifimm_26_o_9(\IDEX|idex_if.imm_26_o [9]),
	.idex_ifimm_26_o_8(\IDEX|idex_if.imm_26_o [8]),
	.idex_ifnext_pc_o_13(\IDEX|idex_if.next_pc_o [13]),
	.idex_ifnext_pc_o_12(\IDEX|idex_if.next_pc_o [12]),
	.idex_ifimm_26_o_11(\IDEX|idex_if.imm_26_o [11]),
	.idex_ifimm_26_o_10(\IDEX|idex_if.imm_26_o [10]),
	.idex_ifnext_pc_o_15(\IDEX|idex_if.next_pc_o [15]),
	.idex_ifnext_pc_o_14(\IDEX|idex_if.next_pc_o [14]),
	.idex_ifimm_26_o_13(\IDEX|idex_if.imm_26_o [13]),
	.idex_ifimm_26_o_12(\IDEX|idex_if.imm_26_o [12]),
	.idex_ifnext_pc_o_17(\IDEX|idex_if.next_pc_o [17]),
	.idex_ifnext_pc_o_16(\IDEX|idex_if.next_pc_o [16]),
	.idex_ifimm_26_o_15(\IDEX|idex_if.imm_26_o [15]),
	.idex_ifimm_26_o_14(\IDEX|idex_if.imm_26_o [14]),
	.idex_ifnext_pc_o_19(\IDEX|idex_if.next_pc_o [19]),
	.idex_ifnext_pc_o_18(\IDEX|idex_if.next_pc_o [18]),
	.idex_ifimm_26_o_17(\IDEX|idex_if.imm_26_o [17]),
	.idex_ifimm_26_o_16(\IDEX|idex_if.imm_26_o [16]),
	.idex_ifnext_pc_o_21(\IDEX|idex_if.next_pc_o [21]),
	.idex_ifnext_pc_o_20(\IDEX|idex_if.next_pc_o [20]),
	.idex_ifimm_26_o_19(\IDEX|idex_if.imm_26_o [19]),
	.idex_ifimm_26_o_18(\IDEX|idex_if.imm_26_o [18]),
	.idex_ifnext_pc_o_23(\IDEX|idex_if.next_pc_o [23]),
	.idex_ifnext_pc_o_22(\IDEX|idex_if.next_pc_o [22]),
	.idex_ifimm_26_o_21(\IDEX|idex_if.imm_26_o [21]),
	.idex_ifimm_26_o_20(\IDEX|idex_if.imm_26_o [20]),
	.idex_ifnext_pc_o_25(\IDEX|idex_if.next_pc_o [25]),
	.idex_ifnext_pc_o_24(\IDEX|idex_if.next_pc_o [24]),
	.idex_ifimm_26_o_23(\IDEX|idex_if.imm_26_o [23]),
	.idex_ifimm_26_o_22(\IDEX|idex_if.imm_26_o [22]),
	.idex_ifnext_pc_o_27(\IDEX|idex_if.next_pc_o [27]),
	.idex_ifnext_pc_o_26(\IDEX|idex_if.next_pc_o [26]),
	.idex_ifimm_26_o_25(\IDEX|idex_if.imm_26_o [25]),
	.idex_ifimm_26_o_24(\IDEX|idex_if.imm_26_o [24]),
	.idex_ifnext_pc_o_29(\IDEX|idex_if.next_pc_o [29]),
	.idex_ifnext_pc_o_28(\IDEX|idex_if.next_pc_o [28]),
	.idex_ifnext_pc_o_31(\IDEX|idex_if.next_pc_o [31]),
	.idex_ifnext_pc_o_30(\IDEX|idex_if.next_pc_o [30]),
	.idex_ifhalt_o(\IDEX|idex_if.halt_o~q ),
	.ifid_ifinstr_o_26(\IFID|ifid_if.instr_o [26]),
	.ifid_ifinstr_o_31(\IFID|ifid_if.instr_o [31]),
	.ifid_ifinstr_o_27(\IFID|ifid_if.instr_o [27]),
	.ifid_ifinstr_o_28(\IFID|ifid_if.instr_o [28]),
	.ifid_ifinstr_o_30(\IFID|ifid_if.instr_o [30]),
	.ifid_ifinstr_o_5(\IFID|ifid_if.instr_o [5]),
	.ifid_ifinstr_o_4(\IFID|ifid_if.instr_o [4]),
	.always0(\CU|always0~0_combout ),
	.ifid_ifinstr_o_29(\IFID|ifid_if.instr_o [29]),
	.ifid_ifinstr_o_1(\IFID|ifid_if.instr_o [1]),
	.ifid_ifinstr_o_3(\IFID|ifid_if.instr_o [3]),
	.ifid_ifinstr_o_2(\IFID|ifid_if.instr_o [2]),
	.idex_ifRegDest_o_1(\IDEX|idex_if.RegDest_o [1]),
	.idex_ifrd_o_1(\IDEX|idex_if.rd_o [1]),
	.idex_ifRegDest_o_0(\IDEX|idex_if.RegDest_o [0]),
	.idex_ifrd_o_0(\IDEX|idex_if.rd_o [0]),
	.idex_ifrd_o_3(\IDEX|idex_if.rd_o [3]),
	.idex_ifrd_o_2(\IDEX|idex_if.rd_o [2]),
	.idex_ifregWEN_o(\IDEX|idex_if.regWEN_o~q ),
	.idex_ifrd_o_4(\IDEX|idex_if.rd_o [4]),
	.cuifregWEN(\CU|cuif.regWEN~0_combout ),
	.Equal0(\CU|Equal0~0_combout ),
	.ifid_ifinstr_o_0(\IFID|ifid_if.instr_o [0]),
	.Equal3(\CU|Equal3~0_combout ),
	.Equal2(\CU|Equal2~0_combout ),
	.idex_ifjal_o(\IDEX|idex_if.jal_o~q ),
	.idex_iflui_o(\IDEX|idex_if.lui_o~q ),
	.idex_ifmemToReg_o(\IDEX|idex_if.memToReg_o~q ),
	.ifid_ifinstr_o_7(\IFID|ifid_if.instr_o [7]),
	.Mux62(\RF|Mux62~9_combout ),
	.Mux621(\RF|Mux62~19_combout ),
	.Mux30(\RF|Mux30~9_combout ),
	.Mux301(\RF|Mux30~19_combout ),
	.ifid_ifinstr_o_6(\IFID|ifid_if.instr_o [6]),
	.Mux63(\RF|Mux63~9_combout ),
	.Mux631(\RF|Mux63~19_combout ),
	.Mux31(\RF|Mux31~9_combout ),
	.Mux311(\RF|Mux31~19_combout ),
	.Equal10(\CU|Equal10~0_combout ),
	.Mux29(\RF|Mux29~9_combout ),
	.Mux291(\RF|Mux29~19_combout ),
	.Mux27(\RF|Mux27~9_combout ),
	.Mux271(\RF|Mux27~19_combout ),
	.Mux28(\RF|Mux28~9_combout ),
	.Mux281(\RF|Mux28~19_combout ),
	.ifid_ifinstr_o_8(\IFID|ifid_if.instr_o [8]),
	.Mux61(\RF|Mux61~9_combout ),
	.Mux611(\RF|Mux61~19_combout ),
	.Mux23(\RF|Mux23~9_combout ),
	.Mux231(\RF|Mux23~19_combout ),
	.Mux24(\RF|Mux24~9_combout ),
	.Mux241(\RF|Mux24~19_combout ),
	.Mux25(\RF|Mux25~9_combout ),
	.Mux251(\RF|Mux25~19_combout ),
	.Mux26(\RF|Mux26~9_combout ),
	.Mux261(\RF|Mux26~19_combout ),
	.Mux60(\RF|Mux60~9_combout ),
	.Mux601(\RF|Mux60~19_combout ),
	.ifid_ifinstr_o_9(\IFID|ifid_if.instr_o [9]),
	.Mux15(\RF|Mux15~9_combout ),
	.Mux151(\RF|Mux15~19_combout ),
	.Mux16(\RF|Mux16~9_combout ),
	.Mux161(\RF|Mux16~19_combout ),
	.Mux17(\RF|Mux17~9_combout ),
	.Mux171(\RF|Mux17~19_combout ),
	.Mux18(\RF|Mux18~9_combout ),
	.Mux181(\RF|Mux18~19_combout ),
	.Mux19(\RF|Mux19~9_combout ),
	.Mux191(\RF|Mux19~19_combout ),
	.Mux20(\RF|Mux20~9_combout ),
	.Mux201(\RF|Mux20~19_combout ),
	.Mux21(\RF|Mux21~9_combout ),
	.Mux211(\RF|Mux21~19_combout ),
	.Mux22(\RF|Mux22~9_combout ),
	.Mux221(\RF|Mux22~19_combout ),
	.Mux59(\RF|Mux59~9_combout ),
	.Mux591(\RF|Mux59~19_combout ),
	.ifid_ifinstr_o_10(\IFID|ifid_if.instr_o [10]),
	.Mux0(\RF|Mux0~9_combout ),
	.Mux01(\RF|Mux0~19_combout ),
	.Mux2(\RF|Mux2~9_combout ),
	.Mux210(\RF|Mux2~19_combout ),
	.Mux1(\RF|Mux1~9_combout ),
	.Mux11(\RF|Mux1~19_combout ),
	.Mux3(\RF|Mux3~9_combout ),
	.Mux32(\RF|Mux3~19_combout ),
	.Mux5(\RF|Mux5~9_combout ),
	.Mux51(\RF|Mux5~19_combout ),
	.Mux4(\RF|Mux4~9_combout ),
	.Mux41(\RF|Mux4~19_combout ),
	.Mux6(\RF|Mux6~9_combout ),
	.Mux64(\RF|Mux6~19_combout ),
	.Mux7(\RF|Mux7~9_combout ),
	.Mux71(\RF|Mux7~19_combout ),
	.Mux9(\RF|Mux9~9_combout ),
	.Mux91(\RF|Mux9~19_combout ),
	.Mux8(\RF|Mux8~9_combout ),
	.Mux81(\RF|Mux8~19_combout ),
	.Mux10(\RF|Mux10~9_combout ),
	.Mux101(\RF|Mux10~19_combout ),
	.Mux111(\RF|Mux11~9_combout ),
	.Mux112(\RF|Mux11~19_combout ),
	.Mux13(\RF|Mux13~9_combout ),
	.Mux131(\RF|Mux13~19_combout ),
	.Mux12(\RF|Mux12~9_combout ),
	.Mux121(\RF|Mux12~19_combout ),
	.Mux14(\RF|Mux14~9_combout ),
	.Mux141(\RF|Mux14~19_combout ),
	.ifid_ifinstr_o_15(\IFID|ifid_if.instr_o [15]),
	.Mux321(\RF|Mux32~9_combout ),
	.Mux322(\RF|Mux32~19_combout ),
	.Mux47(\RF|Mux47~9_combout ),
	.Mux471(\RF|Mux47~19_combout ),
	.Mux46(\RF|Mux46~9_combout ),
	.Mux461(\RF|Mux46~19_combout ),
	.Mux45(\RF|Mux45~9_combout ),
	.Mux451(\RF|Mux45~19_combout ),
	.Mux44(\RF|Mux44~9_combout ),
	.Mux441(\RF|Mux44~19_combout ),
	.Mux43(\RF|Mux43~9_combout ),
	.Mux431(\RF|Mux43~19_combout ),
	.Mux42(\RF|Mux42~9_combout ),
	.Mux421(\RF|Mux42~19_combout ),
	.Mux411(\RF|Mux41~9_combout ),
	.Mux412(\RF|Mux41~19_combout ),
	.Mux40(\RF|Mux40~9_combout ),
	.Mux401(\RF|Mux40~19_combout ),
	.Mux39(\RF|Mux39~9_combout ),
	.Mux391(\RF|Mux39~19_combout ),
	.Mux38(\RF|Mux38~9_combout ),
	.Mux381(\RF|Mux38~19_combout ),
	.Mux37(\RF|Mux37~9_combout ),
	.Mux371(\RF|Mux37~19_combout ),
	.Mux58(\RF|Mux58~9_combout ),
	.Mux581(\RF|Mux58~19_combout ),
	.Mux57(\RF|Mux57~9_combout ),
	.Mux571(\RF|Mux57~19_combout ),
	.Mux56(\RF|Mux56~9_combout ),
	.Mux561(\RF|Mux56~19_combout ),
	.Mux55(\RF|Mux55~9_combout ),
	.Mux551(\RF|Mux55~19_combout ),
	.Mux36(\RF|Mux36~9_combout ),
	.Mux361(\RF|Mux36~19_combout ),
	.Mux35(\RF|Mux35~9_combout ),
	.Mux351(\RF|Mux35~19_combout ),
	.Mux34(\RF|Mux34~9_combout ),
	.Mux341(\RF|Mux34~19_combout ),
	.Mux33(\RF|Mux33~9_combout ),
	.Mux331(\RF|Mux33~19_combout ),
	.Mux54(\RF|Mux54~9_combout ),
	.Mux541(\RF|Mux54~19_combout ),
	.Mux49(\RF|Mux49~9_combout ),
	.Mux491(\RF|Mux49~19_combout ),
	.ifid_ifinstr_o_14(\IFID|ifid_if.instr_o [14]),
	.Mux48(\RF|Mux48~9_combout ),
	.Mux481(\RF|Mux48~19_combout ),
	.Mux53(\RF|Mux53~9_combout ),
	.Mux531(\RF|Mux53~19_combout ),
	.Mux52(\RF|Mux52~9_combout ),
	.Mux521(\RF|Mux52~19_combout ),
	.ifid_ifinstr_o_11(\IFID|ifid_if.instr_o [11]),
	.Mux511(\RF|Mux51~9_combout ),
	.Mux512(\RF|Mux51~19_combout ),
	.ifid_ifinstr_o_12(\IFID|ifid_if.instr_o [12]),
	.Mux50(\RF|Mux50~9_combout ),
	.Mux501(\RF|Mux50~19_combout ),
	.ifid_ifinstr_o_13(\IFID|ifid_if.instr_o [13]),
	.Equal14(\CU|Equal14~0_combout ),
	.Equal21(\CU|Equal2~1_combout ),
	.Equal01(\CU|Equal0~1_combout ),
	.ifid_ifnext_pc_o_1(\IFID|ifid_if.next_pc_o [1]),
	.Equal5(\CU|Equal5~0_combout ),
	.ifid_ifnext_pc_o_0(\IFID|ifid_if.next_pc_o [0]),
	.ifid_ifnext_pc_o_3(\IFID|ifid_if.next_pc_o [3]),
	.ifid_ifnext_pc_o_2(\IFID|ifid_if.next_pc_o [2]),
	.ifid_ifnext_pc_o_5(\IFID|ifid_if.next_pc_o [5]),
	.ifid_ifnext_pc_o_4(\IFID|ifid_if.next_pc_o [4]),
	.ifid_ifnext_pc_o_7(\IFID|ifid_if.next_pc_o [7]),
	.ifid_ifnext_pc_o_6(\IFID|ifid_if.next_pc_o [6]),
	.ifid_ifnext_pc_o_9(\IFID|ifid_if.next_pc_o [9]),
	.ifid_ifnext_pc_o_8(\IFID|ifid_if.next_pc_o [8]),
	.ifid_ifnext_pc_o_11(\IFID|ifid_if.next_pc_o [11]),
	.ifid_ifnext_pc_o_10(\IFID|ifid_if.next_pc_o [10]),
	.ifid_ifnext_pc_o_13(\IFID|ifid_if.next_pc_o [13]),
	.ifid_ifnext_pc_o_12(\IFID|ifid_if.next_pc_o [12]),
	.ifid_ifnext_pc_o_15(\IFID|ifid_if.next_pc_o [15]),
	.ifid_ifnext_pc_o_14(\IFID|ifid_if.next_pc_o [14]),
	.ifid_ifnext_pc_o_17(\IFID|ifid_if.next_pc_o [17]),
	.ifid_ifnext_pc_o_16(\IFID|ifid_if.next_pc_o [16]),
	.ifid_ifnext_pc_o_19(\IFID|ifid_if.next_pc_o [19]),
	.ifid_ifnext_pc_o_18(\IFID|ifid_if.next_pc_o [18]),
	.ifid_ifnext_pc_o_21(\IFID|ifid_if.next_pc_o [21]),
	.ifid_ifnext_pc_o_20(\IFID|ifid_if.next_pc_o [20]),
	.ifid_ifnext_pc_o_23(\IFID|ifid_if.next_pc_o [23]),
	.ifid_ifnext_pc_o_22(\IFID|ifid_if.next_pc_o [22]),
	.ifid_ifnext_pc_o_25(\IFID|ifid_if.next_pc_o [25]),
	.ifid_ifnext_pc_o_24(\IFID|ifid_if.next_pc_o [24]),
	.ifid_ifnext_pc_o_27(\IFID|ifid_if.next_pc_o [27]),
	.ifid_ifnext_pc_o_26(\IFID|ifid_if.next_pc_o [26]),
	.ifid_ifnext_pc_o_29(\IFID|ifid_if.next_pc_o [29]),
	.ifid_ifnext_pc_o_28(\IFID|ifid_if.next_pc_o [28]),
	.ifid_ifnext_pc_o_31(\IFID|ifid_if.next_pc_o [31]),
	.ifid_ifnext_pc_o_30(\IFID|ifid_if.next_pc_o [30]),
	.cuifregWEN1(\CU|cuif.regWEN~5_combout ),
	.Equal1(\CU|Equal1~0_combout ),
	.CPUCLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

if_id IFID(
	.nextpc_2(\nextpc[2]~0_combout ),
	.nextpc_3(\nextpc[3]~2_combout ),
	.nextpc_4(\nextpc[4]~4_combout ),
	.nextpc_5(\nextpc[5]~6_combout ),
	.nextpc_6(\nextpc[6]~8_combout ),
	.nextpc_7(\nextpc[7]~10_combout ),
	.nextpc_8(\nextpc[8]~12_combout ),
	.nextpc_9(\nextpc[9]~14_combout ),
	.nextpc_10(\nextpc[10]~16_combout ),
	.nextpc_11(\nextpc[11]~18_combout ),
	.nextpc_12(\nextpc[12]~20_combout ),
	.nextpc_13(\nextpc[13]~22_combout ),
	.nextpc_14(\nextpc[14]~24_combout ),
	.nextpc_15(\nextpc[15]~26_combout ),
	.nextpc_16(\nextpc[16]~28_combout ),
	.nextpc_17(\nextpc[17]~30_combout ),
	.nextpc_18(\nextpc[18]~32_combout ),
	.nextpc_19(\nextpc[19]~34_combout ),
	.nextpc_20(\nextpc[20]~36_combout ),
	.nextpc_21(\nextpc[21]~38_combout ),
	.nextpc_22(\nextpc[22]~40_combout ),
	.nextpc_23(\nextpc[23]~42_combout ),
	.nextpc_24(\nextpc[24]~44_combout ),
	.nextpc_25(\nextpc[25]~46_combout ),
	.nextpc_26(\nextpc[26]~48_combout ),
	.nextpc_27(\nextpc[27]~50_combout ),
	.nextpc_28(\nextpc[28]~52_combout ),
	.nextpc_29(\nextpc[29]~54_combout ),
	.nextpc_30(\nextpc[30]~56_combout ),
	.nextpc_31(\nextpc[31]~58_combout ),
	.ramiframload_0(ramiframload_0),
	.pc_1(pc_1),
	.pc_0(pc_0),
	.ramiframload_1(ramiframload_1),
	.always1(always11),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_111),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.always11(always13),
	.ifid_ifinstr_o_17(\IFID|ifid_if.instr_o [17]),
	.ifid_ifinstr_o_16(\IFID|ifid_if.instr_o [16]),
	.ifid_ifinstr_o_19(\IFID|ifid_if.instr_o [19]),
	.ifid_ifinstr_o_18(\IFID|ifid_if.instr_o [18]),
	.ifid_ifinstr_o_20(\IFID|ifid_if.instr_o [20]),
	.ifid_ifinstr_o_22(\IFID|ifid_if.instr_o [22]),
	.ifid_ifinstr_o_21(\IFID|ifid_if.instr_o [21]),
	.ifid_ifinstr_o_24(\IFID|ifid_if.instr_o [24]),
	.ifid_ifinstr_o_23(\IFID|ifid_if.instr_o [23]),
	.ifid_ifinstr_o_25(\IFID|ifid_if.instr_o [25]),
	.huiffreeze(\HU|huif.freeze~2_combout ),
	.huifflush(\HU|huif.flush~0_combout ),
	.ifid_ifinstr_o_26(\IFID|ifid_if.instr_o [26]),
	.ifid_ifinstr_o_31(\IFID|ifid_if.instr_o [31]),
	.ifid_ifinstr_o_27(\IFID|ifid_if.instr_o [27]),
	.ifid_ifinstr_o_28(\IFID|ifid_if.instr_o [28]),
	.ifid_ifinstr_o_30(\IFID|ifid_if.instr_o [30]),
	.ifid_ifinstr_o_5(\IFID|ifid_if.instr_o [5]),
	.ifid_ifinstr_o_4(\IFID|ifid_if.instr_o [4]),
	.ifid_ifinstr_o_29(\IFID|ifid_if.instr_o [29]),
	.ifid_ifinstr_o_1(\IFID|ifid_if.instr_o [1]),
	.ifid_ifinstr_o_3(\IFID|ifid_if.instr_o [3]),
	.ifid_ifinstr_o_2(\IFID|ifid_if.instr_o [2]),
	.ifid_ifinstr_o_0(\IFID|ifid_if.instr_o [0]),
	.ifid_ifinstr_o_7(\IFID|ifid_if.instr_o [7]),
	.ifid_ifinstr_o_6(\IFID|ifid_if.instr_o [6]),
	.ifid_ifinstr_o_8(\IFID|ifid_if.instr_o [8]),
	.ifid_ifinstr_o_9(\IFID|ifid_if.instr_o [9]),
	.ifid_ifinstr_o_10(\IFID|ifid_if.instr_o [10]),
	.ifid_ifinstr_o_15(\IFID|ifid_if.instr_o [15]),
	.ifid_ifinstr_o_14(\IFID|ifid_if.instr_o [14]),
	.ifid_ifinstr_o_11(\IFID|ifid_if.instr_o [11]),
	.ifid_ifinstr_o_12(\IFID|ifid_if.instr_o [12]),
	.ifid_ifinstr_o_13(\IFID|ifid_if.instr_o [13]),
	.ifid_ifnext_pc_o_1(\IFID|ifid_if.next_pc_o [1]),
	.ifid_ifnext_pc_o_0(\IFID|ifid_if.next_pc_o [0]),
	.ifid_ifnext_pc_o_3(\IFID|ifid_if.next_pc_o [3]),
	.ifid_ifnext_pc_o_2(\IFID|ifid_if.next_pc_o [2]),
	.ifid_ifnext_pc_o_5(\IFID|ifid_if.next_pc_o [5]),
	.ifid_ifnext_pc_o_4(\IFID|ifid_if.next_pc_o [4]),
	.ifid_ifnext_pc_o_7(\IFID|ifid_if.next_pc_o [7]),
	.ifid_ifnext_pc_o_6(\IFID|ifid_if.next_pc_o [6]),
	.ifid_ifnext_pc_o_9(\IFID|ifid_if.next_pc_o [9]),
	.ifid_ifnext_pc_o_8(\IFID|ifid_if.next_pc_o [8]),
	.ifid_ifnext_pc_o_11(\IFID|ifid_if.next_pc_o [11]),
	.ifid_ifnext_pc_o_10(\IFID|ifid_if.next_pc_o [10]),
	.ifid_ifnext_pc_o_13(\IFID|ifid_if.next_pc_o [13]),
	.ifid_ifnext_pc_o_12(\IFID|ifid_if.next_pc_o [12]),
	.ifid_ifnext_pc_o_15(\IFID|ifid_if.next_pc_o [15]),
	.ifid_ifnext_pc_o_14(\IFID|ifid_if.next_pc_o [14]),
	.ifid_ifnext_pc_o_17(\IFID|ifid_if.next_pc_o [17]),
	.ifid_ifnext_pc_o_16(\IFID|ifid_if.next_pc_o [16]),
	.ifid_ifnext_pc_o_19(\IFID|ifid_if.next_pc_o [19]),
	.ifid_ifnext_pc_o_18(\IFID|ifid_if.next_pc_o [18]),
	.ifid_ifnext_pc_o_21(\IFID|ifid_if.next_pc_o [21]),
	.ifid_ifnext_pc_o_20(\IFID|ifid_if.next_pc_o [20]),
	.ifid_ifnext_pc_o_23(\IFID|ifid_if.next_pc_o [23]),
	.ifid_ifnext_pc_o_22(\IFID|ifid_if.next_pc_o [22]),
	.ifid_ifnext_pc_o_25(\IFID|ifid_if.next_pc_o [25]),
	.ifid_ifnext_pc_o_24(\IFID|ifid_if.next_pc_o [24]),
	.ifid_ifnext_pc_o_27(\IFID|ifid_if.next_pc_o [27]),
	.ifid_ifnext_pc_o_26(\IFID|ifid_if.next_pc_o [26]),
	.ifid_ifnext_pc_o_29(\IFID|ifid_if.next_pc_o [29]),
	.ifid_ifnext_pc_o_28(\IFID|ifid_if.next_pc_o [28]),
	.ifid_ifnext_pc_o_31(\IFID|ifid_if.next_pc_o [31]),
	.ifid_ifnext_pc_o_30(\IFID|ifid_if.next_pc_o [30]),
	.CPUCLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

control_unit CU(
	.ifid_ifinstr_o_26(\IFID|ifid_if.instr_o [26]),
	.ifid_ifinstr_o_31(\IFID|ifid_if.instr_o [31]),
	.ifid_ifinstr_o_27(\IFID|ifid_if.instr_o [27]),
	.ifid_ifinstr_o_28(\IFID|ifid_if.instr_o [28]),
	.ifid_ifinstr_o_30(\IFID|ifid_if.instr_o [30]),
	.ifid_ifinstr_o_5(\IFID|ifid_if.instr_o [5]),
	.ifid_ifinstr_o_4(\IFID|ifid_if.instr_o [4]),
	.always0(\CU|always0~0_combout ),
	.ifid_ifinstr_o_29(\IFID|ifid_if.instr_o [29]),
	.ifid_ifinstr_o_1(\IFID|ifid_if.instr_o [1]),
	.ifid_ifinstr_o_3(\IFID|ifid_if.instr_o [3]),
	.ifid_ifinstr_o_2(\IFID|ifid_if.instr_o [2]),
	.cuifregWEN(\CU|cuif.regWEN~0_combout ),
	.Equal0(\CU|Equal0~0_combout ),
	.ifid_ifinstr_o_0(\IFID|ifid_if.instr_o [0]),
	.Equal3(\CU|Equal3~0_combout ),
	.Equal2(\CU|Equal2~0_combout ),
	.Equal10(\CU|Equal10~0_combout ),
	.Equal14(\CU|Equal14~0_combout ),
	.Equal21(\CU|Equal2~1_combout ),
	.Equal01(\CU|Equal0~1_combout ),
	.Equal5(\CU|Equal5~0_combout ),
	.cuifregWEN1(\CU|cuif.regWEN~5_combout ),
	.Equal1(\CU|Equal1~0_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

register_file RF(
	.rwWB(\rwWB~0_combout ),
	.rwWB1(\rwWB~1_combout ),
	.rwWB2(\rwWB~2_combout ),
	.rwWB3(\rwWB~3_combout ),
	.memwb_ifregWEN_o(\MEMWB|memwb_if.regWEN_o~q ),
	.rwWB4(\rwWB~4_combout ),
	.wdat(\wdat~1_combout ),
	.wdat1(\wdat~3_combout ),
	.wdat2(\wdat~5_combout ),
	.wdat3(\wdat~7_combout ),
	.wdat4(\wdat~9_combout ),
	.wdat5(\wdat~11_combout ),
	.wdat6(\wdat~13_combout ),
	.wdat7(\wdat~15_combout ),
	.wdat8(\wdat~17_combout ),
	.wdat9(\wdat~21_combout ),
	.wdat10(\wdat~23_combout ),
	.wdat11(\wdat~25_combout ),
	.wdat12(\wdat~27_combout ),
	.wdat13(\wdat~29_combout ),
	.wdat14(\wdat~31_combout ),
	.wdat15(\wdat~33_combout ),
	.wdat16(\wdat~35_combout ),
	.wdat17(\wdat~37_combout ),
	.wdat18(\wdat~39_combout ),
	.wdat19(\wdat~41_combout ),
	.wdat20(\wdat~43_combout ),
	.wdat21(\wdat~45_combout ),
	.wdat22(\wdat~47_combout ),
	.wdat23(\wdat~49_combout ),
	.wdat24(\wdat~51_combout ),
	.wdat25(\wdat~53_combout ),
	.wdat26(\wdat~55_combout ),
	.wdat27(\wdat~57_combout ),
	.wdat28(\wdat~59_combout ),
	.wdat29(\wdat~61_combout ),
	.wdat30(\wdat~63_combout ),
	.wdat31(\wdat~65_combout ),
	.ifid_ifinstr_o_17(\IFID|ifid_if.instr_o [17]),
	.ifid_ifinstr_o_16(\IFID|ifid_if.instr_o [16]),
	.ifid_ifinstr_o_19(\IFID|ifid_if.instr_o [19]),
	.ifid_ifinstr_o_18(\IFID|ifid_if.instr_o [18]),
	.ifid_ifinstr_o_22(\IFID|ifid_if.instr_o [22]),
	.ifid_ifinstr_o_21(\IFID|ifid_if.instr_o [21]),
	.ifid_ifinstr_o_24(\IFID|ifid_if.instr_o [24]),
	.ifid_ifinstr_o_23(\IFID|ifid_if.instr_o [23]),
	.Mux62(\RF|Mux62~9_combout ),
	.Mux621(\RF|Mux62~19_combout ),
	.Mux30(\RF|Mux30~9_combout ),
	.Mux301(\RF|Mux30~19_combout ),
	.Mux63(\RF|Mux63~9_combout ),
	.Mux631(\RF|Mux63~19_combout ),
	.Mux31(\RF|Mux31~9_combout ),
	.Mux311(\RF|Mux31~19_combout ),
	.Mux29(\RF|Mux29~9_combout ),
	.Mux291(\RF|Mux29~19_combout ),
	.Mux27(\RF|Mux27~9_combout ),
	.Mux271(\RF|Mux27~19_combout ),
	.Mux28(\RF|Mux28~9_combout ),
	.Mux281(\RF|Mux28~19_combout ),
	.Mux61(\RF|Mux61~9_combout ),
	.Mux611(\RF|Mux61~19_combout ),
	.Mux23(\RF|Mux23~9_combout ),
	.Mux231(\RF|Mux23~19_combout ),
	.Mux24(\RF|Mux24~9_combout ),
	.Mux241(\RF|Mux24~19_combout ),
	.Mux25(\RF|Mux25~9_combout ),
	.Mux251(\RF|Mux25~19_combout ),
	.Mux26(\RF|Mux26~9_combout ),
	.Mux261(\RF|Mux26~19_combout ),
	.Mux60(\RF|Mux60~9_combout ),
	.Mux601(\RF|Mux60~19_combout ),
	.Mux15(\RF|Mux15~9_combout ),
	.Mux151(\RF|Mux15~19_combout ),
	.Mux16(\RF|Mux16~9_combout ),
	.Mux161(\RF|Mux16~19_combout ),
	.Mux17(\RF|Mux17~9_combout ),
	.Mux171(\RF|Mux17~19_combout ),
	.Mux18(\RF|Mux18~9_combout ),
	.Mux181(\RF|Mux18~19_combout ),
	.Mux19(\RF|Mux19~9_combout ),
	.Mux191(\RF|Mux19~19_combout ),
	.Mux20(\RF|Mux20~9_combout ),
	.Mux201(\RF|Mux20~19_combout ),
	.Mux21(\RF|Mux21~9_combout ),
	.Mux211(\RF|Mux21~19_combout ),
	.Mux22(\RF|Mux22~9_combout ),
	.Mux221(\RF|Mux22~19_combout ),
	.Mux59(\RF|Mux59~9_combout ),
	.Mux591(\RF|Mux59~19_combout ),
	.Mux0(\RF|Mux0~9_combout ),
	.Mux01(\RF|Mux0~19_combout ),
	.Mux2(\RF|Mux2~9_combout ),
	.Mux210(\RF|Mux2~19_combout ),
	.Mux1(\RF|Mux1~9_combout ),
	.Mux11(\RF|Mux1~19_combout ),
	.Mux3(\RF|Mux3~9_combout ),
	.Mux32(\RF|Mux3~19_combout ),
	.Mux5(\RF|Mux5~9_combout ),
	.Mux51(\RF|Mux5~19_combout ),
	.Mux4(\RF|Mux4~9_combout ),
	.Mux41(\RF|Mux4~19_combout ),
	.Mux6(\RF|Mux6~9_combout ),
	.Mux64(\RF|Mux6~19_combout ),
	.Mux7(\RF|Mux7~9_combout ),
	.Mux71(\RF|Mux7~19_combout ),
	.Mux9(\RF|Mux9~9_combout ),
	.Mux91(\RF|Mux9~19_combout ),
	.Mux8(\RF|Mux8~9_combout ),
	.Mux81(\RF|Mux8~19_combout ),
	.Mux10(\RF|Mux10~9_combout ),
	.Mux101(\RF|Mux10~19_combout ),
	.Mux111(\RF|Mux11~9_combout ),
	.Mux112(\RF|Mux11~19_combout ),
	.Mux13(\RF|Mux13~9_combout ),
	.Mux131(\RF|Mux13~19_combout ),
	.Mux12(\RF|Mux12~9_combout ),
	.Mux121(\RF|Mux12~19_combout ),
	.Mux14(\RF|Mux14~9_combout ),
	.Mux141(\RF|Mux14~19_combout ),
	.Mux321(\RF|Mux32~9_combout ),
	.Mux322(\RF|Mux32~19_combout ),
	.Mux47(\RF|Mux47~9_combout ),
	.Mux471(\RF|Mux47~19_combout ),
	.Mux46(\RF|Mux46~9_combout ),
	.Mux461(\RF|Mux46~19_combout ),
	.Mux45(\RF|Mux45~9_combout ),
	.Mux451(\RF|Mux45~19_combout ),
	.Mux44(\RF|Mux44~9_combout ),
	.Mux441(\RF|Mux44~19_combout ),
	.Mux43(\RF|Mux43~9_combout ),
	.Mux431(\RF|Mux43~19_combout ),
	.Mux42(\RF|Mux42~9_combout ),
	.Mux421(\RF|Mux42~19_combout ),
	.Mux411(\RF|Mux41~9_combout ),
	.Mux412(\RF|Mux41~19_combout ),
	.Mux40(\RF|Mux40~9_combout ),
	.Mux401(\RF|Mux40~19_combout ),
	.Mux39(\RF|Mux39~9_combout ),
	.Mux391(\RF|Mux39~19_combout ),
	.Mux38(\RF|Mux38~9_combout ),
	.Mux381(\RF|Mux38~19_combout ),
	.Mux37(\RF|Mux37~9_combout ),
	.Mux371(\RF|Mux37~19_combout ),
	.Mux58(\RF|Mux58~9_combout ),
	.Mux581(\RF|Mux58~19_combout ),
	.Mux57(\RF|Mux57~9_combout ),
	.Mux571(\RF|Mux57~19_combout ),
	.Mux56(\RF|Mux56~9_combout ),
	.Mux561(\RF|Mux56~19_combout ),
	.Mux55(\RF|Mux55~9_combout ),
	.Mux551(\RF|Mux55~19_combout ),
	.Mux36(\RF|Mux36~9_combout ),
	.Mux361(\RF|Mux36~19_combout ),
	.Mux35(\RF|Mux35~9_combout ),
	.Mux351(\RF|Mux35~19_combout ),
	.Mux34(\RF|Mux34~9_combout ),
	.Mux341(\RF|Mux34~19_combout ),
	.Mux33(\RF|Mux33~9_combout ),
	.Mux331(\RF|Mux33~19_combout ),
	.Mux54(\RF|Mux54~9_combout ),
	.Mux541(\RF|Mux54~19_combout ),
	.Mux49(\RF|Mux49~9_combout ),
	.Mux491(\RF|Mux49~19_combout ),
	.Mux48(\RF|Mux48~9_combout ),
	.Mux481(\RF|Mux48~19_combout ),
	.Mux53(\RF|Mux53~9_combout ),
	.Mux531(\RF|Mux53~19_combout ),
	.Mux52(\RF|Mux52~9_combout ),
	.Mux521(\RF|Mux52~19_combout ),
	.Mux511(\RF|Mux51~9_combout ),
	.Mux512(\RF|Mux51~19_combout ),
	.Mux50(\RF|Mux50~9_combout ),
	.Mux501(\RF|Mux50~19_combout ),
	.CLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

alu_file ALU(
	.idex_ifaluop_o_1(\IDEX|idex_if.aluop_o [1]),
	.port_b(\port_b~0_combout ),
	.fuifrtReplace_1(\FU|fuif.rtReplace[1]~4_combout ),
	.port_b1(\port_b~3_combout ),
	.always0(\FU|always0~15_combout ),
	.rdat1_1(\rdat1[1]~1_combout ),
	.port_b2(\port_b~4_combout ),
	.port_b3(\port_b~6_combout ),
	.fuifrtReplace_0(\FU|fuif.rtReplace[0]~5_combout ),
	.port_b4(\port_b~7_combout ),
	.rdat1_0(\rdat1[0]~3_combout ),
	.idex_ifaluop_o_2(\IDEX|idex_if.aluop_o [2]),
	.rdat1_2(\rdat1[2]~5_combout ),
	.rdat1_4(\rdat1[4]~6_combout ),
	.mem_data(\mem_data~10_combout ),
	.rdat1_41(\rdat1[4]~7_combout ),
	.rdat1_3(\rdat1[3]~8_combout ),
	.mem_data1(\mem_data~12_combout ),
	.rdat1_31(\rdat1[3]~9_combout ),
	.port_b5(\port_b~9_combout ),
	.fuifrtReplace_2(\FU|fuif.rtReplace[2]~6_combout ),
	.port_b6(\port_b~10_combout ),
	.rdat1_8(\rdat1[8]~11_combout ),
	.rdat1_7(\rdat1[7]~13_combout ),
	.rdat1_6(\rdat1[6]~15_combout ),
	.rdat1_5(\rdat1[5]~17_combout ),
	.port_b7(\port_b~14_combout ),
	.rdat1_16(\rdat1[16]~19_combout ),
	.rdat1_15(\rdat1[15]~21_combout ),
	.rdat1_14(\rdat1[14]~23_combout ),
	.rdat1_13(\rdat1[13]~25_combout ),
	.rdat1_12(\rdat1[12]~27_combout ),
	.rdat1_11(\rdat1[11]~29_combout ),
	.rdat1_10(\rdat1[10]~31_combout ),
	.rdat1_9(\rdat1[9]~33_combout ),
	.port_b8(\port_b~17_combout ),
	.rdat1_311(\rdat1[31]~35_combout ),
	.rdat1_29(\rdat1[29]~37_combout ),
	.rdat1_30(\rdat1[30]~39_combout ),
	.rdat1_28(\rdat1[28]~41_combout ),
	.rdat1_26(\rdat1[26]~43_combout ),
	.rdat1_27(\rdat1[27]~45_combout ),
	.rdat1_25(\rdat1[25]~47_combout ),
	.rdat1_24(\rdat1[24]~49_combout ),
	.rdat1_22(\rdat1[22]~51_combout ),
	.rdat1_23(\rdat1[23]~53_combout ),
	.rdat1_21(\rdat1[21]~55_combout ),
	.rdat1_20(\rdat1[20]~57_combout ),
	.rdat1_18(\rdat1[18]~59_combout ),
	.rdat1_19(\rdat1[19]~61_combout ),
	.rdat1_17(\rdat1[17]~63_combout ),
	.port_b9(\port_b~19_combout ),
	.fuifrtReplace_31(\FU|fuif.rtReplace[31]~9_combout ),
	.port_b10(\port_b~20_combout ),
	.port_b11(\port_b~21_combout ),
	.fuifrtReplace_16(\FU|fuif.rtReplace[16]~10_combout ),
	.port_b12(\port_b~22_combout ),
	.port_b13(\port_b~23_combout ),
	.fuifrtReplace_17(\FU|fuif.rtReplace[17]~11_combout ),
	.port_b14(\port_b~24_combout ),
	.port_b15(\port_b~25_combout ),
	.fuifrtReplace_18(\FU|fuif.rtReplace[18]~12_combout ),
	.port_b16(\port_b~26_combout ),
	.port_b17(\port_b~27_combout ),
	.fuifrtReplace_19(\FU|fuif.rtReplace[19]~13_combout ),
	.port_b18(\port_b~28_combout ),
	.port_b19(\port_b~29_combout ),
	.fuifrtReplace_20(\FU|fuif.rtReplace[20]~14_combout ),
	.port_b20(\port_b~30_combout ),
	.port_b21(\port_b~31_combout ),
	.fuifrtReplace_21(\FU|fuif.rtReplace[21]~15_combout ),
	.port_b22(\port_b~32_combout ),
	.port_b23(\port_b~33_combout ),
	.fuifrtReplace_22(\FU|fuif.rtReplace[22]~16_combout ),
	.port_b24(\port_b~34_combout ),
	.port_b25(\port_b~35_combout ),
	.fuifrtReplace_23(\FU|fuif.rtReplace[23]~17_combout ),
	.port_b26(\port_b~36_combout ),
	.port_b27(\port_b~37_combout ),
	.fuifrtReplace_24(\FU|fuif.rtReplace[24]~18_combout ),
	.port_b28(\port_b~38_combout ),
	.port_b29(\port_b~39_combout ),
	.fuifrtReplace_25(\FU|fuif.rtReplace[25]~19_combout ),
	.port_b30(\port_b~40_combout ),
	.port_b31(\port_b~41_combout ),
	.fuifrtReplace_26(\FU|fuif.rtReplace[26]~20_combout ),
	.port_b32(\port_b~42_combout ),
	.port_b33(\port_b~43_combout ),
	.fuifrtReplace_5(\FU|fuif.rtReplace[5]~21_combout ),
	.port_b34(\port_b~44_combout ),
	.port_b35(\port_b~45_combout ),
	.fuifrtReplace_6(\FU|fuif.rtReplace[6]~22_combout ),
	.port_b36(\port_b~46_combout ),
	.port_b37(\port_b~47_combout ),
	.fuifrtReplace_7(\FU|fuif.rtReplace[7]~23_combout ),
	.port_b38(\port_b~48_combout ),
	.port_b39(\port_b~49_combout ),
	.fuifrtReplace_8(\FU|fuif.rtReplace[8]~24_combout ),
	.port_b40(\port_b~50_combout ),
	.port_b41(\port_b~51_combout ),
	.fuifrtReplace_27(\FU|fuif.rtReplace[27]~25_combout ),
	.port_b42(\port_b~52_combout ),
	.port_b43(\port_b~53_combout ),
	.fuifrtReplace_28(\FU|fuif.rtReplace[28]~26_combout ),
	.port_b44(\port_b~54_combout ),
	.port_b45(\port_b~55_combout ),
	.fuifrtReplace_29(\FU|fuif.rtReplace[29]~27_combout ),
	.port_b46(\port_b~56_combout ),
	.port_b47(\port_b~57_combout ),
	.fuifrtReplace_30(\FU|fuif.rtReplace[30]~28_combout ),
	.port_b48(\port_b~58_combout ),
	.port_b49(\port_b~59_combout ),
	.fuifrtReplace_9(\FU|fuif.rtReplace[9]~29_combout ),
	.port_b50(\port_b~60_combout ),
	.port_b51(\port_b~61_combout ),
	.fuifrtReplace_14(\FU|fuif.rtReplace[14]~30_combout ),
	.port_b52(\port_b~62_combout ),
	.fuifrtReplace_15(\FU|fuif.rtReplace[15]~31_combout ),
	.port_b53(\port_b~63_combout ),
	.port_b54(\port_b~64_combout ),
	.fuifrtReplace_10(\FU|fuif.rtReplace[10]~32_combout ),
	.port_b55(\port_b~65_combout ),
	.port_b56(\port_b~66_combout ),
	.fuifrtReplace_11(\FU|fuif.rtReplace[11]~33_combout ),
	.port_b57(\port_b~67_combout ),
	.port_b58(\port_b~68_combout ),
	.fuifrtReplace_12(\FU|fuif.rtReplace[12]~34_combout ),
	.port_b59(\port_b~69_combout ),
	.fuifrtReplace_13(\FU|fuif.rtReplace[13]~35_combout ),
	.port_b60(\port_b~70_combout ),
	.idex_ifaluop_o_0(\IDEX|idex_if.aluop_o [0]),
	.idex_ifaluop_o_3(\IDEX|idex_if.aluop_o [3]),
	.myifout_1(\ALU|myif.out[1]~15_combout ),
	.myifout_6(\ALU|myif.out[6]~26_combout ),
	.myifout_4(\ALU|myif.out[4]~33_combout ),
	.port_b61(\port_b~71_combout ),
	.port_b62(\port_b~72_combout ),
	.myifout_24(\ALU|myif.out[24]~40_combout ),
	.myifout_26(\ALU|myif.out[26]~47_combout ),
	.myifout_25(\ALU|myif.out[25]~54_combout ),
	.myifout_27(\ALU|myif.out[27]~61_combout ),
	.myifout_5(\ALU|myif.out[5]~68_combout ),
	.myifout_7(\ALU|myif.out[7]~81_combout ),
	.myifout_13(\ALU|myif.out[13]~92_combout ),
	.myifout_9(\ALU|myif.out[9]~98_combout ),
	.myifout_8(\ALU|myif.out[8]~104_combout ),
	.myifout_14(\ALU|myif.out[14]~110_combout ),
	.myifout_12(\ALU|myif.out[12]~116_combout ),
	.myifout_15(\ALU|myif.out[15]~122_combout ),
	.myifout_10(\ALU|myif.out[10]~128_combout ),
	.myifout_11(\ALU|myif.out[11]~134_combout ),
	.myifout_23(\ALU|myif.out[23]~152_combout ),
	.myifout_16(\ALU|myif.out[16]~158_combout ),
	.myifout_17(\ALU|myif.out[17]~174_combout ),
	.myifout_18(\ALU|myif.out[18]~180_combout ),
	.myifout_19(\ALU|myif.out[19]~196_combout ),
	.myifout_30(\ALU|myif.out[30]~204_combout ),
	.myifout_21(\ALU|myif.out[21]~220_combout ),
	.myifnegative(\ALU|myif.negative~8_combout ),
	.myifout_22(\ALU|myif.out[22]~226_combout ),
	.myifout_20(\ALU|myif.out[20]~232_combout ),
	.myifout_0(\ALU|myif.out[0]~239_combout ),
	.Equal10(\ALU|Equal10~10_combout ),
	.myifout_28(\ALU|myif.out[28]~252_combout ),
	.myifout_29(\ALU|myif.out[29]~264_combout ),
	.myifout_2(\ALU|myif.out[2]~274_combout ),
	.myifout_3(\ALU|myif.out[3]~283_combout ),
	.myifout_31(\ALU|myif.out[3]~285_combout ),
	.myifout_210(\ALU|myif.out[2]~289_combout ),
	.Equal101(\ALU|Equal10~12_combout ),
	.myifout_32(\ALU|myif.out[3]~291_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

forward_unit FU(
	.idex_ifrt_o_0(\IDEX|idex_if.rt_o [0]),
	.idex_ifrt_o_1(\IDEX|idex_if.rt_o [1]),
	.rwMEM(\rwMEM~0_combout ),
	.rwMEM1(\rwMEM~1_combout ),
	.idex_ifrt_o_2(\IDEX|idex_if.rt_o [2]),
	.idex_ifrt_o_3(\IDEX|idex_if.rt_o [3]),
	.rwMEM2(\rwMEM~2_combout ),
	.rwMEM3(\rwMEM~3_combout ),
	.exmem_ifregWEN_o(\EXMEM|exmem_if.regWEN_o~q ),
	.idex_ifrt_o_4(\IDEX|idex_if.rt_o [4]),
	.rwMEM4(\rwMEM~4_combout ),
	.always0(\FU|always0~3_combout ),
	.rwWB(\rwWB~0_combout ),
	.rwWB1(\rwWB~1_combout ),
	.rwWB2(\rwWB~2_combout ),
	.rwWB3(\rwWB~3_combout ),
	.memwb_ifregWEN_o(\MEMWB|memwb_if.regWEN_o~q ),
	.rwWB4(\rwWB~4_combout ),
	.always01(\FU|always0~7_combout ),
	.wdat(\wdat~1_combout ),
	.mem_data(\mem_data~4_combout ),
	.fuifrtReplace_1(\FU|fuif.rtReplace[1]~4_combout ),
	.idex_ifrs_o_1(\IDEX|idex_if.rs_o [1]),
	.idex_ifrs_o_0(\IDEX|idex_if.rs_o [0]),
	.idex_ifrs_o_3(\IDEX|idex_if.rs_o [3]),
	.idex_ifrs_o_2(\IDEX|idex_if.rs_o [2]),
	.idex_ifrs_o_4(\IDEX|idex_if.rs_o [4]),
	.always02(\FU|always0~11_combout ),
	.always03(\FU|always0~15_combout ),
	.mem_data1(\mem_data~6_combout ),
	.wdat1(\wdat~3_combout ),
	.fuifrtReplace_0(\FU|fuif.rtReplace[0]~5_combout ),
	.wdat2(\wdat~5_combout ),
	.mem_data2(\mem_data~8_combout ),
	.wdat3(\wdat~7_combout ),
	.mem_data3(\mem_data~10_combout ),
	.wdat4(\wdat~9_combout ),
	.mem_data4(\mem_data~12_combout ),
	.fuifrtReplace_2(\FU|fuif.rtReplace[2]~6_combout ),
	.wdat5(\wdat~11_combout ),
	.mem_data5(\mem_data~14_combout ),
	.wdat6(\wdat~13_combout ),
	.mem_data6(\mem_data~16_combout ),
	.wdat7(\wdat~15_combout ),
	.mem_data7(\mem_data~18_combout ),
	.wdat8(\wdat~17_combout ),
	.mem_data8(\mem_data~20_combout ),
	.fuifrtReplace_3(\FU|fuif.rtReplace[3]~7_combout ),
	.wdat9(\wdat~21_combout ),
	.mem_data9(\mem_data~24_combout ),
	.wdat10(\wdat~23_combout ),
	.mem_data10(\mem_data~26_combout ),
	.wdat11(\wdat~25_combout ),
	.mem_data11(\mem_data~28_combout ),
	.wdat12(\wdat~27_combout ),
	.mem_data12(\mem_data~30_combout ),
	.wdat13(\wdat~29_combout ),
	.mem_data13(\mem_data~32_combout ),
	.wdat14(\wdat~31_combout ),
	.mem_data14(\mem_data~34_combout ),
	.wdat15(\wdat~33_combout ),
	.mem_data15(\mem_data~36_combout ),
	.wdat16(\wdat~35_combout ),
	.mem_data16(\mem_data~38_combout ),
	.fuifrtReplace_4(\FU|fuif.rtReplace[4]~8_combout ),
	.wdat17(\wdat~37_combout ),
	.mem_data17(\mem_data~40_combout ),
	.wdat18(\wdat~39_combout ),
	.mem_data18(\mem_data~42_combout ),
	.wdat19(\wdat~41_combout ),
	.mem_data19(\mem_data~44_combout ),
	.wdat20(\wdat~43_combout ),
	.mem_data20(\mem_data~46_combout ),
	.wdat21(\wdat~45_combout ),
	.mem_data21(\mem_data~48_combout ),
	.wdat22(\wdat~47_combout ),
	.mem_data22(\mem_data~50_combout ),
	.wdat23(\wdat~49_combout ),
	.mem_data23(\mem_data~52_combout ),
	.wdat24(\wdat~51_combout ),
	.mem_data24(\mem_data~54_combout ),
	.wdat25(\wdat~53_combout ),
	.mem_data25(\mem_data~56_combout ),
	.wdat26(\wdat~55_combout ),
	.mem_data26(\mem_data~58_combout ),
	.wdat27(\wdat~57_combout ),
	.mem_data27(\mem_data~60_combout ),
	.wdat28(\wdat~59_combout ),
	.mem_data28(\mem_data~62_combout ),
	.wdat29(\wdat~61_combout ),
	.mem_data29(\mem_data~64_combout ),
	.wdat30(\wdat~63_combout ),
	.mem_data30(\mem_data~66_combout ),
	.wdat31(\wdat~65_combout ),
	.mem_data31(\mem_data~68_combout ),
	.fuifrtReplace_31(\FU|fuif.rtReplace[31]~9_combout ),
	.fuifrtReplace_16(\FU|fuif.rtReplace[16]~10_combout ),
	.fuifrtReplace_17(\FU|fuif.rtReplace[17]~11_combout ),
	.fuifrtReplace_18(\FU|fuif.rtReplace[18]~12_combout ),
	.fuifrtReplace_19(\FU|fuif.rtReplace[19]~13_combout ),
	.fuifrtReplace_20(\FU|fuif.rtReplace[20]~14_combout ),
	.fuifrtReplace_21(\FU|fuif.rtReplace[21]~15_combout ),
	.fuifrtReplace_22(\FU|fuif.rtReplace[22]~16_combout ),
	.fuifrtReplace_23(\FU|fuif.rtReplace[23]~17_combout ),
	.fuifrtReplace_24(\FU|fuif.rtReplace[24]~18_combout ),
	.fuifrtReplace_25(\FU|fuif.rtReplace[25]~19_combout ),
	.fuifrtReplace_26(\FU|fuif.rtReplace[26]~20_combout ),
	.fuifrtReplace_5(\FU|fuif.rtReplace[5]~21_combout ),
	.fuifrtReplace_6(\FU|fuif.rtReplace[6]~22_combout ),
	.fuifrtReplace_7(\FU|fuif.rtReplace[7]~23_combout ),
	.fuifrtReplace_8(\FU|fuif.rtReplace[8]~24_combout ),
	.fuifrtReplace_27(\FU|fuif.rtReplace[27]~25_combout ),
	.fuifrtReplace_28(\FU|fuif.rtReplace[28]~26_combout ),
	.fuifrtReplace_29(\FU|fuif.rtReplace[29]~27_combout ),
	.fuifrtReplace_30(\FU|fuif.rtReplace[30]~28_combout ),
	.fuifrtReplace_9(\FU|fuif.rtReplace[9]~29_combout ),
	.fuifrtReplace_14(\FU|fuif.rtReplace[14]~30_combout ),
	.fuifrtReplace_15(\FU|fuif.rtReplace[15]~31_combout ),
	.fuifrtReplace_10(\FU|fuif.rtReplace[10]~32_combout ),
	.fuifrtReplace_11(\FU|fuif.rtReplace[11]~33_combout ),
	.fuifrtReplace_12(\FU|fuif.rtReplace[12]~34_combout ),
	.fuifrtReplace_13(\FU|fuif.rtReplace[13]~35_combout ),
	.fuifrdat2_ow(\FU|fuif.rdat2_ow~0_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X52_Y29_N30
cycloneive_lcell_comb \nextpc[16]~28 (
// Equation(s):
// \nextpc[16]~28_combout  = (pc_16 & (\nextpc[15]~27  $ (GND))) # (!pc_16 & (!\nextpc[15]~27  & VCC))
// \nextpc[16]~29  = CARRY((pc_16 & !\nextpc[15]~27 ))

	.dataa(gnd),
	.datab(pc_16),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[15]~27 ),
	.combout(\nextpc[16]~28_combout ),
	.cout(\nextpc[16]~29 ));
// synopsys translate_off
defparam \nextpc[16]~28 .lut_mask = 16'hC30C;
defparam \nextpc[16]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N2
cycloneive_lcell_comb \nextpc[18]~32 (
// Equation(s):
// \nextpc[18]~32_combout  = (pc_18 & (\nextpc[17]~31  $ (GND))) # (!pc_18 & (!\nextpc[17]~31  & VCC))
// \nextpc[18]~33  = CARRY((pc_18 & !\nextpc[17]~31 ))

	.dataa(pc_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[17]~31 ),
	.combout(\nextpc[18]~32_combout ),
	.cout(\nextpc[18]~33 ));
// synopsys translate_off
defparam \nextpc[18]~32 .lut_mask = 16'hA50A;
defparam \nextpc[18]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N14
cycloneive_lcell_comb \nextpc[24]~44 (
// Equation(s):
// \nextpc[24]~44_combout  = (pc_24 & (\nextpc[23]~43  $ (GND))) # (!pc_24 & (!\nextpc[23]~43  & VCC))
// \nextpc[24]~45  = CARRY((pc_24 & !\nextpc[23]~43 ))

	.dataa(gnd),
	.datab(pc_24),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[23]~43 ),
	.combout(\nextpc[24]~44_combout ),
	.cout(\nextpc[24]~45 ));
// synopsys translate_off
defparam \nextpc[24]~44 .lut_mask = 16'hC30C;
defparam \nextpc[24]~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N18
cycloneive_lcell_comb \nextpc[26]~48 (
// Equation(s):
// \nextpc[26]~48_combout  = (pc_26 & (\nextpc[25]~47  $ (GND))) # (!pc_26 & (!\nextpc[25]~47  & VCC))
// \nextpc[26]~49  = CARRY((pc_26 & !\nextpc[25]~47 ))

	.dataa(gnd),
	.datab(pc_26),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[25]~47 ),
	.combout(\nextpc[26]~48_combout ),
	.cout(\nextpc[26]~49 ));
// synopsys translate_off
defparam \nextpc[26]~48 .lut_mask = 16'hC30C;
defparam \nextpc[26]~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N22
cycloneive_lcell_comb \nextpc[28]~52 (
// Equation(s):
// \nextpc[28]~52_combout  = (pc_28 & (\nextpc[27]~51  $ (GND))) # (!pc_28 & (!\nextpc[27]~51  & VCC))
// \nextpc[28]~53  = CARRY((pc_28 & !\nextpc[27]~51 ))

	.dataa(pc_28),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[27]~51 ),
	.combout(\nextpc[28]~52_combout ),
	.cout(\nextpc[28]~53 ));
// synopsys translate_off
defparam \nextpc[28]~52 .lut_mask = 16'hA50A;
defparam \nextpc[28]~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N18
cycloneive_lcell_comb \rwMEM~0 (
// Equation(s):
// \rwMEM~0_combout  = (exmem_ifRegDest_o_1) # ((exmem_ifRegDest_o_0 & (exmem_ifrt_o_1)) # (!exmem_ifRegDest_o_0 & ((exmem_ifrd_o_1))))

	.dataa(\EXMEM|exmem_if.RegDest_o [0]),
	.datab(\EXMEM|exmem_if.rt_o [1]),
	.datac(\EXMEM|exmem_if.rd_o [1]),
	.datad(\EXMEM|exmem_if.RegDest_o [1]),
	.cin(gnd),
	.combout(\rwMEM~0_combout ),
	.cout());
// synopsys translate_off
defparam \rwMEM~0 .lut_mask = 16'hFFD8;
defparam \rwMEM~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N28
cycloneive_lcell_comb \rwMEM~1 (
// Equation(s):
// \rwMEM~1_combout  = (exmem_ifRegDest_o_1) # ((exmem_ifRegDest_o_0 & (exmem_ifrt_o_0)) # (!exmem_ifRegDest_o_0 & ((exmem_ifrd_o_0))))

	.dataa(\EXMEM|exmem_if.RegDest_o [0]),
	.datab(\EXMEM|exmem_if.rt_o [0]),
	.datac(\EXMEM|exmem_if.rd_o [0]),
	.datad(\EXMEM|exmem_if.RegDest_o [1]),
	.cin(gnd),
	.combout(\rwMEM~1_combout ),
	.cout());
// synopsys translate_off
defparam \rwMEM~1 .lut_mask = 16'hFFD8;
defparam \rwMEM~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N14
cycloneive_lcell_comb \rwMEM~2 (
// Equation(s):
// \rwMEM~2_combout  = (exmem_ifRegDest_o_1) # ((exmem_ifRegDest_o_0 & (exmem_ifrt_o_3)) # (!exmem_ifRegDest_o_0 & ((exmem_ifrd_o_3))))

	.dataa(\EXMEM|exmem_if.RegDest_o [0]),
	.datab(\EXMEM|exmem_if.RegDest_o [1]),
	.datac(\EXMEM|exmem_if.rt_o [3]),
	.datad(\EXMEM|exmem_if.rd_o [3]),
	.cin(gnd),
	.combout(\rwMEM~2_combout ),
	.cout());
// synopsys translate_off
defparam \rwMEM~2 .lut_mask = 16'hFDEC;
defparam \rwMEM~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N24
cycloneive_lcell_comb \rwMEM~3 (
// Equation(s):
// \rwMEM~3_combout  = (exmem_ifRegDest_o_1) # ((exmem_ifRegDest_o_0 & ((exmem_ifrt_o_2))) # (!exmem_ifRegDest_o_0 & (exmem_ifrd_o_2)))

	.dataa(\EXMEM|exmem_if.rd_o [2]),
	.datab(\EXMEM|exmem_if.RegDest_o [1]),
	.datac(\EXMEM|exmem_if.rt_o [2]),
	.datad(\EXMEM|exmem_if.RegDest_o [0]),
	.cin(gnd),
	.combout(\rwMEM~3_combout ),
	.cout());
// synopsys translate_off
defparam \rwMEM~3 .lut_mask = 16'hFCEE;
defparam \rwMEM~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N4
cycloneive_lcell_comb \rwMEM~4 (
// Equation(s):
// \rwMEM~4_combout  = (exmem_ifRegDest_o_1) # ((exmem_ifRegDest_o_0 & (exmem_ifrt_o_4)) # (!exmem_ifRegDest_o_0 & ((exmem_ifrd_o_4))))

	.dataa(\EXMEM|exmem_if.rt_o [4]),
	.datab(\EXMEM|exmem_if.RegDest_o [0]),
	.datac(\EXMEM|exmem_if.rd_o [4]),
	.datad(\EXMEM|exmem_if.RegDest_o [1]),
	.cin(gnd),
	.combout(\rwMEM~4_combout ),
	.cout());
// synopsys translate_off
defparam \rwMEM~4 .lut_mask = 16'hFFB8;
defparam \rwMEM~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N16
cycloneive_lcell_comb \rwWB~0 (
// Equation(s):
// \rwWB~0_combout  = (memwb_ifRegDest_o_1) # ((memwb_ifRegDest_o_0 & (memwb_ifrt_o_1)) # (!memwb_ifRegDest_o_0 & ((memwb_ifrd_o_1))))

	.dataa(\MEMWB|memwb_if.RegDest_o [0]),
	.datab(\MEMWB|memwb_if.rt_o [1]),
	.datac(\MEMWB|memwb_if.rd_o [1]),
	.datad(\MEMWB|memwb_if.RegDest_o [1]),
	.cin(gnd),
	.combout(\rwWB~0_combout ),
	.cout());
// synopsys translate_off
defparam \rwWB~0 .lut_mask = 16'hFFD8;
defparam \rwWB~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N14
cycloneive_lcell_comb \rwWB~1 (
// Equation(s):
// \rwWB~1_combout  = (memwb_ifRegDest_o_1) # ((memwb_ifRegDest_o_0 & (memwb_ifrt_o_0)) # (!memwb_ifRegDest_o_0 & ((memwb_ifrd_o_0))))

	.dataa(\MEMWB|memwb_if.RegDest_o [0]),
	.datab(\MEMWB|memwb_if.rt_o [0]),
	.datac(\MEMWB|memwb_if.rd_o [0]),
	.datad(\MEMWB|memwb_if.RegDest_o [1]),
	.cin(gnd),
	.combout(\rwWB~1_combout ),
	.cout());
// synopsys translate_off
defparam \rwWB~1 .lut_mask = 16'hFFD8;
defparam \rwWB~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N10
cycloneive_lcell_comb \rwWB~2 (
// Equation(s):
// \rwWB~2_combout  = (memwb_ifRegDest_o_1) # ((memwb_ifRegDest_o_0 & (memwb_ifrt_o_3)) # (!memwb_ifRegDest_o_0 & ((memwb_ifrd_o_3))))

	.dataa(\MEMWB|memwb_if.RegDest_o [0]),
	.datab(\MEMWB|memwb_if.rt_o [3]),
	.datac(\MEMWB|memwb_if.rd_o [3]),
	.datad(\MEMWB|memwb_if.RegDest_o [1]),
	.cin(gnd),
	.combout(\rwWB~2_combout ),
	.cout());
// synopsys translate_off
defparam \rwWB~2 .lut_mask = 16'hFFD8;
defparam \rwWB~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N6
cycloneive_lcell_comb \rwWB~3 (
// Equation(s):
// \rwWB~3_combout  = (memwb_ifRegDest_o_1) # ((memwb_ifRegDest_o_0 & (memwb_ifrt_o_2)) # (!memwb_ifRegDest_o_0 & ((memwb_ifrd_o_2))))

	.dataa(\MEMWB|memwb_if.rt_o [2]),
	.datab(\MEMWB|memwb_if.RegDest_o [1]),
	.datac(\MEMWB|memwb_if.rd_o [2]),
	.datad(\MEMWB|memwb_if.RegDest_o [0]),
	.cin(gnd),
	.combout(\rwWB~3_combout ),
	.cout());
// synopsys translate_off
defparam \rwWB~3 .lut_mask = 16'hEEFC;
defparam \rwWB~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N2
cycloneive_lcell_comb \rwWB~4 (
// Equation(s):
// \rwWB~4_combout  = (memwb_ifRegDest_o_1) # ((memwb_ifRegDest_o_0 & (memwb_ifrt_o_4)) # (!memwb_ifRegDest_o_0 & ((memwb_ifrd_o_4))))

	.dataa(\MEMWB|memwb_if.RegDest_o [0]),
	.datab(\MEMWB|memwb_if.rt_o [4]),
	.datac(\MEMWB|memwb_if.rd_o [4]),
	.datad(\MEMWB|memwb_if.RegDest_o [1]),
	.cin(gnd),
	.combout(\rwWB~4_combout ),
	.cout());
// synopsys translate_off
defparam \rwWB~4 .lut_mask = 16'hFFD8;
defparam \rwWB~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N20
cycloneive_lcell_comb \port_b~0 (
// Equation(s):
// \port_b~0_combout  = (!idex_ifALUSel_o_1 & (!idex_ifALUSel_o_0 & ((always0) # (always01))))

	.dataa(\IDEX|idex_if.ALUSel_o [1]),
	.datab(\FU|always0~3_combout ),
	.datac(\IDEX|idex_if.ALUSel_o [0]),
	.datad(\FU|always0~7_combout ),
	.cin(gnd),
	.combout(\port_b~0_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~0 .lut_mask = 16'h0504;
defparam \port_b~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N18
cycloneive_lcell_comb \wdat~0 (
// Equation(s):
// \wdat~0_combout  = (!memwb_ifjal_o & ((memwb_ifmemToReg_o & (memwb_ifdmemload_o_1)) # (!memwb_ifmemToReg_o & ((memwb_ifout_o_1)))))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.dmemload_o [1]),
	.datac(\MEMWB|memwb_if.out_o [1]),
	.datad(\MEMWB|memwb_if.memToReg_o~q ),
	.cin(gnd),
	.combout(\wdat~0_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~0 .lut_mask = 16'h4450;
defparam \wdat~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N28
cycloneive_lcell_comb \wdat~1 (
// Equation(s):
// \wdat~1_combout  = (!memwb_iflui_o & ((\wdat~0_combout ) # ((memwb_ifjal_o & memwb_ifnext_pc_o_1))))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.lui_o~q ),
	.datac(\MEMWB|memwb_if.next_pc_o [1]),
	.datad(\wdat~0_combout ),
	.cin(gnd),
	.combout(\wdat~1_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~1 .lut_mask = 16'h3320;
defparam \wdat~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N26
cycloneive_lcell_comb \mem_data~0 (
// Equation(s):
// \mem_data~0_combout  = (!exmem_iflui_o & exmem_ifjal_o)

	.dataa(\EXMEM|exmem_if.lui_o~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\EXMEM|exmem_if.jal_o~q ),
	.cin(gnd),
	.combout(\mem_data~0_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~0 .lut_mask = 16'h5500;
defparam \mem_data~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N2
cycloneive_lcell_comb \mem_data~1 (
// Equation(s):
// \mem_data~1_combout  = (!exmem_iflui_o & (!exmem_ifjal_o & !exmem_ifmemToReg_o))

	.dataa(\EXMEM|exmem_if.lui_o~q ),
	.datab(\EXMEM|exmem_if.jal_o~q ),
	.datac(\EXMEM|exmem_if.memToReg_o~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_data~1_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~1 .lut_mask = 16'h0101;
defparam \mem_data~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N4
cycloneive_lcell_comb \mem_data~2 (
// Equation(s):
// \mem_data~2_combout  = (\mem_data~0_combout  & ((exmem_ifnext_pc_o_1) # ((exmem_ifout_o_1 & \mem_data~1_combout )))) # (!\mem_data~0_combout  & (((exmem_ifout_o_1 & \mem_data~1_combout ))))

	.dataa(\mem_data~0_combout ),
	.datab(\EXMEM|exmem_if.next_pc_o [1]),
	.datac(exmem_ifout_o_1),
	.datad(\mem_data~1_combout ),
	.cin(gnd),
	.combout(\mem_data~2_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~2 .lut_mask = 16'hF888;
defparam \mem_data~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N14
cycloneive_lcell_comb \mem_data~3 (
// Equation(s):
// \mem_data~3_combout  = (!exmem_iflui_o & (!exmem_ifjal_o & exmem_ifmemToReg_o))

	.dataa(\EXMEM|exmem_if.lui_o~q ),
	.datab(\EXMEM|exmem_if.jal_o~q ),
	.datac(gnd),
	.datad(\EXMEM|exmem_if.memToReg_o~q ),
	.cin(gnd),
	.combout(\mem_data~3_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~3 .lut_mask = 16'h1100;
defparam \mem_data~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N2
cycloneive_lcell_comb \mem_data~4 (
// Equation(s):
// \mem_data~4_combout  = (\mem_data~2_combout ) # ((always11 & (\mem_data~3_combout  & ramiframload_1)))

	.dataa(always11),
	.datab(\mem_data~3_combout ),
	.datac(ramiframload_1),
	.datad(\mem_data~2_combout ),
	.cin(gnd),
	.combout(\mem_data~4_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~4 .lut_mask = 16'hFF80;
defparam \mem_data~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N2
cycloneive_lcell_comb \port_b~1 (
// Equation(s):
// \port_b~1_combout  = (idex_ifALUSel_o_1 & (((idex_ifimm_o_1)))) # (!idex_ifALUSel_o_1 & (idex_ifALUSel_o_0 & (idex_ifshamt_o_1)))

	.dataa(\IDEX|idex_if.ALUSel_o [1]),
	.datab(\IDEX|idex_if.ALUSel_o [0]),
	.datac(\IDEX|idex_if.shamt_o [1]),
	.datad(\IDEX|idex_if.imm_o [1]),
	.cin(gnd),
	.combout(\port_b~1_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~1 .lut_mask = 16'hEA40;
defparam \port_b~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N14
cycloneive_lcell_comb \port_b~2 (
// Equation(s):
// \port_b~2_combout  = (!idex_ifALUSel_o_1 & (!always0 & (!idex_ifALUSel_o_0 & !always01)))

	.dataa(\IDEX|idex_if.ALUSel_o [1]),
	.datab(\FU|always0~3_combout ),
	.datac(\IDEX|idex_if.ALUSel_o [0]),
	.datad(\FU|always0~7_combout ),
	.cin(gnd),
	.combout(\port_b~2_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~2 .lut_mask = 16'h0001;
defparam \port_b~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N6
cycloneive_lcell_comb \port_b~3 (
// Equation(s):
// \port_b~3_combout  = (\port_b~1_combout ) # ((idex_ifrdat2_o_1 & \port_b~2_combout ))

	.dataa(gnd),
	.datab(\IDEX|idex_if.rdat2_o [1]),
	.datac(\port_b~2_combout ),
	.datad(\port_b~1_combout ),
	.cin(gnd),
	.combout(\port_b~3_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~3 .lut_mask = 16'hFFC0;
defparam \port_b~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N8
cycloneive_lcell_comb \rdat1[1]~0 (
// Equation(s):
// \rdat1[1]~0_combout  = (!always03 & ((always02 & (\wdat~1_combout )) # (!always02 & ((idex_ifrdat1_o_1)))))

	.dataa(\FU|always0~11_combout ),
	.datab(\FU|always0~15_combout ),
	.datac(\wdat~1_combout ),
	.datad(\IDEX|idex_if.rdat1_o [1]),
	.cin(gnd),
	.combout(\rdat1[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[1]~0 .lut_mask = 16'h3120;
defparam \rdat1[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N24
cycloneive_lcell_comb \rdat1[1]~1 (
// Equation(s):
// \rdat1[1]~1_combout  = (\rdat1[1]~0_combout ) # ((always03 & \mem_data~4_combout ))

	.dataa(\rdat1[1]~0_combout ),
	.datab(gnd),
	.datac(\FU|always0~15_combout ),
	.datad(\mem_data~4_combout ),
	.cin(gnd),
	.combout(\rdat1[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[1]~1 .lut_mask = 16'hFAAA;
defparam \rdat1[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N8
cycloneive_lcell_comb \port_b~4 (
// Equation(s):
// \port_b~4_combout  = (\port_b~3_combout ) # ((\port_b~0_combout  & fuifrtReplace_1))

	.dataa(\port_b~3_combout ),
	.datab(\port_b~0_combout ),
	.datac(gnd),
	.datad(\FU|fuif.rtReplace[1]~4_combout ),
	.cin(gnd),
	.combout(\port_b~4_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~4 .lut_mask = 16'hEEAA;
defparam \port_b~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N0
cycloneive_lcell_comb \port_b~5 (
// Equation(s):
// \port_b~5_combout  = (idex_ifALUSel_o_1 & (((idex_ifimm_o_0)))) # (!idex_ifALUSel_o_1 & (idex_ifALUSel_o_0 & (idex_ifshamt_o_0)))

	.dataa(\IDEX|idex_if.ALUSel_o [1]),
	.datab(\IDEX|idex_if.ALUSel_o [0]),
	.datac(\IDEX|idex_if.shamt_o [0]),
	.datad(\IDEX|idex_if.imm_o [0]),
	.cin(gnd),
	.combout(\port_b~5_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~5 .lut_mask = 16'hEA40;
defparam \port_b~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N14
cycloneive_lcell_comb \port_b~6 (
// Equation(s):
// \port_b~6_combout  = (\port_b~5_combout ) # ((idex_ifrdat2_o_0 & \port_b~2_combout ))

	.dataa(\IDEX|idex_if.rdat2_o [0]),
	.datab(gnd),
	.datac(\port_b~5_combout ),
	.datad(\port_b~2_combout ),
	.cin(gnd),
	.combout(\port_b~6_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~6 .lut_mask = 16'hFAF0;
defparam \port_b~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N12
cycloneive_lcell_comb \mem_data~5 (
// Equation(s):
// \mem_data~5_combout  = (\mem_data~1_combout  & ((exmem_ifout_o_0) # ((\mem_data~0_combout  & exmem_ifnext_pc_o_0)))) # (!\mem_data~1_combout  & (((\mem_data~0_combout  & exmem_ifnext_pc_o_0))))

	.dataa(\mem_data~1_combout ),
	.datab(exmem_ifout_o_0),
	.datac(\mem_data~0_combout ),
	.datad(\EXMEM|exmem_if.next_pc_o [0]),
	.cin(gnd),
	.combout(\mem_data~5_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~5 .lut_mask = 16'hF888;
defparam \mem_data~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N8
cycloneive_lcell_comb \mem_data~6 (
// Equation(s):
// \mem_data~6_combout  = (\mem_data~5_combout ) # ((\mem_data~3_combout  & ((ramiframload_0) # (!always11))))

	.dataa(\mem_data~5_combout ),
	.datab(\mem_data~3_combout ),
	.datac(always11),
	.datad(ramiframload_0),
	.cin(gnd),
	.combout(\mem_data~6_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~6 .lut_mask = 16'hEEAE;
defparam \mem_data~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N18
cycloneive_lcell_comb \wdat~2 (
// Equation(s):
// \wdat~2_combout  = (!memwb_ifjal_o & ((memwb_ifmemToReg_o & (memwb_ifdmemload_o_0)) # (!memwb_ifmemToReg_o & ((memwb_ifout_o_0)))))

	.dataa(\MEMWB|memwb_if.memToReg_o~q ),
	.datab(\MEMWB|memwb_if.dmemload_o [0]),
	.datac(\MEMWB|memwb_if.out_o [0]),
	.datad(\MEMWB|memwb_if.jal_o~q ),
	.cin(gnd),
	.combout(\wdat~2_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~2 .lut_mask = 16'h00D8;
defparam \wdat~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N20
cycloneive_lcell_comb \wdat~3 (
// Equation(s):
// \wdat~3_combout  = (!memwb_iflui_o & ((\wdat~2_combout ) # ((memwb_ifjal_o & memwb_ifnext_pc_o_0))))

	.dataa(\MEMWB|memwb_if.lui_o~q ),
	.datab(\MEMWB|memwb_if.jal_o~q ),
	.datac(\MEMWB|memwb_if.next_pc_o [0]),
	.datad(\wdat~2_combout ),
	.cin(gnd),
	.combout(\wdat~3_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~3 .lut_mask = 16'h5540;
defparam \wdat~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N12
cycloneive_lcell_comb \port_b~7 (
// Equation(s):
// \port_b~7_combout  = (\port_b~6_combout ) # ((\port_b~0_combout  & fuifrtReplace_0))

	.dataa(gnd),
	.datab(\port_b~0_combout ),
	.datac(\port_b~6_combout ),
	.datad(\FU|fuif.rtReplace[0]~5_combout ),
	.cin(gnd),
	.combout(\port_b~7_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~7 .lut_mask = 16'hFCF0;
defparam \port_b~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N2
cycloneive_lcell_comb \rdat1[0]~2 (
// Equation(s):
// \rdat1[0]~2_combout  = (!always03 & ((always02 & ((\wdat~3_combout ))) # (!always02 & (idex_ifrdat1_o_0))))

	.dataa(\FU|always0~11_combout ),
	.datab(\IDEX|idex_if.rdat1_o [0]),
	.datac(\wdat~3_combout ),
	.datad(\FU|always0~15_combout ),
	.cin(gnd),
	.combout(\rdat1[0]~2_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[0]~2 .lut_mask = 16'h00E4;
defparam \rdat1[0]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N16
cycloneive_lcell_comb \rdat1[0]~3 (
// Equation(s):
// \rdat1[0]~3_combout  = (\rdat1[0]~2_combout ) # ((always03 & \mem_data~6_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(gnd),
	.datac(\mem_data~6_combout ),
	.datad(\rdat1[0]~2_combout ),
	.cin(gnd),
	.combout(\rdat1[0]~3_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[0]~3 .lut_mask = 16'hFFA0;
defparam \rdat1[0]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N12
cycloneive_lcell_comb \wdat~4 (
// Equation(s):
// \wdat~4_combout  = (!memwb_ifjal_o & ((memwb_ifmemToReg_o & ((memwb_ifdmemload_o_2))) # (!memwb_ifmemToReg_o & (memwb_ifout_o_2))))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.memToReg_o~q ),
	.datac(\MEMWB|memwb_if.out_o [2]),
	.datad(\MEMWB|memwb_if.dmemload_o [2]),
	.cin(gnd),
	.combout(\wdat~4_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~4 .lut_mask = 16'h5410;
defparam \wdat~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N30
cycloneive_lcell_comb \wdat~5 (
// Equation(s):
// \wdat~5_combout  = (!memwb_iflui_o & ((\wdat~4_combout ) # ((memwb_ifjal_o & memwb_ifnext_pc_o_2))))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.lui_o~q ),
	.datac(\MEMWB|memwb_if.next_pc_o [2]),
	.datad(\wdat~4_combout ),
	.cin(gnd),
	.combout(\wdat~5_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~5 .lut_mask = 16'h3320;
defparam \wdat~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N8
cycloneive_lcell_comb \rdat1[2]~4 (
// Equation(s):
// \rdat1[2]~4_combout  = (!always03 & ((always02 & (\wdat~5_combout )) # (!always02 & ((idex_ifrdat1_o_2)))))

	.dataa(\FU|always0~15_combout ),
	.datab(\wdat~5_combout ),
	.datac(\FU|always0~11_combout ),
	.datad(\IDEX|idex_if.rdat1_o [2]),
	.cin(gnd),
	.combout(\rdat1[2]~4_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[2]~4 .lut_mask = 16'h4540;
defparam \rdat1[2]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N30
cycloneive_lcell_comb \mem_data~7 (
// Equation(s):
// \mem_data~7_combout  = (\mem_data~1_combout  & ((exmem_ifout_o_2) # ((\mem_data~0_combout  & exmem_ifnext_pc_o_2)))) # (!\mem_data~1_combout  & (((\mem_data~0_combout  & exmem_ifnext_pc_o_2))))

	.dataa(\mem_data~1_combout ),
	.datab(exmem_ifout_o_2),
	.datac(\mem_data~0_combout ),
	.datad(\EXMEM|exmem_if.next_pc_o [2]),
	.cin(gnd),
	.combout(\mem_data~7_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~7 .lut_mask = 16'hF888;
defparam \mem_data~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N4
cycloneive_lcell_comb \mem_data~8 (
// Equation(s):
// \mem_data~8_combout  = (\mem_data~7_combout ) # ((\mem_data~3_combout  & ramiframload_2))

	.dataa(\mem_data~3_combout ),
	.datab(gnd),
	.datac(\mem_data~7_combout ),
	.datad(ramiframload_2),
	.cin(gnd),
	.combout(\mem_data~8_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~8 .lut_mask = 16'hFAF0;
defparam \mem_data~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N18
cycloneive_lcell_comb \rdat1[2]~5 (
// Equation(s):
// \rdat1[2]~5_combout  = (\rdat1[2]~4_combout ) # ((always03 & \mem_data~8_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(gnd),
	.datac(\rdat1[2]~4_combout ),
	.datad(\mem_data~8_combout ),
	.cin(gnd),
	.combout(\rdat1[2]~5_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[2]~5 .lut_mask = 16'hFAF0;
defparam \rdat1[2]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N8
cycloneive_lcell_comb \wdat~6 (
// Equation(s):
// \wdat~6_combout  = (!memwb_ifjal_o & ((memwb_ifmemToReg_o & (memwb_ifdmemload_o_4)) # (!memwb_ifmemToReg_o & ((memwb_ifout_o_4)))))

	.dataa(\MEMWB|memwb_if.dmemload_o [4]),
	.datab(\MEMWB|memwb_if.memToReg_o~q ),
	.datac(\MEMWB|memwb_if.out_o [4]),
	.datad(\MEMWB|memwb_if.jal_o~q ),
	.cin(gnd),
	.combout(\wdat~6_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~6 .lut_mask = 16'h00B8;
defparam \wdat~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N12
cycloneive_lcell_comb \wdat~7 (
// Equation(s):
// \wdat~7_combout  = (!memwb_iflui_o & ((\wdat~6_combout ) # ((memwb_ifnext_pc_o_4 & memwb_ifjal_o))))

	.dataa(\MEMWB|memwb_if.next_pc_o [4]),
	.datab(\MEMWB|memwb_if.jal_o~q ),
	.datac(\MEMWB|memwb_if.lui_o~q ),
	.datad(\wdat~6_combout ),
	.cin(gnd),
	.combout(\wdat~7_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~7 .lut_mask = 16'h0F08;
defparam \wdat~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N30
cycloneive_lcell_comb \rdat1[4]~6 (
// Equation(s):
// \rdat1[4]~6_combout  = (!always03 & ((always02 & ((\wdat~7_combout ))) # (!always02 & (idex_ifrdat1_o_4))))

	.dataa(\FU|always0~15_combout ),
	.datab(\FU|always0~11_combout ),
	.datac(\IDEX|idex_if.rdat1_o [4]),
	.datad(\wdat~7_combout ),
	.cin(gnd),
	.combout(\rdat1[4]~6_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[4]~6 .lut_mask = 16'h5410;
defparam \rdat1[4]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N2
cycloneive_lcell_comb \mem_data~9 (
// Equation(s):
// \mem_data~9_combout  = (\mem_data~1_combout  & ((exmem_ifout_o_4) # ((exmem_ifnext_pc_o_4 & \mem_data~0_combout )))) # (!\mem_data~1_combout  & (exmem_ifnext_pc_o_4 & (\mem_data~0_combout )))

	.dataa(\mem_data~1_combout ),
	.datab(\EXMEM|exmem_if.next_pc_o [4]),
	.datac(\mem_data~0_combout ),
	.datad(exmem_ifout_o_4),
	.cin(gnd),
	.combout(\mem_data~9_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~9 .lut_mask = 16'hEAC0;
defparam \mem_data~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N0
cycloneive_lcell_comb \mem_data~10 (
// Equation(s):
// \mem_data~10_combout  = (\mem_data~9_combout ) # ((\mem_data~3_combout  & ramiframload_4))

	.dataa(gnd),
	.datab(\mem_data~3_combout ),
	.datac(ramiframload_4),
	.datad(\mem_data~9_combout ),
	.cin(gnd),
	.combout(\mem_data~10_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~10 .lut_mask = 16'hFFC0;
defparam \mem_data~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N6
cycloneive_lcell_comb \rdat1[4]~7 (
// Equation(s):
// \rdat1[4]~7_combout  = (\rdat1[4]~6_combout ) # ((always03 & \mem_data~10_combout ))

	.dataa(gnd),
	.datab(\FU|always0~15_combout ),
	.datac(\rdat1[4]~6_combout ),
	.datad(\mem_data~10_combout ),
	.cin(gnd),
	.combout(\rdat1[4]~7_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[4]~7 .lut_mask = 16'hFCF0;
defparam \rdat1[4]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N16
cycloneive_lcell_comb \wdat~8 (
// Equation(s):
// \wdat~8_combout  = (!memwb_ifjal_o & ((memwb_ifmemToReg_o & (memwb_ifdmemload_o_3)) # (!memwb_ifmemToReg_o & ((memwb_ifout_o_3)))))

	.dataa(\MEMWB|memwb_if.dmemload_o [3]),
	.datab(\MEMWB|memwb_if.jal_o~q ),
	.datac(\MEMWB|memwb_if.out_o [3]),
	.datad(\MEMWB|memwb_if.memToReg_o~q ),
	.cin(gnd),
	.combout(\wdat~8_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~8 .lut_mask = 16'h2230;
defparam \wdat~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N2
cycloneive_lcell_comb \wdat~9 (
// Equation(s):
// \wdat~9_combout  = (!memwb_iflui_o & ((\wdat~8_combout ) # ((memwb_ifjal_o & memwb_ifnext_pc_o_3))))

	.dataa(\MEMWB|memwb_if.lui_o~q ),
	.datab(\MEMWB|memwb_if.jal_o~q ),
	.datac(\MEMWB|memwb_if.next_pc_o [3]),
	.datad(\wdat~8_combout ),
	.cin(gnd),
	.combout(\wdat~9_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~9 .lut_mask = 16'h5540;
defparam \wdat~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N2
cycloneive_lcell_comb \rdat1[3]~8 (
// Equation(s):
// \rdat1[3]~8_combout  = (!always03 & ((always02 & ((\wdat~9_combout ))) # (!always02 & (idex_ifrdat1_o_3))))

	.dataa(\FU|always0~11_combout ),
	.datab(\FU|always0~15_combout ),
	.datac(\IDEX|idex_if.rdat1_o [3]),
	.datad(\wdat~9_combout ),
	.cin(gnd),
	.combout(\rdat1[3]~8_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[3]~8 .lut_mask = 16'h3210;
defparam \rdat1[3]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N18
cycloneive_lcell_comb \mem_data~11 (
// Equation(s):
// \mem_data~11_combout  = (exmem_ifnext_pc_o_3 & ((\mem_data~0_combout ) # ((exmem_ifout_o_3 & \mem_data~1_combout )))) # (!exmem_ifnext_pc_o_3 & (exmem_ifout_o_3 & (\mem_data~1_combout )))

	.dataa(\EXMEM|exmem_if.next_pc_o [3]),
	.datab(exmem_ifout_o_3),
	.datac(\mem_data~1_combout ),
	.datad(\mem_data~0_combout ),
	.cin(gnd),
	.combout(\mem_data~11_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~11 .lut_mask = 16'hEAC0;
defparam \mem_data~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N6
cycloneive_lcell_comb \mem_data~12 (
// Equation(s):
// \mem_data~12_combout  = (\mem_data~11_combout ) # ((\mem_data~3_combout  & ramiframload_3))

	.dataa(\mem_data~3_combout ),
	.datab(\mem_data~11_combout ),
	.datac(gnd),
	.datad(ramiframload_3),
	.cin(gnd),
	.combout(\mem_data~12_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~12 .lut_mask = 16'hEECC;
defparam \mem_data~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N16
cycloneive_lcell_comb \rdat1[3]~9 (
// Equation(s):
// \rdat1[3]~9_combout  = (\rdat1[3]~8_combout ) # ((\mem_data~12_combout  & always03))

	.dataa(\mem_data~12_combout ),
	.datab(\rdat1[3]~8_combout ),
	.datac(gnd),
	.datad(\FU|always0~15_combout ),
	.cin(gnd),
	.combout(\rdat1[3]~9_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[3]~9 .lut_mask = 16'hEECC;
defparam \rdat1[3]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N14
cycloneive_lcell_comb \port_b~8 (
// Equation(s):
// \port_b~8_combout  = (idex_ifALUSel_o_1 & (((idex_ifimm_o_2)))) # (!idex_ifALUSel_o_1 & (idex_ifALUSel_o_0 & (idex_ifshamt_o_2)))

	.dataa(\IDEX|idex_if.ALUSel_o [0]),
	.datab(\IDEX|idex_if.shamt_o [2]),
	.datac(\IDEX|idex_if.ALUSel_o [1]),
	.datad(\IDEX|idex_if.imm_o [2]),
	.cin(gnd),
	.combout(\port_b~8_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~8 .lut_mask = 16'hF808;
defparam \port_b~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N28
cycloneive_lcell_comb \port_b~9 (
// Equation(s):
// \port_b~9_combout  = (\port_b~8_combout ) # ((idex_ifrdat2_o_2 & \port_b~2_combout ))

	.dataa(gnd),
	.datab(\IDEX|idex_if.rdat2_o [2]),
	.datac(\port_b~8_combout ),
	.datad(\port_b~2_combout ),
	.cin(gnd),
	.combout(\port_b~9_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~9 .lut_mask = 16'hFCF0;
defparam \port_b~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N0
cycloneive_lcell_comb \port_b~10 (
// Equation(s):
// \port_b~10_combout  = (\port_b~9_combout ) # ((\port_b~0_combout  & fuifrtReplace_2))

	.dataa(\port_b~9_combout ),
	.datab(\port_b~0_combout ),
	.datac(gnd),
	.datad(\FU|fuif.rtReplace[2]~6_combout ),
	.cin(gnd),
	.combout(\port_b~10_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~10 .lut_mask = 16'hEEAA;
defparam \port_b~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N2
cycloneive_lcell_comb \wdat~10 (
// Equation(s):
// \wdat~10_combout  = (!memwb_ifjal_o & ((memwb_ifmemToReg_o & (memwb_ifdmemload_o_8)) # (!memwb_ifmemToReg_o & ((memwb_ifout_o_8)))))

	.dataa(\MEMWB|memwb_if.dmemload_o [8]),
	.datab(\MEMWB|memwb_if.jal_o~q ),
	.datac(\MEMWB|memwb_if.out_o [8]),
	.datad(\MEMWB|memwb_if.memToReg_o~q ),
	.cin(gnd),
	.combout(\wdat~10_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~10 .lut_mask = 16'h2230;
defparam \wdat~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N6
cycloneive_lcell_comb \wdat~11 (
// Equation(s):
// \wdat~11_combout  = (!memwb_iflui_o & ((\wdat~10_combout ) # ((memwb_ifjal_o & memwb_ifnext_pc_o_8))))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.lui_o~q ),
	.datac(\MEMWB|memwb_if.next_pc_o [8]),
	.datad(\wdat~10_combout ),
	.cin(gnd),
	.combout(\wdat~11_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~11 .lut_mask = 16'h3320;
defparam \wdat~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N4
cycloneive_lcell_comb \rdat1[8]~10 (
// Equation(s):
// \rdat1[8]~10_combout  = (!always03 & ((always02 & ((\wdat~11_combout ))) # (!always02 & (idex_ifrdat1_o_8))))

	.dataa(\FU|always0~11_combout ),
	.datab(\IDEX|idex_if.rdat1_o [8]),
	.datac(\FU|always0~15_combout ),
	.datad(\wdat~11_combout ),
	.cin(gnd),
	.combout(\rdat1[8]~10_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[8]~10 .lut_mask = 16'h0E04;
defparam \rdat1[8]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N0
cycloneive_lcell_comb \mem_data~13 (
// Equation(s):
// \mem_data~13_combout  = (\mem_data~1_combout  & ((exmem_ifout_o_8) # ((exmem_ifnext_pc_o_8 & \mem_data~0_combout )))) # (!\mem_data~1_combout  & (((exmem_ifnext_pc_o_8 & \mem_data~0_combout ))))

	.dataa(\mem_data~1_combout ),
	.datab(exmem_ifout_o_8),
	.datac(\EXMEM|exmem_if.next_pc_o [8]),
	.datad(\mem_data~0_combout ),
	.cin(gnd),
	.combout(\mem_data~13_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~13 .lut_mask = 16'hF888;
defparam \mem_data~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N20
cycloneive_lcell_comb \mem_data~14 (
// Equation(s):
// \mem_data~14_combout  = (\mem_data~13_combout ) # ((\mem_data~3_combout  & ramiframload_8))

	.dataa(\mem_data~3_combout ),
	.datab(gnd),
	.datac(\mem_data~13_combout ),
	.datad(ramiframload_8),
	.cin(gnd),
	.combout(\mem_data~14_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~14 .lut_mask = 16'hFAF0;
defparam \mem_data~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N30
cycloneive_lcell_comb \rdat1[8]~11 (
// Equation(s):
// \rdat1[8]~11_combout  = (\rdat1[8]~10_combout ) # ((always03 & \mem_data~14_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(gnd),
	.datac(\rdat1[8]~10_combout ),
	.datad(\mem_data~14_combout ),
	.cin(gnd),
	.combout(\rdat1[8]~11_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[8]~11 .lut_mask = 16'hFAF0;
defparam \rdat1[8]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N14
cycloneive_lcell_comb \wdat~12 (
// Equation(s):
// \wdat~12_combout  = (!memwb_ifjal_o & ((memwb_ifmemToReg_o & (memwb_ifdmemload_o_7)) # (!memwb_ifmemToReg_o & ((memwb_ifout_o_7)))))

	.dataa(\MEMWB|memwb_if.memToReg_o~q ),
	.datab(\MEMWB|memwb_if.dmemload_o [7]),
	.datac(\MEMWB|memwb_if.out_o [7]),
	.datad(\MEMWB|memwb_if.jal_o~q ),
	.cin(gnd),
	.combout(\wdat~12_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~12 .lut_mask = 16'h00D8;
defparam \wdat~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N0
cycloneive_lcell_comb \wdat~13 (
// Equation(s):
// \wdat~13_combout  = (!memwb_iflui_o & ((\wdat~12_combout ) # ((memwb_ifnext_pc_o_7 & memwb_ifjal_o))))

	.dataa(\MEMWB|memwb_if.next_pc_o [7]),
	.datab(\MEMWB|memwb_if.jal_o~q ),
	.datac(\wdat~12_combout ),
	.datad(\MEMWB|memwb_if.lui_o~q ),
	.cin(gnd),
	.combout(\wdat~13_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~13 .lut_mask = 16'h00F8;
defparam \wdat~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N18
cycloneive_lcell_comb \rdat1[7]~12 (
// Equation(s):
// \rdat1[7]~12_combout  = (!always03 & ((always02 & ((\wdat~13_combout ))) # (!always02 & (idex_ifrdat1_o_7))))

	.dataa(\IDEX|idex_if.rdat1_o [7]),
	.datab(\FU|always0~15_combout ),
	.datac(\FU|always0~11_combout ),
	.datad(\wdat~13_combout ),
	.cin(gnd),
	.combout(\rdat1[7]~12_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[7]~12 .lut_mask = 16'h3202;
defparam \rdat1[7]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N14
cycloneive_lcell_comb \mem_data~15 (
// Equation(s):
// \mem_data~15_combout  = (exmem_ifout_o_7 & ((\mem_data~1_combout ) # ((exmem_ifnext_pc_o_7 & \mem_data~0_combout )))) # (!exmem_ifout_o_7 & (((exmem_ifnext_pc_o_7 & \mem_data~0_combout ))))

	.dataa(exmem_ifout_o_7),
	.datab(\mem_data~1_combout ),
	.datac(\EXMEM|exmem_if.next_pc_o [7]),
	.datad(\mem_data~0_combout ),
	.cin(gnd),
	.combout(\mem_data~15_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~15 .lut_mask = 16'hF888;
defparam \mem_data~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N8
cycloneive_lcell_comb \mem_data~16 (
// Equation(s):
// \mem_data~16_combout  = (\mem_data~15_combout ) # ((\mem_data~3_combout  & ramiframload_7))

	.dataa(\mem_data~3_combout ),
	.datab(gnd),
	.datac(ramiframload_7),
	.datad(\mem_data~15_combout ),
	.cin(gnd),
	.combout(\mem_data~16_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~16 .lut_mask = 16'hFFA0;
defparam \mem_data~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N6
cycloneive_lcell_comb \rdat1[7]~13 (
// Equation(s):
// \rdat1[7]~13_combout  = (\rdat1[7]~12_combout ) # ((always03 & \mem_data~16_combout ))

	.dataa(gnd),
	.datab(\FU|always0~15_combout ),
	.datac(\mem_data~16_combout ),
	.datad(\rdat1[7]~12_combout ),
	.cin(gnd),
	.combout(\rdat1[7]~13_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[7]~13 .lut_mask = 16'hFFC0;
defparam \rdat1[7]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N6
cycloneive_lcell_comb \wdat~14 (
// Equation(s):
// \wdat~14_combout  = (!memwb_ifjal_o & ((memwb_ifmemToReg_o & (memwb_ifdmemload_o_6)) # (!memwb_ifmemToReg_o & ((memwb_ifout_o_6)))))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.dmemload_o [6]),
	.datac(\MEMWB|memwb_if.out_o [6]),
	.datad(\MEMWB|memwb_if.memToReg_o~q ),
	.cin(gnd),
	.combout(\wdat~14_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~14 .lut_mask = 16'h4450;
defparam \wdat~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N4
cycloneive_lcell_comb \wdat~15 (
// Equation(s):
// \wdat~15_combout  = (!memwb_iflui_o & ((\wdat~14_combout ) # ((memwb_ifjal_o & memwb_ifnext_pc_o_6))))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.lui_o~q ),
	.datac(\MEMWB|memwb_if.next_pc_o [6]),
	.datad(\wdat~14_combout ),
	.cin(gnd),
	.combout(\wdat~15_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~15 .lut_mask = 16'h3320;
defparam \wdat~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N26
cycloneive_lcell_comb \rdat1[6]~14 (
// Equation(s):
// \rdat1[6]~14_combout  = (!always03 & ((always02 & ((\wdat~15_combout ))) # (!always02 & (idex_ifrdat1_o_6))))

	.dataa(\FU|always0~11_combout ),
	.datab(\IDEX|idex_if.rdat1_o [6]),
	.datac(\FU|always0~15_combout ),
	.datad(\wdat~15_combout ),
	.cin(gnd),
	.combout(\rdat1[6]~14_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[6]~14 .lut_mask = 16'h0E04;
defparam \rdat1[6]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N10
cycloneive_lcell_comb \mem_data~17 (
// Equation(s):
// \mem_data~17_combout  = (exmem_ifout_o_6 & ((\mem_data~1_combout ) # ((exmem_ifnext_pc_o_6 & \mem_data~0_combout )))) # (!exmem_ifout_o_6 & (exmem_ifnext_pc_o_6 & ((\mem_data~0_combout ))))

	.dataa(exmem_ifout_o_6),
	.datab(\EXMEM|exmem_if.next_pc_o [6]),
	.datac(\mem_data~1_combout ),
	.datad(\mem_data~0_combout ),
	.cin(gnd),
	.combout(\mem_data~17_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~17 .lut_mask = 16'hECA0;
defparam \mem_data~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N28
cycloneive_lcell_comb \mem_data~18 (
// Equation(s):
// \mem_data~18_combout  = (\mem_data~17_combout ) # ((\mem_data~3_combout  & ramiframload_6))

	.dataa(\mem_data~3_combout ),
	.datab(gnd),
	.datac(\mem_data~17_combout ),
	.datad(ramiframload_6),
	.cin(gnd),
	.combout(\mem_data~18_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~18 .lut_mask = 16'hFAF0;
defparam \mem_data~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N6
cycloneive_lcell_comb \rdat1[6]~15 (
// Equation(s):
// \rdat1[6]~15_combout  = (\rdat1[6]~14_combout ) # ((always03 & \mem_data~18_combout ))

	.dataa(gnd),
	.datab(\FU|always0~15_combout ),
	.datac(\rdat1[6]~14_combout ),
	.datad(\mem_data~18_combout ),
	.cin(gnd),
	.combout(\rdat1[6]~15_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[6]~15 .lut_mask = 16'hFCF0;
defparam \rdat1[6]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N24
cycloneive_lcell_comb \wdat~16 (
// Equation(s):
// \wdat~16_combout  = (!memwb_ifjal_o & ((memwb_ifmemToReg_o & (memwb_ifdmemload_o_5)) # (!memwb_ifmemToReg_o & ((memwb_ifout_o_5)))))

	.dataa(\MEMWB|memwb_if.dmemload_o [5]),
	.datab(\MEMWB|memwb_if.memToReg_o~q ),
	.datac(\MEMWB|memwb_if.out_o [5]),
	.datad(\MEMWB|memwb_if.jal_o~q ),
	.cin(gnd),
	.combout(\wdat~16_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~16 .lut_mask = 16'h00B8;
defparam \wdat~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N26
cycloneive_lcell_comb \wdat~17 (
// Equation(s):
// \wdat~17_combout  = (!memwb_iflui_o & ((\wdat~16_combout ) # ((memwb_ifnext_pc_o_5 & memwb_ifjal_o))))

	.dataa(\MEMWB|memwb_if.lui_o~q ),
	.datab(\wdat~16_combout ),
	.datac(\MEMWB|memwb_if.next_pc_o [5]),
	.datad(\MEMWB|memwb_if.jal_o~q ),
	.cin(gnd),
	.combout(\wdat~17_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~17 .lut_mask = 16'h5444;
defparam \wdat~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N12
cycloneive_lcell_comb \rdat1[5]~16 (
// Equation(s):
// \rdat1[5]~16_combout  = (!always03 & ((always02 & (\wdat~17_combout )) # (!always02 & ((idex_ifrdat1_o_5)))))

	.dataa(\FU|always0~11_combout ),
	.datab(\FU|always0~15_combout ),
	.datac(\wdat~17_combout ),
	.datad(\IDEX|idex_if.rdat1_o [5]),
	.cin(gnd),
	.combout(\rdat1[5]~16_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[5]~16 .lut_mask = 16'h3120;
defparam \rdat1[5]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N2
cycloneive_lcell_comb \mem_data~19 (
// Equation(s):
// \mem_data~19_combout  = (exmem_ifout_o_5 & ((\mem_data~1_combout ) # ((exmem_ifnext_pc_o_5 & \mem_data~0_combout )))) # (!exmem_ifout_o_5 & (exmem_ifnext_pc_o_5 & ((\mem_data~0_combout ))))

	.dataa(exmem_ifout_o_5),
	.datab(\EXMEM|exmem_if.next_pc_o [5]),
	.datac(\mem_data~1_combout ),
	.datad(\mem_data~0_combout ),
	.cin(gnd),
	.combout(\mem_data~19_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~19 .lut_mask = 16'hECA0;
defparam \mem_data~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N6
cycloneive_lcell_comb \mem_data~20 (
// Equation(s):
// \mem_data~20_combout  = (\mem_data~19_combout ) # ((\mem_data~3_combout  & ramiframload_5))

	.dataa(gnd),
	.datab(\mem_data~3_combout ),
	.datac(\mem_data~19_combout ),
	.datad(ramiframload_5),
	.cin(gnd),
	.combout(\mem_data~20_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~20 .lut_mask = 16'hFCF0;
defparam \mem_data~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N12
cycloneive_lcell_comb \rdat1[5]~17 (
// Equation(s):
// \rdat1[5]~17_combout  = (\rdat1[5]~16_combout ) # ((always03 & \mem_data~20_combout ))

	.dataa(gnd),
	.datab(\FU|always0~15_combout ),
	.datac(\rdat1[5]~16_combout ),
	.datad(\mem_data~20_combout ),
	.cin(gnd),
	.combout(\rdat1[5]~17_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[5]~17 .lut_mask = 16'hFCF0;
defparam \rdat1[5]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N12
cycloneive_lcell_comb \port_b~11 (
// Equation(s):
// \port_b~11_combout  = (!idex_ifALUSel_o_0 & !idex_ifALUSel_o_1)

	.dataa(gnd),
	.datab(gnd),
	.datac(\IDEX|idex_if.ALUSel_o [0]),
	.datad(\IDEX|idex_if.ALUSel_o [1]),
	.cin(gnd),
	.combout(\port_b~11_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~11 .lut_mask = 16'h000F;
defparam \port_b~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N26
cycloneive_lcell_comb \port_b~12 (
// Equation(s):
// \port_b~12_combout  = (\port_b~11_combout  & (idex_ifrdat2_o_3 & (!always01 & !always0)))

	.dataa(\port_b~11_combout ),
	.datab(\IDEX|idex_if.rdat2_o [3]),
	.datac(\FU|always0~7_combout ),
	.datad(\FU|always0~3_combout ),
	.cin(gnd),
	.combout(\port_b~12_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~12 .lut_mask = 16'h0008;
defparam \port_b~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N6
cycloneive_lcell_comb \port_b~13 (
// Equation(s):
// \port_b~13_combout  = (idex_ifALUSel_o_1 & (((idex_ifimm_o_3)))) # (!idex_ifALUSel_o_1 & (idex_ifALUSel_o_0 & (idex_ifshamt_o_3)))

	.dataa(\IDEX|idex_if.ALUSel_o [1]),
	.datab(\IDEX|idex_if.ALUSel_o [0]),
	.datac(\IDEX|idex_if.shamt_o [3]),
	.datad(\IDEX|idex_if.imm_o [3]),
	.cin(gnd),
	.combout(\port_b~13_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~13 .lut_mask = 16'hEA40;
defparam \port_b~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N2
cycloneive_lcell_comb \port_b~14 (
// Equation(s):
// \port_b~14_combout  = (\port_b~13_combout ) # ((\port_b~12_combout ) # ((\port_b~0_combout  & fuifrtReplace_3)))

	.dataa(\port_b~0_combout ),
	.datab(\port_b~13_combout ),
	.datac(\port_b~12_combout ),
	.datad(\FU|fuif.rtReplace[3]~7_combout ),
	.cin(gnd),
	.combout(\port_b~14_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~14 .lut_mask = 16'hFEFC;
defparam \port_b~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N24
cycloneive_lcell_comb \wdat~18 (
// Equation(s):
// \wdat~18_combout  = (memwb_iflui_o) # ((!memwb_ifjal_o & memwb_ifmemToReg_o))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.lui_o~q ),
	.datac(gnd),
	.datad(\MEMWB|memwb_if.memToReg_o~q ),
	.cin(gnd),
	.combout(\wdat~18_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~18 .lut_mask = 16'hDDCC;
defparam \wdat~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N6
cycloneive_lcell_comb \wdat~19 (
// Equation(s):
// \wdat~19_combout  = (memwb_ifjal_o) # (memwb_iflui_o)

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.lui_o~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wdat~19_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~19 .lut_mask = 16'hEEEE;
defparam \wdat~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N26
cycloneive_lcell_comb \wdat~20 (
// Equation(s):
// \wdat~20_combout  = (\wdat~19_combout  & ((memwb_ifnext_pc_o_16) # ((\wdat~18_combout )))) # (!\wdat~19_combout  & (((memwb_ifout_o_16 & !\wdat~18_combout ))))

	.dataa(\MEMWB|memwb_if.next_pc_o [16]),
	.datab(\wdat~19_combout ),
	.datac(\MEMWB|memwb_if.out_o [16]),
	.datad(\wdat~18_combout ),
	.cin(gnd),
	.combout(\wdat~20_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~20 .lut_mask = 16'hCCB8;
defparam \wdat~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N4
cycloneive_lcell_comb \wdat~21 (
// Equation(s):
// \wdat~21_combout  = (\wdat~18_combout  & ((\wdat~20_combout  & ((memwb_ifimm_o_0))) # (!\wdat~20_combout  & (memwb_ifdmemload_o_16)))) # (!\wdat~18_combout  & (((\wdat~20_combout ))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.dmemload_o [16]),
	.datac(\MEMWB|memwb_if.imm_o [0]),
	.datad(\wdat~20_combout ),
	.cin(gnd),
	.combout(\wdat~21_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~21 .lut_mask = 16'hF588;
defparam \wdat~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N8
cycloneive_lcell_comb \rdat1[16]~18 (
// Equation(s):
// \rdat1[16]~18_combout  = (!always03 & ((always02 & (\wdat~21_combout )) # (!always02 & ((idex_ifrdat1_o_16)))))

	.dataa(\FU|always0~15_combout ),
	.datab(\FU|always0~11_combout ),
	.datac(\wdat~21_combout ),
	.datad(\IDEX|idex_if.rdat1_o [16]),
	.cin(gnd),
	.combout(\rdat1[16]~18_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[16]~18 .lut_mask = 16'h5140;
defparam \rdat1[16]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N22
cycloneive_lcell_comb \mem_data~21 (
// Equation(s):
// \mem_data~21_combout  = (exmem_iflui_o) # ((!exmem_ifjal_o & exmem_ifmemToReg_o))

	.dataa(\EXMEM|exmem_if.lui_o~q ),
	.datab(\EXMEM|exmem_if.jal_o~q ),
	.datac(\EXMEM|exmem_if.memToReg_o~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_data~21_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~21 .lut_mask = 16'hBABA;
defparam \mem_data~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N10
cycloneive_lcell_comb \mem_data~22 (
// Equation(s):
// \mem_data~22_combout  = (!exmem_ifjal_o & !exmem_iflui_o)

	.dataa(gnd),
	.datab(\EXMEM|exmem_if.jal_o~q ),
	.datac(\EXMEM|exmem_if.lui_o~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_data~22_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~22 .lut_mask = 16'h0303;
defparam \mem_data~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N12
cycloneive_lcell_comb \mem_data~23 (
// Equation(s):
// \mem_data~23_combout  = (\mem_data~21_combout  & (((\mem_data~22_combout )))) # (!\mem_data~21_combout  & ((\mem_data~22_combout  & (exmem_ifout_o_16)) # (!\mem_data~22_combout  & ((exmem_ifnext_pc_o_16)))))

	.dataa(exmem_ifout_o_16),
	.datab(\mem_data~21_combout ),
	.datac(\EXMEM|exmem_if.next_pc_o [16]),
	.datad(\mem_data~22_combout ),
	.cin(gnd),
	.combout(\mem_data~23_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~23 .lut_mask = 16'hEE30;
defparam \mem_data~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N2
cycloneive_lcell_comb \mem_data~24 (
// Equation(s):
// \mem_data~24_combout  = (\mem_data~23_combout  & (((ramiframload_16)) # (!\mem_data~21_combout ))) # (!\mem_data~23_combout  & (\mem_data~21_combout  & (exmem_ifimm_o_0)))

	.dataa(\mem_data~23_combout ),
	.datab(\mem_data~21_combout ),
	.datac(\EXMEM|exmem_if.imm_o [0]),
	.datad(ramiframload_16),
	.cin(gnd),
	.combout(\mem_data~24_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~24 .lut_mask = 16'hEA62;
defparam \mem_data~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N20
cycloneive_lcell_comb \rdat1[16]~19 (
// Equation(s):
// \rdat1[16]~19_combout  = (\rdat1[16]~18_combout ) # ((always03 & \mem_data~24_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(gnd),
	.datac(\rdat1[16]~18_combout ),
	.datad(\mem_data~24_combout ),
	.cin(gnd),
	.combout(\rdat1[16]~19_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[16]~19 .lut_mask = 16'hFAF0;
defparam \rdat1[16]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N8
cycloneive_lcell_comb \wdat~22 (
// Equation(s):
// \wdat~22_combout  = (!memwb_ifjal_o & ((memwb_ifmemToReg_o & ((memwb_ifdmemload_o_15))) # (!memwb_ifmemToReg_o & (memwb_ifout_o_15))))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.memToReg_o~q ),
	.datac(\MEMWB|memwb_if.out_o [15]),
	.datad(\MEMWB|memwb_if.dmemload_o [15]),
	.cin(gnd),
	.combout(\wdat~22_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~22 .lut_mask = 16'h5410;
defparam \wdat~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N28
cycloneive_lcell_comb \wdat~23 (
// Equation(s):
// \wdat~23_combout  = (!memwb_iflui_o & ((\wdat~22_combout ) # ((memwb_ifjal_o & memwb_ifnext_pc_o_15))))

	.dataa(\wdat~22_combout ),
	.datab(\MEMWB|memwb_if.jal_o~q ),
	.datac(\MEMWB|memwb_if.next_pc_o [15]),
	.datad(\MEMWB|memwb_if.lui_o~q ),
	.cin(gnd),
	.combout(\wdat~23_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~23 .lut_mask = 16'h00EA;
defparam \wdat~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N26
cycloneive_lcell_comb \rdat1[15]~20 (
// Equation(s):
// \rdat1[15]~20_combout  = (!always03 & ((always02 & (\wdat~23_combout )) # (!always02 & ((idex_ifrdat1_o_15)))))

	.dataa(\wdat~23_combout ),
	.datab(\FU|always0~11_combout ),
	.datac(\FU|always0~15_combout ),
	.datad(\IDEX|idex_if.rdat1_o [15]),
	.cin(gnd),
	.combout(\rdat1[15]~20_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[15]~20 .lut_mask = 16'h0B08;
defparam \rdat1[15]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N28
cycloneive_lcell_comb \mem_data~25 (
// Equation(s):
// \mem_data~25_combout  = (\mem_data~1_combout  & ((exmem_ifout_o_15) # ((exmem_ifnext_pc_o_15 & \mem_data~0_combout )))) # (!\mem_data~1_combout  & (exmem_ifnext_pc_o_15 & ((\mem_data~0_combout ))))

	.dataa(\mem_data~1_combout ),
	.datab(\EXMEM|exmem_if.next_pc_o [15]),
	.datac(exmem_ifout_o_15),
	.datad(\mem_data~0_combout ),
	.cin(gnd),
	.combout(\mem_data~25_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~25 .lut_mask = 16'hECA0;
defparam \mem_data~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N0
cycloneive_lcell_comb \mem_data~26 (
// Equation(s):
// \mem_data~26_combout  = (\mem_data~25_combout ) # ((\mem_data~3_combout  & ramiframload_15))

	.dataa(gnd),
	.datab(\mem_data~3_combout ),
	.datac(ramiframload_15),
	.datad(\mem_data~25_combout ),
	.cin(gnd),
	.combout(\mem_data~26_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~26 .lut_mask = 16'hFFC0;
defparam \mem_data~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N14
cycloneive_lcell_comb \rdat1[15]~21 (
// Equation(s):
// \rdat1[15]~21_combout  = (\rdat1[15]~20_combout ) # ((always03 & \mem_data~26_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(gnd),
	.datac(\rdat1[15]~20_combout ),
	.datad(\mem_data~26_combout ),
	.cin(gnd),
	.combout(\rdat1[15]~21_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[15]~21 .lut_mask = 16'hFAF0;
defparam \rdat1[15]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N18
cycloneive_lcell_comb \wdat~24 (
// Equation(s):
// \wdat~24_combout  = (!memwb_ifjal_o & ((memwb_ifmemToReg_o & (memwb_ifdmemload_o_14)) # (!memwb_ifmemToReg_o & ((memwb_ifout_o_14)))))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.dmemload_o [14]),
	.datac(\MEMWB|memwb_if.out_o [14]),
	.datad(\MEMWB|memwb_if.memToReg_o~q ),
	.cin(gnd),
	.combout(\wdat~24_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~24 .lut_mask = 16'h4450;
defparam \wdat~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N0
cycloneive_lcell_comb \wdat~25 (
// Equation(s):
// \wdat~25_combout  = (!memwb_iflui_o & ((\wdat~24_combout ) # ((memwb_ifjal_o & memwb_ifnext_pc_o_14))))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.lui_o~q ),
	.datac(\MEMWB|memwb_if.next_pc_o [14]),
	.datad(\wdat~24_combout ),
	.cin(gnd),
	.combout(\wdat~25_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~25 .lut_mask = 16'h3320;
defparam \wdat~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N8
cycloneive_lcell_comb \rdat1[14]~22 (
// Equation(s):
// \rdat1[14]~22_combout  = (!always03 & ((always02 & ((\wdat~25_combout ))) # (!always02 & (idex_ifrdat1_o_14))))

	.dataa(\FU|always0~15_combout ),
	.datab(\IDEX|idex_if.rdat1_o [14]),
	.datac(\FU|always0~11_combout ),
	.datad(\wdat~25_combout ),
	.cin(gnd),
	.combout(\rdat1[14]~22_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[14]~22 .lut_mask = 16'h5404;
defparam \rdat1[14]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N12
cycloneive_lcell_comb \mem_data~27 (
// Equation(s):
// \mem_data~27_combout  = (\mem_data~1_combout  & ((exmem_ifout_o_14) # ((exmem_ifnext_pc_o_14 & \mem_data~0_combout )))) # (!\mem_data~1_combout  & (((exmem_ifnext_pc_o_14 & \mem_data~0_combout ))))

	.dataa(\mem_data~1_combout ),
	.datab(exmem_ifout_o_14),
	.datac(\EXMEM|exmem_if.next_pc_o [14]),
	.datad(\mem_data~0_combout ),
	.cin(gnd),
	.combout(\mem_data~27_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~27 .lut_mask = 16'hF888;
defparam \mem_data~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N20
cycloneive_lcell_comb \mem_data~28 (
// Equation(s):
// \mem_data~28_combout  = (\mem_data~27_combout ) # ((\mem_data~3_combout  & ramiframload_14))

	.dataa(gnd),
	.datab(\mem_data~3_combout ),
	.datac(ramiframload_14),
	.datad(\mem_data~27_combout ),
	.cin(gnd),
	.combout(\mem_data~28_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~28 .lut_mask = 16'hFFC0;
defparam \mem_data~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N14
cycloneive_lcell_comb \rdat1[14]~23 (
// Equation(s):
// \rdat1[14]~23_combout  = (\rdat1[14]~22_combout ) # ((always03 & \mem_data~28_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(gnd),
	.datac(\rdat1[14]~22_combout ),
	.datad(\mem_data~28_combout ),
	.cin(gnd),
	.combout(\rdat1[14]~23_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[14]~23 .lut_mask = 16'hFAF0;
defparam \rdat1[14]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N10
cycloneive_lcell_comb \wdat~26 (
// Equation(s):
// \wdat~26_combout  = (!memwb_ifjal_o & ((memwb_ifmemToReg_o & (memwb_ifdmemload_o_13)) # (!memwb_ifmemToReg_o & ((memwb_ifout_o_13)))))

	.dataa(\MEMWB|memwb_if.dmemload_o [13]),
	.datab(\MEMWB|memwb_if.jal_o~q ),
	.datac(\MEMWB|memwb_if.out_o [13]),
	.datad(\MEMWB|memwb_if.memToReg_o~q ),
	.cin(gnd),
	.combout(\wdat~26_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~26 .lut_mask = 16'h2230;
defparam \wdat~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N20
cycloneive_lcell_comb \wdat~27 (
// Equation(s):
// \wdat~27_combout  = (!memwb_iflui_o & ((\wdat~26_combout ) # ((memwb_ifnext_pc_o_13 & memwb_ifjal_o))))

	.dataa(\wdat~26_combout ),
	.datab(\MEMWB|memwb_if.lui_o~q ),
	.datac(\MEMWB|memwb_if.next_pc_o [13]),
	.datad(\MEMWB|memwb_if.jal_o~q ),
	.cin(gnd),
	.combout(\wdat~27_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~27 .lut_mask = 16'h3222;
defparam \wdat~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N4
cycloneive_lcell_comb \rdat1[13]~24 (
// Equation(s):
// \rdat1[13]~24_combout  = (!always03 & ((always02 & (\wdat~27_combout )) # (!always02 & ((idex_ifrdat1_o_13)))))

	.dataa(\FU|always0~15_combout ),
	.datab(\wdat~27_combout ),
	.datac(\IDEX|idex_if.rdat1_o [13]),
	.datad(\FU|always0~11_combout ),
	.cin(gnd),
	.combout(\rdat1[13]~24_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[13]~24 .lut_mask = 16'h4450;
defparam \rdat1[13]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N16
cycloneive_lcell_comb \mem_data~29 (
// Equation(s):
// \mem_data~29_combout  = (exmem_ifnext_pc_o_13 & ((\mem_data~0_combout ) # ((\mem_data~1_combout  & exmem_ifout_o_13)))) # (!exmem_ifnext_pc_o_13 & (((\mem_data~1_combout  & exmem_ifout_o_13))))

	.dataa(\EXMEM|exmem_if.next_pc_o [13]),
	.datab(\mem_data~0_combout ),
	.datac(\mem_data~1_combout ),
	.datad(exmem_ifout_o_13),
	.cin(gnd),
	.combout(\mem_data~29_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~29 .lut_mask = 16'hF888;
defparam \mem_data~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N30
cycloneive_lcell_comb \mem_data~30 (
// Equation(s):
// \mem_data~30_combout  = (\mem_data~29_combout ) # ((\mem_data~3_combout  & ramiframload_13))

	.dataa(gnd),
	.datab(\mem_data~3_combout ),
	.datac(ramiframload_13),
	.datad(\mem_data~29_combout ),
	.cin(gnd),
	.combout(\mem_data~30_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~30 .lut_mask = 16'hFFC0;
defparam \mem_data~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N12
cycloneive_lcell_comb \rdat1[13]~25 (
// Equation(s):
// \rdat1[13]~25_combout  = (\rdat1[13]~24_combout ) # ((always03 & \mem_data~30_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(gnd),
	.datac(\rdat1[13]~24_combout ),
	.datad(\mem_data~30_combout ),
	.cin(gnd),
	.combout(\rdat1[13]~25_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[13]~25 .lut_mask = 16'hFAF0;
defparam \rdat1[13]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N20
cycloneive_lcell_comb \wdat~28 (
// Equation(s):
// \wdat~28_combout  = (!memwb_ifjal_o & ((memwb_ifmemToReg_o & (memwb_ifdmemload_o_12)) # (!memwb_ifmemToReg_o & ((memwb_ifout_o_12)))))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.dmemload_o [12]),
	.datac(\MEMWB|memwb_if.out_o [12]),
	.datad(\MEMWB|memwb_if.memToReg_o~q ),
	.cin(gnd),
	.combout(\wdat~28_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~28 .lut_mask = 16'h4450;
defparam \wdat~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N8
cycloneive_lcell_comb \wdat~29 (
// Equation(s):
// \wdat~29_combout  = (!memwb_iflui_o & ((\wdat~28_combout ) # ((memwb_ifjal_o & memwb_ifnext_pc_o_12))))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.lui_o~q ),
	.datac(\MEMWB|memwb_if.next_pc_o [12]),
	.datad(\wdat~28_combout ),
	.cin(gnd),
	.combout(\wdat~29_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~29 .lut_mask = 16'h3320;
defparam \wdat~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N16
cycloneive_lcell_comb \rdat1[12]~26 (
// Equation(s):
// \rdat1[12]~26_combout  = (!always03 & ((always02 & ((\wdat~29_combout ))) # (!always02 & (idex_ifrdat1_o_12))))

	.dataa(\IDEX|idex_if.rdat1_o [12]),
	.datab(\wdat~29_combout ),
	.datac(\FU|always0~15_combout ),
	.datad(\FU|always0~11_combout ),
	.cin(gnd),
	.combout(\rdat1[12]~26_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[12]~26 .lut_mask = 16'h0C0A;
defparam \rdat1[12]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N10
cycloneive_lcell_comb \mem_data~31 (
// Equation(s):
// \mem_data~31_combout  = (\mem_data~0_combout  & ((exmem_ifnext_pc_o_12) # ((exmem_ifout_o_12 & \mem_data~1_combout )))) # (!\mem_data~0_combout  & (exmem_ifout_o_12 & ((\mem_data~1_combout ))))

	.dataa(\mem_data~0_combout ),
	.datab(exmem_ifout_o_12),
	.datac(\EXMEM|exmem_if.next_pc_o [12]),
	.datad(\mem_data~1_combout ),
	.cin(gnd),
	.combout(\mem_data~31_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~31 .lut_mask = 16'hECA0;
defparam \mem_data~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N18
cycloneive_lcell_comb \mem_data~32 (
// Equation(s):
// \mem_data~32_combout  = (\mem_data~31_combout ) # ((\mem_data~3_combout  & ramiframload_12))

	.dataa(\mem_data~3_combout ),
	.datab(gnd),
	.datac(\mem_data~31_combout ),
	.datad(ramiframload_12),
	.cin(gnd),
	.combout(\mem_data~32_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~32 .lut_mask = 16'hFAF0;
defparam \mem_data~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N28
cycloneive_lcell_comb \rdat1[12]~27 (
// Equation(s):
// \rdat1[12]~27_combout  = (\rdat1[12]~26_combout ) # ((always03 & \mem_data~32_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(gnd),
	.datac(\rdat1[12]~26_combout ),
	.datad(\mem_data~32_combout ),
	.cin(gnd),
	.combout(\rdat1[12]~27_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[12]~27 .lut_mask = 16'hFAF0;
defparam \rdat1[12]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N10
cycloneive_lcell_comb \wdat~30 (
// Equation(s):
// \wdat~30_combout  = (!memwb_ifjal_o & ((memwb_ifmemToReg_o & ((memwb_ifdmemload_o_11))) # (!memwb_ifmemToReg_o & (memwb_ifout_o_11))))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.memToReg_o~q ),
	.datac(\MEMWB|memwb_if.out_o [11]),
	.datad(\MEMWB|memwb_if.dmemload_o [11]),
	.cin(gnd),
	.combout(\wdat~30_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~30 .lut_mask = 16'h5410;
defparam \wdat~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N28
cycloneive_lcell_comb \wdat~31 (
// Equation(s):
// \wdat~31_combout  = (!memwb_iflui_o & ((\wdat~30_combout ) # ((memwb_ifjal_o & memwb_ifnext_pc_o_11))))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.lui_o~q ),
	.datac(\MEMWB|memwb_if.next_pc_o [11]),
	.datad(\wdat~30_combout ),
	.cin(gnd),
	.combout(\wdat~31_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~31 .lut_mask = 16'h3320;
defparam \wdat~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N14
cycloneive_lcell_comb \rdat1[11]~28 (
// Equation(s):
// \rdat1[11]~28_combout  = (!always03 & ((always02 & (\wdat~31_combout )) # (!always02 & ((idex_ifrdat1_o_11)))))

	.dataa(\FU|always0~11_combout ),
	.datab(\wdat~31_combout ),
	.datac(\IDEX|idex_if.rdat1_o [11]),
	.datad(\FU|always0~15_combout ),
	.cin(gnd),
	.combout(\rdat1[11]~28_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[11]~28 .lut_mask = 16'h00D8;
defparam \rdat1[11]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N0
cycloneive_lcell_comb \mem_data~33 (
// Equation(s):
// \mem_data~33_combout  = (exmem_ifout_o_11 & ((\mem_data~1_combout ) # ((exmem_ifnext_pc_o_11 & \mem_data~0_combout )))) # (!exmem_ifout_o_11 & (exmem_ifnext_pc_o_11 & (\mem_data~0_combout )))

	.dataa(exmem_ifout_o_11),
	.datab(\EXMEM|exmem_if.next_pc_o [11]),
	.datac(\mem_data~0_combout ),
	.datad(\mem_data~1_combout ),
	.cin(gnd),
	.combout(\mem_data~33_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~33 .lut_mask = 16'hEAC0;
defparam \mem_data~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N18
cycloneive_lcell_comb \mem_data~34 (
// Equation(s):
// \mem_data~34_combout  = (\mem_data~33_combout ) # ((\mem_data~3_combout  & ramiframload_111))

	.dataa(gnd),
	.datab(\mem_data~3_combout ),
	.datac(ramiframload_111),
	.datad(\mem_data~33_combout ),
	.cin(gnd),
	.combout(\mem_data~34_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~34 .lut_mask = 16'hFFC0;
defparam \mem_data~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N0
cycloneive_lcell_comb \rdat1[11]~29 (
// Equation(s):
// \rdat1[11]~29_combout  = (\rdat1[11]~28_combout ) # ((always03 & \mem_data~34_combout ))

	.dataa(\rdat1[11]~28_combout ),
	.datab(gnd),
	.datac(\FU|always0~15_combout ),
	.datad(\mem_data~34_combout ),
	.cin(gnd),
	.combout(\rdat1[11]~29_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[11]~29 .lut_mask = 16'hFAAA;
defparam \rdat1[11]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N12
cycloneive_lcell_comb \wdat~32 (
// Equation(s):
// \wdat~32_combout  = (!memwb_ifjal_o & ((memwb_ifmemToReg_o & (memwb_ifdmemload_o_10)) # (!memwb_ifmemToReg_o & ((memwb_ifout_o_10)))))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.dmemload_o [10]),
	.datac(\MEMWB|memwb_if.out_o [10]),
	.datad(\MEMWB|memwb_if.memToReg_o~q ),
	.cin(gnd),
	.combout(\wdat~32_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~32 .lut_mask = 16'h4450;
defparam \wdat~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N26
cycloneive_lcell_comb \wdat~33 (
// Equation(s):
// \wdat~33_combout  = (!memwb_iflui_o & ((\wdat~32_combout ) # ((memwb_ifjal_o & memwb_ifnext_pc_o_10))))

	.dataa(\MEMWB|memwb_if.jal_o~q ),
	.datab(\MEMWB|memwb_if.lui_o~q ),
	.datac(\MEMWB|memwb_if.next_pc_o [10]),
	.datad(\wdat~32_combout ),
	.cin(gnd),
	.combout(\wdat~33_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~33 .lut_mask = 16'h3320;
defparam \wdat~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N24
cycloneive_lcell_comb \rdat1[10]~30 (
// Equation(s):
// \rdat1[10]~30_combout  = (!always03 & ((always02 & ((\wdat~33_combout ))) # (!always02 & (idex_ifrdat1_o_10))))

	.dataa(\IDEX|idex_if.rdat1_o [10]),
	.datab(\FU|always0~15_combout ),
	.datac(\wdat~33_combout ),
	.datad(\FU|always0~11_combout ),
	.cin(gnd),
	.combout(\rdat1[10]~30_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[10]~30 .lut_mask = 16'h3022;
defparam \rdat1[10]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N30
cycloneive_lcell_comb \mem_data~35 (
// Equation(s):
// \mem_data~35_combout  = (exmem_ifout_o_10 & ((\mem_data~1_combout ) # ((exmem_ifnext_pc_o_10 & \mem_data~0_combout )))) # (!exmem_ifout_o_10 & (((exmem_ifnext_pc_o_10 & \mem_data~0_combout ))))

	.dataa(exmem_ifout_o_10),
	.datab(\mem_data~1_combout ),
	.datac(\EXMEM|exmem_if.next_pc_o [10]),
	.datad(\mem_data~0_combout ),
	.cin(gnd),
	.combout(\mem_data~35_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~35 .lut_mask = 16'hF888;
defparam \mem_data~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N6
cycloneive_lcell_comb \mem_data~36 (
// Equation(s):
// \mem_data~36_combout  = (\mem_data~35_combout ) # ((\mem_data~3_combout  & ramiframload_10))

	.dataa(gnd),
	.datab(\mem_data~35_combout ),
	.datac(\mem_data~3_combout ),
	.datad(ramiframload_10),
	.cin(gnd),
	.combout(\mem_data~36_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~36 .lut_mask = 16'hFCCC;
defparam \mem_data~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N0
cycloneive_lcell_comb \rdat1[10]~31 (
// Equation(s):
// \rdat1[10]~31_combout  = (\rdat1[10]~30_combout ) # ((always03 & \mem_data~36_combout ))

	.dataa(\rdat1[10]~30_combout ),
	.datab(gnd),
	.datac(\FU|always0~15_combout ),
	.datad(\mem_data~36_combout ),
	.cin(gnd),
	.combout(\rdat1[10]~31_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[10]~31 .lut_mask = 16'hFAAA;
defparam \rdat1[10]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N22
cycloneive_lcell_comb \wdat~34 (
// Equation(s):
// \wdat~34_combout  = (!memwb_ifjal_o & ((memwb_ifmemToReg_o & (memwb_ifdmemload_o_9)) # (!memwb_ifmemToReg_o & ((memwb_ifout_o_9)))))

	.dataa(\MEMWB|memwb_if.dmemload_o [9]),
	.datab(\MEMWB|memwb_if.jal_o~q ),
	.datac(\MEMWB|memwb_if.out_o [9]),
	.datad(\MEMWB|memwb_if.memToReg_o~q ),
	.cin(gnd),
	.combout(\wdat~34_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~34 .lut_mask = 16'h2230;
defparam \wdat~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N4
cycloneive_lcell_comb \wdat~35 (
// Equation(s):
// \wdat~35_combout  = (!memwb_iflui_o & ((\wdat~34_combout ) # ((memwb_ifnext_pc_o_9 & memwb_ifjal_o))))

	.dataa(\wdat~34_combout ),
	.datab(\MEMWB|memwb_if.lui_o~q ),
	.datac(\MEMWB|memwb_if.next_pc_o [9]),
	.datad(\MEMWB|memwb_if.jal_o~q ),
	.cin(gnd),
	.combout(\wdat~35_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~35 .lut_mask = 16'h3222;
defparam \wdat~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N22
cycloneive_lcell_comb \rdat1[9]~32 (
// Equation(s):
// \rdat1[9]~32_combout  = (!always03 & ((always02 & ((\wdat~35_combout ))) # (!always02 & (idex_ifrdat1_o_9))))

	.dataa(\IDEX|idex_if.rdat1_o [9]),
	.datab(\wdat~35_combout ),
	.datac(\FU|always0~11_combout ),
	.datad(\FU|always0~15_combout ),
	.cin(gnd),
	.combout(\rdat1[9]~32_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[9]~32 .lut_mask = 16'h00CA;
defparam \rdat1[9]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N24
cycloneive_lcell_comb \mem_data~37 (
// Equation(s):
// \mem_data~37_combout  = (exmem_ifout_o_9 & ((\mem_data~1_combout ) # ((exmem_ifnext_pc_o_9 & \mem_data~0_combout )))) # (!exmem_ifout_o_9 & (exmem_ifnext_pc_o_9 & ((\mem_data~0_combout ))))

	.dataa(exmem_ifout_o_9),
	.datab(\EXMEM|exmem_if.next_pc_o [9]),
	.datac(\mem_data~1_combout ),
	.datad(\mem_data~0_combout ),
	.cin(gnd),
	.combout(\mem_data~37_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~37 .lut_mask = 16'hECA0;
defparam \mem_data~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N24
cycloneive_lcell_comb \mem_data~38 (
// Equation(s):
// \mem_data~38_combout  = (\mem_data~37_combout ) # ((\mem_data~3_combout  & ramiframload_9))

	.dataa(gnd),
	.datab(\mem_data~3_combout ),
	.datac(ramiframload_9),
	.datad(\mem_data~37_combout ),
	.cin(gnd),
	.combout(\mem_data~38_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~38 .lut_mask = 16'hFFC0;
defparam \mem_data~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N18
cycloneive_lcell_comb \rdat1[9]~33 (
// Equation(s):
// \rdat1[9]~33_combout  = (\rdat1[9]~32_combout ) # ((always03 & \mem_data~38_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(gnd),
	.datac(\rdat1[9]~32_combout ),
	.datad(\mem_data~38_combout ),
	.cin(gnd),
	.combout(\rdat1[9]~33_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[9]~33 .lut_mask = 16'hFAF0;
defparam \rdat1[9]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N14
cycloneive_lcell_comb \port_b~15 (
// Equation(s):
// \port_b~15_combout  = (idex_ifrdat2_o_4 & (!always01 & (!always0 & \port_b~11_combout )))

	.dataa(\IDEX|idex_if.rdat2_o [4]),
	.datab(\FU|always0~7_combout ),
	.datac(\FU|always0~3_combout ),
	.datad(\port_b~11_combout ),
	.cin(gnd),
	.combout(\port_b~15_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~15 .lut_mask = 16'h0200;
defparam \port_b~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N10
cycloneive_lcell_comb \port_b~16 (
// Equation(s):
// \port_b~16_combout  = (idex_ifALUSel_o_1 & (((idex_ifimm_o_4)))) # (!idex_ifALUSel_o_1 & (idex_ifALUSel_o_0 & (idex_ifshamt_o_4)))

	.dataa(\IDEX|idex_if.ALUSel_o [1]),
	.datab(\IDEX|idex_if.ALUSel_o [0]),
	.datac(\IDEX|idex_if.shamt_o [4]),
	.datad(\IDEX|idex_if.imm_o [4]),
	.cin(gnd),
	.combout(\port_b~16_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~16 .lut_mask = 16'hEA40;
defparam \port_b~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N18
cycloneive_lcell_comb \port_b~17 (
// Equation(s):
// \port_b~17_combout  = (\port_b~16_combout ) # ((\port_b~15_combout ) # ((\port_b~0_combout  & fuifrtReplace_4)))

	.dataa(\port_b~16_combout ),
	.datab(\port_b~0_combout ),
	.datac(\port_b~15_combout ),
	.datad(\FU|fuif.rtReplace[4]~8_combout ),
	.cin(gnd),
	.combout(\port_b~17_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~17 .lut_mask = 16'hFEFA;
defparam \port_b~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N18
cycloneive_lcell_comb \wdat~36 (
// Equation(s):
// \wdat~36_combout  = (\wdat~18_combout  & ((memwb_ifdmemload_o_31) # ((\wdat~19_combout )))) # (!\wdat~18_combout  & (((memwb_ifout_o_31 & !\wdat~19_combout ))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.dmemload_o [31]),
	.datac(\MEMWB|memwb_if.out_o [31]),
	.datad(\wdat~19_combout ),
	.cin(gnd),
	.combout(\wdat~36_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~36 .lut_mask = 16'hAAD8;
defparam \wdat~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N2
cycloneive_lcell_comb \wdat~37 (
// Equation(s):
// \wdat~37_combout  = (\wdat~19_combout  & ((\wdat~36_combout  & (memwb_ifimm_o_15)) # (!\wdat~36_combout  & ((memwb_ifnext_pc_o_31))))) # (!\wdat~19_combout  & (((\wdat~36_combout ))))

	.dataa(\wdat~19_combout ),
	.datab(\MEMWB|memwb_if.imm_o [15]),
	.datac(\MEMWB|memwb_if.next_pc_o [31]),
	.datad(\wdat~36_combout ),
	.cin(gnd),
	.combout(\wdat~37_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~37 .lut_mask = 16'hDDA0;
defparam \wdat~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N28
cycloneive_lcell_comb \rdat1[31]~34 (
// Equation(s):
// \rdat1[31]~34_combout  = (!always03 & ((always02 & ((\wdat~37_combout ))) # (!always02 & (idex_ifrdat1_o_31))))

	.dataa(\FU|always0~15_combout ),
	.datab(\IDEX|idex_if.rdat1_o [31]),
	.datac(\FU|always0~11_combout ),
	.datad(\wdat~37_combout ),
	.cin(gnd),
	.combout(\rdat1[31]~34_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[31]~34 .lut_mask = 16'h5404;
defparam \rdat1[31]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N14
cycloneive_lcell_comb \mem_data~39 (
// Equation(s):
// \mem_data~39_combout  = (\mem_data~21_combout  & (((!\mem_data~22_combout )))) # (!\mem_data~21_combout  & ((\mem_data~22_combout  & (exmem_ifout_o_31)) # (!\mem_data~22_combout  & ((exmem_ifnext_pc_o_31)))))

	.dataa(\mem_data~21_combout ),
	.datab(exmem_ifout_o_31),
	.datac(\EXMEM|exmem_if.next_pc_o [31]),
	.datad(\mem_data~22_combout ),
	.cin(gnd),
	.combout(\mem_data~39_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~39 .lut_mask = 16'h44FA;
defparam \mem_data~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N22
cycloneive_lcell_comb \mem_data~40 (
// Equation(s):
// \mem_data~40_combout  = (\mem_data~39_combout  & (((exmem_ifimm_o_15)) # (!\mem_data~21_combout ))) # (!\mem_data~39_combout  & (\mem_data~21_combout  & (ramiframload_31)))

	.dataa(\mem_data~39_combout ),
	.datab(\mem_data~21_combout ),
	.datac(ramiframload_31),
	.datad(\EXMEM|exmem_if.imm_o [15]),
	.cin(gnd),
	.combout(\mem_data~40_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~40 .lut_mask = 16'hEA62;
defparam \mem_data~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N16
cycloneive_lcell_comb \rdat1[31]~35 (
// Equation(s):
// \rdat1[31]~35_combout  = (\rdat1[31]~34_combout ) # ((always03 & \mem_data~40_combout ))

	.dataa(gnd),
	.datab(\FU|always0~15_combout ),
	.datac(\mem_data~40_combout ),
	.datad(\rdat1[31]~34_combout ),
	.cin(gnd),
	.combout(\rdat1[31]~35_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[31]~35 .lut_mask = 16'hFFC0;
defparam \rdat1[31]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N16
cycloneive_lcell_comb \wdat~38 (
// Equation(s):
// \wdat~38_combout  = (\wdat~18_combout  & ((memwb_ifdmemload_o_29) # ((\wdat~19_combout )))) # (!\wdat~18_combout  & (((memwb_ifout_o_29 & !\wdat~19_combout ))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.dmemload_o [29]),
	.datac(\MEMWB|memwb_if.out_o [29]),
	.datad(\wdat~19_combout ),
	.cin(gnd),
	.combout(\wdat~38_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~38 .lut_mask = 16'hAAD8;
defparam \wdat~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N12
cycloneive_lcell_comb \wdat~39 (
// Equation(s):
// \wdat~39_combout  = (\wdat~19_combout  & ((\wdat~38_combout  & (memwb_ifimm_o_13)) # (!\wdat~38_combout  & ((memwb_ifnext_pc_o_29))))) # (!\wdat~19_combout  & (((\wdat~38_combout ))))

	.dataa(\MEMWB|memwb_if.imm_o [13]),
	.datab(\wdat~19_combout ),
	.datac(\MEMWB|memwb_if.next_pc_o [29]),
	.datad(\wdat~38_combout ),
	.cin(gnd),
	.combout(\wdat~39_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~39 .lut_mask = 16'hBBC0;
defparam \wdat~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N26
cycloneive_lcell_comb \rdat1[29]~36 (
// Equation(s):
// \rdat1[29]~36_combout  = (!always03 & ((always02 & ((\wdat~39_combout ))) # (!always02 & (idex_ifrdat1_o_29))))

	.dataa(\FU|always0~15_combout ),
	.datab(\IDEX|idex_if.rdat1_o [29]),
	.datac(\wdat~39_combout ),
	.datad(\FU|always0~11_combout ),
	.cin(gnd),
	.combout(\rdat1[29]~36_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[29]~36 .lut_mask = 16'h5044;
defparam \rdat1[29]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N10
cycloneive_lcell_comb \mem_data~41 (
// Equation(s):
// \mem_data~41_combout  = (\mem_data~21_combout  & (((!\mem_data~22_combout )))) # (!\mem_data~21_combout  & ((\mem_data~22_combout  & ((exmem_ifout_o_29))) # (!\mem_data~22_combout  & (exmem_ifnext_pc_o_29))))

	.dataa(\EXMEM|exmem_if.next_pc_o [29]),
	.datab(exmem_ifout_o_29),
	.datac(\mem_data~21_combout ),
	.datad(\mem_data~22_combout ),
	.cin(gnd),
	.combout(\mem_data~41_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~41 .lut_mask = 16'h0CFA;
defparam \mem_data~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N0
cycloneive_lcell_comb \mem_data~42 (
// Equation(s):
// \mem_data~42_combout  = (\mem_data~21_combout  & ((\mem_data~41_combout  & (exmem_ifimm_o_13)) # (!\mem_data~41_combout  & ((ramiframload_29))))) # (!\mem_data~21_combout  & (((\mem_data~41_combout ))))

	.dataa(\mem_data~21_combout ),
	.datab(\EXMEM|exmem_if.imm_o [13]),
	.datac(ramiframload_29),
	.datad(\mem_data~41_combout ),
	.cin(gnd),
	.combout(\mem_data~42_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~42 .lut_mask = 16'hDDA0;
defparam \mem_data~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N2
cycloneive_lcell_comb \rdat1[29]~37 (
// Equation(s):
// \rdat1[29]~37_combout  = (\rdat1[29]~36_combout ) # ((always03 & \mem_data~42_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(gnd),
	.datac(\rdat1[29]~36_combout ),
	.datad(\mem_data~42_combout ),
	.cin(gnd),
	.combout(\rdat1[29]~37_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[29]~37 .lut_mask = 16'hFAF0;
defparam \rdat1[29]~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N28
cycloneive_lcell_comb \wdat~40 (
// Equation(s):
// \wdat~40_combout  = (\wdat~18_combout  & (((\wdat~19_combout )))) # (!\wdat~18_combout  & ((\wdat~19_combout  & (memwb_ifnext_pc_o_30)) # (!\wdat~19_combout  & ((memwb_ifout_o_30)))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.next_pc_o [30]),
	.datac(\MEMWB|memwb_if.out_o [30]),
	.datad(\wdat~19_combout ),
	.cin(gnd),
	.combout(\wdat~40_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~40 .lut_mask = 16'hEE50;
defparam \wdat~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N30
cycloneive_lcell_comb \wdat~41 (
// Equation(s):
// \wdat~41_combout  = (\wdat~18_combout  & ((\wdat~40_combout  & (memwb_ifimm_o_14)) # (!\wdat~40_combout  & ((memwb_ifdmemload_o_30))))) # (!\wdat~18_combout  & (((\wdat~40_combout ))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.imm_o [14]),
	.datac(\MEMWB|memwb_if.dmemload_o [30]),
	.datad(\wdat~40_combout ),
	.cin(gnd),
	.combout(\wdat~41_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~41 .lut_mask = 16'hDDA0;
defparam \wdat~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N26
cycloneive_lcell_comb \rdat1[30]~38 (
// Equation(s):
// \rdat1[30]~38_combout  = (!always03 & ((always02 & (\wdat~41_combout )) # (!always02 & ((idex_ifrdat1_o_30)))))

	.dataa(\FU|always0~11_combout ),
	.datab(\wdat~41_combout ),
	.datac(\IDEX|idex_if.rdat1_o [30]),
	.datad(\FU|always0~15_combout ),
	.cin(gnd),
	.combout(\rdat1[30]~38_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[30]~38 .lut_mask = 16'h00D8;
defparam \rdat1[30]~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N0
cycloneive_lcell_comb \mem_data~43 (
// Equation(s):
// \mem_data~43_combout  = (\mem_data~22_combout  & ((exmem_ifout_o_30) # ((\mem_data~21_combout )))) # (!\mem_data~22_combout  & (((!\mem_data~21_combout  & exmem_ifnext_pc_o_30))))

	.dataa(\mem_data~22_combout ),
	.datab(exmem_ifout_o_30),
	.datac(\mem_data~21_combout ),
	.datad(\EXMEM|exmem_if.next_pc_o [30]),
	.cin(gnd),
	.combout(\mem_data~43_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~43 .lut_mask = 16'hADA8;
defparam \mem_data~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N10
cycloneive_lcell_comb \mem_data~44 (
// Equation(s):
// \mem_data~44_combout  = (\mem_data~43_combout  & (((ramiframload_30)) # (!\mem_data~21_combout ))) # (!\mem_data~43_combout  & (\mem_data~21_combout  & (exmem_ifimm_o_14)))

	.dataa(\mem_data~43_combout ),
	.datab(\mem_data~21_combout ),
	.datac(\EXMEM|exmem_if.imm_o [14]),
	.datad(ramiframload_30),
	.cin(gnd),
	.combout(\mem_data~44_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~44 .lut_mask = 16'hEA62;
defparam \mem_data~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N0
cycloneive_lcell_comb \rdat1[30]~39 (
// Equation(s):
// \rdat1[30]~39_combout  = (\rdat1[30]~38_combout ) # ((always03 & \mem_data~44_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(gnd),
	.datac(\rdat1[30]~38_combout ),
	.datad(\mem_data~44_combout ),
	.cin(gnd),
	.combout(\rdat1[30]~39_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[30]~39 .lut_mask = 16'hFAF0;
defparam \rdat1[30]~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N0
cycloneive_lcell_comb \wdat~42 (
// Equation(s):
// \wdat~42_combout  = (\wdat~18_combout  & (((\wdat~19_combout )))) # (!\wdat~18_combout  & ((\wdat~19_combout  & (memwb_ifnext_pc_o_28)) # (!\wdat~19_combout  & ((memwb_ifout_o_28)))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.next_pc_o [28]),
	.datac(\MEMWB|memwb_if.out_o [28]),
	.datad(\wdat~19_combout ),
	.cin(gnd),
	.combout(\wdat~42_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~42 .lut_mask = 16'hEE50;
defparam \wdat~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N22
cycloneive_lcell_comb \wdat~43 (
// Equation(s):
// \wdat~43_combout  = (\wdat~18_combout  & ((\wdat~42_combout  & (memwb_ifimm_o_12)) # (!\wdat~42_combout  & ((memwb_ifdmemload_o_28))))) # (!\wdat~18_combout  & (((\wdat~42_combout ))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.imm_o [12]),
	.datac(\MEMWB|memwb_if.dmemload_o [28]),
	.datad(\wdat~42_combout ),
	.cin(gnd),
	.combout(\wdat~43_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~43 .lut_mask = 16'hDDA0;
defparam \wdat~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N30
cycloneive_lcell_comb \rdat1[28]~40 (
// Equation(s):
// \rdat1[28]~40_combout  = (!always03 & ((always02 & ((\wdat~43_combout ))) # (!always02 & (idex_ifrdat1_o_28))))

	.dataa(\FU|always0~15_combout ),
	.datab(\IDEX|idex_if.rdat1_o [28]),
	.datac(\FU|always0~11_combout ),
	.datad(\wdat~43_combout ),
	.cin(gnd),
	.combout(\rdat1[28]~40_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[28]~40 .lut_mask = 16'h5404;
defparam \rdat1[28]~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N14
cycloneive_lcell_comb \mem_data~45 (
// Equation(s):
// \mem_data~45_combout  = (\mem_data~21_combout  & (((\mem_data~22_combout )))) # (!\mem_data~21_combout  & ((\mem_data~22_combout  & ((exmem_ifout_o_28))) # (!\mem_data~22_combout  & (exmem_ifnext_pc_o_28))))

	.dataa(\EXMEM|exmem_if.next_pc_o [28]),
	.datab(\mem_data~21_combout ),
	.datac(exmem_ifout_o_28),
	.datad(\mem_data~22_combout ),
	.cin(gnd),
	.combout(\mem_data~45_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~45 .lut_mask = 16'hFC22;
defparam \mem_data~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N20
cycloneive_lcell_comb \mem_data~46 (
// Equation(s):
// \mem_data~46_combout  = (\mem_data~45_combout  & (((ramiframload_28)) # (!\mem_data~21_combout ))) # (!\mem_data~45_combout  & (\mem_data~21_combout  & ((exmem_ifimm_o_12))))

	.dataa(\mem_data~45_combout ),
	.datab(\mem_data~21_combout ),
	.datac(ramiframload_28),
	.datad(\EXMEM|exmem_if.imm_o [12]),
	.cin(gnd),
	.combout(\mem_data~46_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~46 .lut_mask = 16'hE6A2;
defparam \mem_data~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N26
cycloneive_lcell_comb \rdat1[28]~41 (
// Equation(s):
// \rdat1[28]~41_combout  = (\rdat1[28]~40_combout ) # ((always03 & \mem_data~46_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(gnd),
	.datac(\rdat1[28]~40_combout ),
	.datad(\mem_data~46_combout ),
	.cin(gnd),
	.combout(\rdat1[28]~41_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[28]~41 .lut_mask = 16'hFAF0;
defparam \rdat1[28]~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N24
cycloneive_lcell_comb \wdat~44 (
// Equation(s):
// \wdat~44_combout  = (\wdat~18_combout  & (((\wdat~19_combout )))) # (!\wdat~18_combout  & ((\wdat~19_combout  & (memwb_ifnext_pc_o_26)) # (!\wdat~19_combout  & ((memwb_ifout_o_26)))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.next_pc_o [26]),
	.datac(\MEMWB|memwb_if.out_o [26]),
	.datad(\wdat~19_combout ),
	.cin(gnd),
	.combout(\wdat~44_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~44 .lut_mask = 16'hEE50;
defparam \wdat~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N20
cycloneive_lcell_comb \wdat~45 (
// Equation(s):
// \wdat~45_combout  = (\wdat~18_combout  & ((\wdat~44_combout  & (memwb_ifimm_o_10)) # (!\wdat~44_combout  & ((memwb_ifdmemload_o_26))))) # (!\wdat~18_combout  & (((\wdat~44_combout ))))

	.dataa(\MEMWB|memwb_if.imm_o [10]),
	.datab(\wdat~18_combout ),
	.datac(\MEMWB|memwb_if.dmemload_o [26]),
	.datad(\wdat~44_combout ),
	.cin(gnd),
	.combout(\wdat~45_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~45 .lut_mask = 16'hBBC0;
defparam \wdat~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N26
cycloneive_lcell_comb \rdat1[26]~42 (
// Equation(s):
// \rdat1[26]~42_combout  = (!always03 & ((always02 & ((\wdat~45_combout ))) # (!always02 & (idex_ifrdat1_o_26))))

	.dataa(\FU|always0~15_combout ),
	.datab(\IDEX|idex_if.rdat1_o [26]),
	.datac(\FU|always0~11_combout ),
	.datad(\wdat~45_combout ),
	.cin(gnd),
	.combout(\rdat1[26]~42_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[26]~42 .lut_mask = 16'h5404;
defparam \rdat1[26]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N4
cycloneive_lcell_comb \mem_data~47 (
// Equation(s):
// \mem_data~47_combout  = (\mem_data~21_combout  & (((\mem_data~22_combout )))) # (!\mem_data~21_combout  & ((\mem_data~22_combout  & ((exmem_ifout_o_26))) # (!\mem_data~22_combout  & (exmem_ifnext_pc_o_26))))

	.dataa(\mem_data~21_combout ),
	.datab(\EXMEM|exmem_if.next_pc_o [26]),
	.datac(\mem_data~22_combout ),
	.datad(exmem_ifout_o_26),
	.cin(gnd),
	.combout(\mem_data~47_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~47 .lut_mask = 16'hF4A4;
defparam \mem_data~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N14
cycloneive_lcell_comb \mem_data~48 (
// Equation(s):
// \mem_data~48_combout  = (\mem_data~21_combout  & ((\mem_data~47_combout  & ((ramiframload_26))) # (!\mem_data~47_combout  & (exmem_ifimm_o_10)))) # (!\mem_data~21_combout  & (((\mem_data~47_combout ))))

	.dataa(\mem_data~21_combout ),
	.datab(\EXMEM|exmem_if.imm_o [10]),
	.datac(\mem_data~47_combout ),
	.datad(ramiframload_26),
	.cin(gnd),
	.combout(\mem_data~48_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~48 .lut_mask = 16'hF858;
defparam \mem_data~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N8
cycloneive_lcell_comb \rdat1[26]~43 (
// Equation(s):
// \rdat1[26]~43_combout  = (\rdat1[26]~42_combout ) # ((always03 & \mem_data~48_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(\mem_data~48_combout ),
	.datac(gnd),
	.datad(\rdat1[26]~42_combout ),
	.cin(gnd),
	.combout(\rdat1[26]~43_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[26]~43 .lut_mask = 16'hFF88;
defparam \rdat1[26]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N20
cycloneive_lcell_comb \wdat~46 (
// Equation(s):
// \wdat~46_combout  = (\wdat~18_combout  & ((memwb_ifdmemload_o_27) # ((\wdat~19_combout )))) # (!\wdat~18_combout  & (((memwb_ifout_o_27 & !\wdat~19_combout ))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.dmemload_o [27]),
	.datac(\MEMWB|memwb_if.out_o [27]),
	.datad(\wdat~19_combout ),
	.cin(gnd),
	.combout(\wdat~46_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~46 .lut_mask = 16'hAAD8;
defparam \wdat~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N16
cycloneive_lcell_comb \wdat~47 (
// Equation(s):
// \wdat~47_combout  = (\wdat~46_combout  & ((memwb_ifimm_o_11) # ((!\wdat~19_combout )))) # (!\wdat~46_combout  & (((memwb_ifnext_pc_o_27 & \wdat~19_combout ))))

	.dataa(\MEMWB|memwb_if.imm_o [11]),
	.datab(\wdat~46_combout ),
	.datac(\MEMWB|memwb_if.next_pc_o [27]),
	.datad(\wdat~19_combout ),
	.cin(gnd),
	.combout(\wdat~47_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~47 .lut_mask = 16'hB8CC;
defparam \wdat~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N28
cycloneive_lcell_comb \rdat1[27]~44 (
// Equation(s):
// \rdat1[27]~44_combout  = (!always03 & ((always02 & (\wdat~47_combout )) # (!always02 & ((idex_ifrdat1_o_27)))))

	.dataa(\FU|always0~11_combout ),
	.datab(\wdat~47_combout ),
	.datac(\FU|always0~15_combout ),
	.datad(\IDEX|idex_if.rdat1_o [27]),
	.cin(gnd),
	.combout(\rdat1[27]~44_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[27]~44 .lut_mask = 16'h0D08;
defparam \rdat1[27]~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N10
cycloneive_lcell_comb \mem_data~49 (
// Equation(s):
// \mem_data~49_combout  = (\mem_data~22_combout  & (((exmem_ifout_o_27 & !\mem_data~21_combout )))) # (!\mem_data~22_combout  & ((exmem_ifnext_pc_o_27) # ((\mem_data~21_combout ))))

	.dataa(\EXMEM|exmem_if.next_pc_o [27]),
	.datab(exmem_ifout_o_27),
	.datac(\mem_data~22_combout ),
	.datad(\mem_data~21_combout ),
	.cin(gnd),
	.combout(\mem_data~49_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~49 .lut_mask = 16'h0FCA;
defparam \mem_data~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N6
cycloneive_lcell_comb \mem_data~50 (
// Equation(s):
// \mem_data~50_combout  = (\mem_data~21_combout  & ((\mem_data~49_combout  & (exmem_ifimm_o_11)) # (!\mem_data~49_combout  & ((ramiframload_27))))) # (!\mem_data~21_combout  & (\mem_data~49_combout ))

	.dataa(\mem_data~21_combout ),
	.datab(\mem_data~49_combout ),
	.datac(\EXMEM|exmem_if.imm_o [11]),
	.datad(ramiframload_27),
	.cin(gnd),
	.combout(\mem_data~50_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~50 .lut_mask = 16'hE6C4;
defparam \mem_data~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N4
cycloneive_lcell_comb \rdat1[27]~45 (
// Equation(s):
// \rdat1[27]~45_combout  = (\rdat1[27]~44_combout ) # ((always03 & \mem_data~50_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(\rdat1[27]~44_combout ),
	.datac(gnd),
	.datad(\mem_data~50_combout ),
	.cin(gnd),
	.combout(\rdat1[27]~45_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[27]~45 .lut_mask = 16'hEECC;
defparam \rdat1[27]~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N0
cycloneive_lcell_comb \wdat~48 (
// Equation(s):
// \wdat~48_combout  = (\wdat~18_combout  & ((\wdat~19_combout ) # ((memwb_ifdmemload_o_25)))) # (!\wdat~18_combout  & (!\wdat~19_combout  & (memwb_ifout_o_25)))

	.dataa(\wdat~18_combout ),
	.datab(\wdat~19_combout ),
	.datac(\MEMWB|memwb_if.out_o [25]),
	.datad(\MEMWB|memwb_if.dmemload_o [25]),
	.cin(gnd),
	.combout(\wdat~48_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~48 .lut_mask = 16'hBA98;
defparam \wdat~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N24
cycloneive_lcell_comb \wdat~49 (
// Equation(s):
// \wdat~49_combout  = (\wdat~48_combout  & ((memwb_ifimm_o_9) # ((!\wdat~19_combout )))) # (!\wdat~48_combout  & (((memwb_ifnext_pc_o_25 & \wdat~19_combout ))))

	.dataa(\MEMWB|memwb_if.imm_o [9]),
	.datab(\wdat~48_combout ),
	.datac(\MEMWB|memwb_if.next_pc_o [25]),
	.datad(\wdat~19_combout ),
	.cin(gnd),
	.combout(\wdat~49_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~49 .lut_mask = 16'hB8CC;
defparam \wdat~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N24
cycloneive_lcell_comb \rdat1[25]~46 (
// Equation(s):
// \rdat1[25]~46_combout  = (!always03 & ((always02 & ((\wdat~49_combout ))) # (!always02 & (idex_ifrdat1_o_25))))

	.dataa(\FU|always0~11_combout ),
	.datab(\IDEX|idex_if.rdat1_o [25]),
	.datac(\wdat~49_combout ),
	.datad(\FU|always0~15_combout ),
	.cin(gnd),
	.combout(\rdat1[25]~46_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[25]~46 .lut_mask = 16'h00E4;
defparam \rdat1[25]~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N6
cycloneive_lcell_comb \mem_data~51 (
// Equation(s):
// \mem_data~51_combout  = (\mem_data~21_combout  & (((!\mem_data~22_combout )))) # (!\mem_data~21_combout  & ((\mem_data~22_combout  & (exmem_ifout_o_25)) # (!\mem_data~22_combout  & ((exmem_ifnext_pc_o_25)))))

	.dataa(\mem_data~21_combout ),
	.datab(exmem_ifout_o_25),
	.datac(\mem_data~22_combout ),
	.datad(\EXMEM|exmem_if.next_pc_o [25]),
	.cin(gnd),
	.combout(\mem_data~51_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~51 .lut_mask = 16'h4F4A;
defparam \mem_data~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N6
cycloneive_lcell_comb \mem_data~52 (
// Equation(s):
// \mem_data~52_combout  = (\mem_data~51_combout  & (((exmem_ifimm_o_9)) # (!\mem_data~21_combout ))) # (!\mem_data~51_combout  & (\mem_data~21_combout  & ((ramiframload_25))))

	.dataa(\mem_data~51_combout ),
	.datab(\mem_data~21_combout ),
	.datac(\EXMEM|exmem_if.imm_o [9]),
	.datad(ramiframload_25),
	.cin(gnd),
	.combout(\mem_data~52_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~52 .lut_mask = 16'hE6A2;
defparam \mem_data~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N28
cycloneive_lcell_comb \rdat1[25]~47 (
// Equation(s):
// \rdat1[25]~47_combout  = (\rdat1[25]~46_combout ) # ((always03 & \mem_data~52_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(\rdat1[25]~46_combout ),
	.datac(gnd),
	.datad(\mem_data~52_combout ),
	.cin(gnd),
	.combout(\rdat1[25]~47_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[25]~47 .lut_mask = 16'hEECC;
defparam \rdat1[25]~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N20
cycloneive_lcell_comb \wdat~50 (
// Equation(s):
// \wdat~50_combout  = (\wdat~18_combout  & (((\wdat~19_combout )))) # (!\wdat~18_combout  & ((\wdat~19_combout  & (memwb_ifnext_pc_o_24)) # (!\wdat~19_combout  & ((memwb_ifout_o_24)))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.next_pc_o [24]),
	.datac(\MEMWB|memwb_if.out_o [24]),
	.datad(\wdat~19_combout ),
	.cin(gnd),
	.combout(\wdat~50_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~50 .lut_mask = 16'hEE50;
defparam \wdat~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N28
cycloneive_lcell_comb \wdat~51 (
// Equation(s):
// \wdat~51_combout  = (\wdat~18_combout  & ((\wdat~50_combout  & (memwb_ifimm_o_8)) # (!\wdat~50_combout  & ((memwb_ifdmemload_o_24))))) # (!\wdat~18_combout  & (((\wdat~50_combout ))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.imm_o [8]),
	.datac(\MEMWB|memwb_if.dmemload_o [24]),
	.datad(\wdat~50_combout ),
	.cin(gnd),
	.combout(\wdat~51_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~51 .lut_mask = 16'hDDA0;
defparam \wdat~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N4
cycloneive_lcell_comb \rdat1[24]~48 (
// Equation(s):
// \rdat1[24]~48_combout  = (!always03 & ((always02 & (\wdat~51_combout )) # (!always02 & ((idex_ifrdat1_o_24)))))

	.dataa(\FU|always0~15_combout ),
	.datab(\wdat~51_combout ),
	.datac(\FU|always0~11_combout ),
	.datad(\IDEX|idex_if.rdat1_o [24]),
	.cin(gnd),
	.combout(\rdat1[24]~48_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[24]~48 .lut_mask = 16'h4540;
defparam \rdat1[24]~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N6
cycloneive_lcell_comb \mem_data~53 (
// Equation(s):
// \mem_data~53_combout  = (\mem_data~22_combout  & ((\mem_data~21_combout ) # ((exmem_ifout_o_24)))) # (!\mem_data~22_combout  & (!\mem_data~21_combout  & ((exmem_ifnext_pc_o_24))))

	.dataa(\mem_data~22_combout ),
	.datab(\mem_data~21_combout ),
	.datac(exmem_ifout_o_24),
	.datad(\EXMEM|exmem_if.next_pc_o [24]),
	.cin(gnd),
	.combout(\mem_data~53_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~53 .lut_mask = 16'hB9A8;
defparam \mem_data~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N22
cycloneive_lcell_comb \mem_data~54 (
// Equation(s):
// \mem_data~54_combout  = (\mem_data~21_combout  & ((\mem_data~53_combout  & ((ramiframload_24))) # (!\mem_data~53_combout  & (exmem_ifimm_o_8)))) # (!\mem_data~21_combout  & (\mem_data~53_combout ))

	.dataa(\mem_data~21_combout ),
	.datab(\mem_data~53_combout ),
	.datac(\EXMEM|exmem_if.imm_o [8]),
	.datad(ramiframload_24),
	.cin(gnd),
	.combout(\mem_data~54_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~54 .lut_mask = 16'hEC64;
defparam \mem_data~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N28
cycloneive_lcell_comb \rdat1[24]~49 (
// Equation(s):
// \rdat1[24]~49_combout  = (\rdat1[24]~48_combout ) # ((always03 & \mem_data~54_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(\rdat1[24]~48_combout ),
	.datac(\mem_data~54_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdat1[24]~49_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[24]~49 .lut_mask = 16'hECEC;
defparam \rdat1[24]~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N4
cycloneive_lcell_comb \wdat~52 (
// Equation(s):
// \wdat~52_combout  = (\wdat~18_combout  & (((\wdat~19_combout )))) # (!\wdat~18_combout  & ((\wdat~19_combout  & (memwb_ifnext_pc_o_22)) # (!\wdat~19_combout  & ((memwb_ifout_o_22)))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.next_pc_o [22]),
	.datac(\MEMWB|memwb_if.out_o [22]),
	.datad(\wdat~19_combout ),
	.cin(gnd),
	.combout(\wdat~52_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~52 .lut_mask = 16'hEE50;
defparam \wdat~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N16
cycloneive_lcell_comb \wdat~53 (
// Equation(s):
// \wdat~53_combout  = (\wdat~18_combout  & ((\wdat~52_combout  & (memwb_ifimm_o_6)) # (!\wdat~52_combout  & ((memwb_ifdmemload_o_22))))) # (!\wdat~18_combout  & (\wdat~52_combout ))

	.dataa(\wdat~18_combout ),
	.datab(\wdat~52_combout ),
	.datac(\MEMWB|memwb_if.imm_o [6]),
	.datad(\MEMWB|memwb_if.dmemload_o [22]),
	.cin(gnd),
	.combout(\wdat~53_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~53 .lut_mask = 16'hE6C4;
defparam \wdat~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N4
cycloneive_lcell_comb \rdat1[22]~50 (
// Equation(s):
// \rdat1[22]~50_combout  = (!always03 & ((always02 & ((\wdat~53_combout ))) # (!always02 & (idex_ifrdat1_o_22))))

	.dataa(\FU|always0~11_combout ),
	.datab(\FU|always0~15_combout ),
	.datac(\IDEX|idex_if.rdat1_o [22]),
	.datad(\wdat~53_combout ),
	.cin(gnd),
	.combout(\rdat1[22]~50_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[22]~50 .lut_mask = 16'h3210;
defparam \rdat1[22]~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N22
cycloneive_lcell_comb \mem_data~55 (
// Equation(s):
// \mem_data~55_combout  = (\mem_data~21_combout  & (((\mem_data~22_combout )))) # (!\mem_data~21_combout  & ((\mem_data~22_combout  & ((exmem_ifout_o_22))) # (!\mem_data~22_combout  & (exmem_ifnext_pc_o_22))))

	.dataa(\mem_data~21_combout ),
	.datab(\EXMEM|exmem_if.next_pc_o [22]),
	.datac(\mem_data~22_combout ),
	.datad(exmem_ifout_o_22),
	.cin(gnd),
	.combout(\mem_data~55_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~55 .lut_mask = 16'hF4A4;
defparam \mem_data~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N16
cycloneive_lcell_comb \mem_data~56 (
// Equation(s):
// \mem_data~56_combout  = (\mem_data~21_combout  & ((\mem_data~55_combout  & ((ramiframload_22))) # (!\mem_data~55_combout  & (exmem_ifimm_o_6)))) # (!\mem_data~21_combout  & (((\mem_data~55_combout ))))

	.dataa(\EXMEM|exmem_if.imm_o [6]),
	.datab(\mem_data~21_combout ),
	.datac(\mem_data~55_combout ),
	.datad(ramiframload_22),
	.cin(gnd),
	.combout(\mem_data~56_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~56 .lut_mask = 16'hF838;
defparam \mem_data~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N14
cycloneive_lcell_comb \rdat1[22]~51 (
// Equation(s):
// \rdat1[22]~51_combout  = (\rdat1[22]~50_combout ) # ((always03 & \mem_data~56_combout ))

	.dataa(gnd),
	.datab(\FU|always0~15_combout ),
	.datac(\rdat1[22]~50_combout ),
	.datad(\mem_data~56_combout ),
	.cin(gnd),
	.combout(\rdat1[22]~51_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[22]~51 .lut_mask = 16'hFCF0;
defparam \rdat1[22]~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N10
cycloneive_lcell_comb \wdat~54 (
// Equation(s):
// \wdat~54_combout  = (\wdat~18_combout  & ((memwb_ifdmemload_o_23) # ((\wdat~19_combout )))) # (!\wdat~18_combout  & (((memwb_ifout_o_23 & !\wdat~19_combout ))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.dmemload_o [23]),
	.datac(\MEMWB|memwb_if.out_o [23]),
	.datad(\wdat~19_combout ),
	.cin(gnd),
	.combout(\wdat~54_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~54 .lut_mask = 16'hAAD8;
defparam \wdat~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N26
cycloneive_lcell_comb \wdat~55 (
// Equation(s):
// \wdat~55_combout  = (\wdat~19_combout  & ((\wdat~54_combout  & (memwb_ifimm_o_7)) # (!\wdat~54_combout  & ((memwb_ifnext_pc_o_23))))) # (!\wdat~19_combout  & (((\wdat~54_combout ))))

	.dataa(\wdat~19_combout ),
	.datab(\MEMWB|memwb_if.imm_o [7]),
	.datac(\MEMWB|memwb_if.next_pc_o [23]),
	.datad(\wdat~54_combout ),
	.cin(gnd),
	.combout(\wdat~55_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~55 .lut_mask = 16'hDDA0;
defparam \wdat~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N26
cycloneive_lcell_comb \rdat1[23]~52 (
// Equation(s):
// \rdat1[23]~52_combout  = (!always03 & ((always02 & (\wdat~55_combout )) # (!always02 & ((idex_ifrdat1_o_23)))))

	.dataa(\FU|always0~11_combout ),
	.datab(\wdat~55_combout ),
	.datac(\IDEX|idex_if.rdat1_o [23]),
	.datad(\FU|always0~15_combout ),
	.cin(gnd),
	.combout(\rdat1[23]~52_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[23]~52 .lut_mask = 16'h00D8;
defparam \rdat1[23]~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N12
cycloneive_lcell_comb \mem_data~57 (
// Equation(s):
// \mem_data~57_combout  = (\mem_data~22_combout  & (exmem_ifout_o_23 & ((!\mem_data~21_combout )))) # (!\mem_data~22_combout  & (((exmem_ifnext_pc_o_23) # (\mem_data~21_combout ))))

	.dataa(exmem_ifout_o_23),
	.datab(\mem_data~22_combout ),
	.datac(\EXMEM|exmem_if.next_pc_o [23]),
	.datad(\mem_data~21_combout ),
	.cin(gnd),
	.combout(\mem_data~57_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~57 .lut_mask = 16'h33B8;
defparam \mem_data~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N18
cycloneive_lcell_comb \mem_data~58 (
// Equation(s):
// \mem_data~58_combout  = (\mem_data~57_combout  & (((exmem_ifimm_o_7)) # (!\mem_data~21_combout ))) # (!\mem_data~57_combout  & (\mem_data~21_combout  & ((ramiframload_23))))

	.dataa(\mem_data~57_combout ),
	.datab(\mem_data~21_combout ),
	.datac(\EXMEM|exmem_if.imm_o [7]),
	.datad(ramiframload_23),
	.cin(gnd),
	.combout(\mem_data~58_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~58 .lut_mask = 16'hE6A2;
defparam \mem_data~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N16
cycloneive_lcell_comb \rdat1[23]~53 (
// Equation(s):
// \rdat1[23]~53_combout  = (\rdat1[23]~52_combout ) # ((always03 & \mem_data~58_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(gnd),
	.datac(\rdat1[23]~52_combout ),
	.datad(\mem_data~58_combout ),
	.cin(gnd),
	.combout(\rdat1[23]~53_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[23]~53 .lut_mask = 16'hFAF0;
defparam \rdat1[23]~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N14
cycloneive_lcell_comb \wdat~56 (
// Equation(s):
// \wdat~56_combout  = (\wdat~18_combout  & ((memwb_ifdmemload_o_21) # ((\wdat~19_combout )))) # (!\wdat~18_combout  & (((memwb_ifout_o_21 & !\wdat~19_combout ))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.dmemload_o [21]),
	.datac(\MEMWB|memwb_if.out_o [21]),
	.datad(\wdat~19_combout ),
	.cin(gnd),
	.combout(\wdat~56_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~56 .lut_mask = 16'hAAD8;
defparam \wdat~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N26
cycloneive_lcell_comb \wdat~57 (
// Equation(s):
// \wdat~57_combout  = (\wdat~56_combout  & ((memwb_ifimm_o_5) # ((!\wdat~19_combout )))) # (!\wdat~56_combout  & (((memwb_ifnext_pc_o_21 & \wdat~19_combout ))))

	.dataa(\MEMWB|memwb_if.imm_o [5]),
	.datab(\wdat~56_combout ),
	.datac(\MEMWB|memwb_if.next_pc_o [21]),
	.datad(\wdat~19_combout ),
	.cin(gnd),
	.combout(\wdat~57_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~57 .lut_mask = 16'hB8CC;
defparam \wdat~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N8
cycloneive_lcell_comb \rdat1[21]~54 (
// Equation(s):
// \rdat1[21]~54_combout  = (!always03 & ((always02 & ((\wdat~57_combout ))) # (!always02 & (idex_ifrdat1_o_21))))

	.dataa(\FU|always0~15_combout ),
	.datab(\IDEX|idex_if.rdat1_o [21]),
	.datac(\FU|always0~11_combout ),
	.datad(\wdat~57_combout ),
	.cin(gnd),
	.combout(\rdat1[21]~54_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[21]~54 .lut_mask = 16'h5404;
defparam \rdat1[21]~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N20
cycloneive_lcell_comb \mem_data~59 (
// Equation(s):
// \mem_data~59_combout  = (\mem_data~21_combout  & (((!\mem_data~22_combout )))) # (!\mem_data~21_combout  & ((\mem_data~22_combout  & (exmem_ifout_o_21)) # (!\mem_data~22_combout  & ((exmem_ifnext_pc_o_21)))))

	.dataa(\mem_data~21_combout ),
	.datab(exmem_ifout_o_21),
	.datac(\EXMEM|exmem_if.next_pc_o [21]),
	.datad(\mem_data~22_combout ),
	.cin(gnd),
	.combout(\mem_data~59_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~59 .lut_mask = 16'h44FA;
defparam \mem_data~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N24
cycloneive_lcell_comb \mem_data~60 (
// Equation(s):
// \mem_data~60_combout  = (\mem_data~59_combout  & (((exmem_ifimm_o_5)) # (!\mem_data~21_combout ))) # (!\mem_data~59_combout  & (\mem_data~21_combout  & ((ramiframload_21))))

	.dataa(\mem_data~59_combout ),
	.datab(\mem_data~21_combout ),
	.datac(\EXMEM|exmem_if.imm_o [5]),
	.datad(ramiframload_21),
	.cin(gnd),
	.combout(\mem_data~60_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~60 .lut_mask = 16'hE6A2;
defparam \mem_data~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N14
cycloneive_lcell_comb \rdat1[21]~55 (
// Equation(s):
// \rdat1[21]~55_combout  = (\rdat1[21]~54_combout ) # ((always03 & \mem_data~60_combout ))

	.dataa(\rdat1[21]~54_combout ),
	.datab(gnd),
	.datac(\FU|always0~15_combout ),
	.datad(\mem_data~60_combout ),
	.cin(gnd),
	.combout(\rdat1[21]~55_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[21]~55 .lut_mask = 16'hFAAA;
defparam \rdat1[21]~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N18
cycloneive_lcell_comb \wdat~58 (
// Equation(s):
// \wdat~58_combout  = (\wdat~18_combout  & (((\wdat~19_combout )))) # (!\wdat~18_combout  & ((\wdat~19_combout  & (memwb_ifnext_pc_o_20)) # (!\wdat~19_combout  & ((memwb_ifout_o_20)))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.next_pc_o [20]),
	.datac(\MEMWB|memwb_if.out_o [20]),
	.datad(\wdat~19_combout ),
	.cin(gnd),
	.combout(\wdat~58_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~58 .lut_mask = 16'hEE50;
defparam \wdat~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N30
cycloneive_lcell_comb \wdat~59 (
// Equation(s):
// \wdat~59_combout  = (\wdat~18_combout  & ((\wdat~58_combout  & (memwb_ifimm_o_4)) # (!\wdat~58_combout  & ((memwb_ifdmemload_o_20))))) # (!\wdat~18_combout  & (((\wdat~58_combout ))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.imm_o [4]),
	.datac(\MEMWB|memwb_if.dmemload_o [20]),
	.datad(\wdat~58_combout ),
	.cin(gnd),
	.combout(\wdat~59_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~59 .lut_mask = 16'hDDA0;
defparam \wdat~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N26
cycloneive_lcell_comb \rdat1[20]~56 (
// Equation(s):
// \rdat1[20]~56_combout  = (!always03 & ((always02 & ((\wdat~59_combout ))) # (!always02 & (idex_ifrdat1_o_20))))

	.dataa(\FU|always0~11_combout ),
	.datab(\FU|always0~15_combout ),
	.datac(\IDEX|idex_if.rdat1_o [20]),
	.datad(\wdat~59_combout ),
	.cin(gnd),
	.combout(\rdat1[20]~56_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[20]~56 .lut_mask = 16'h3210;
defparam \rdat1[20]~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N6
cycloneive_lcell_comb \mem_data~61 (
// Equation(s):
// \mem_data~61_combout  = (\mem_data~22_combout  & ((\mem_data~21_combout ) # ((exmem_ifout_o_20)))) # (!\mem_data~22_combout  & (!\mem_data~21_combout  & (exmem_ifnext_pc_o_20)))

	.dataa(\mem_data~22_combout ),
	.datab(\mem_data~21_combout ),
	.datac(\EXMEM|exmem_if.next_pc_o [20]),
	.datad(exmem_ifout_o_20),
	.cin(gnd),
	.combout(\mem_data~61_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~61 .lut_mask = 16'hBA98;
defparam \mem_data~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N24
cycloneive_lcell_comb \mem_data~62 (
// Equation(s):
// \mem_data~62_combout  = (\mem_data~21_combout  & ((\mem_data~61_combout  & ((ramiframload_20))) # (!\mem_data~61_combout  & (exmem_ifimm_o_4)))) # (!\mem_data~21_combout  & (((\mem_data~61_combout ))))

	.dataa(\EXMEM|exmem_if.imm_o [4]),
	.datab(\mem_data~21_combout ),
	.datac(ramiframload_20),
	.datad(\mem_data~61_combout ),
	.cin(gnd),
	.combout(\mem_data~62_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~62 .lut_mask = 16'hF388;
defparam \mem_data~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N20
cycloneive_lcell_comb \rdat1[20]~57 (
// Equation(s):
// \rdat1[20]~57_combout  = (\rdat1[20]~56_combout ) # ((always03 & \mem_data~62_combout ))

	.dataa(gnd),
	.datab(\FU|always0~15_combout ),
	.datac(\rdat1[20]~56_combout ),
	.datad(\mem_data~62_combout ),
	.cin(gnd),
	.combout(\rdat1[20]~57_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[20]~57 .lut_mask = 16'hFCF0;
defparam \rdat1[20]~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N26
cycloneive_lcell_comb \wdat~60 (
// Equation(s):
// \wdat~60_combout  = (\wdat~18_combout  & (((\wdat~19_combout )))) # (!\wdat~18_combout  & ((\wdat~19_combout  & (memwb_ifnext_pc_o_18)) # (!\wdat~19_combout  & ((memwb_ifout_o_18)))))

	.dataa(\wdat~18_combout ),
	.datab(\MEMWB|memwb_if.next_pc_o [18]),
	.datac(\MEMWB|memwb_if.out_o [18]),
	.datad(\wdat~19_combout ),
	.cin(gnd),
	.combout(\wdat~60_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~60 .lut_mask = 16'hEE50;
defparam \wdat~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N6
cycloneive_lcell_comb \wdat~61 (
// Equation(s):
// \wdat~61_combout  = (\wdat~60_combout  & ((memwb_ifimm_o_2) # ((!\wdat~18_combout )))) # (!\wdat~60_combout  & (((memwb_ifdmemload_o_18 & \wdat~18_combout ))))

	.dataa(\wdat~60_combout ),
	.datab(\MEMWB|memwb_if.imm_o [2]),
	.datac(\MEMWB|memwb_if.dmemload_o [18]),
	.datad(\wdat~18_combout ),
	.cin(gnd),
	.combout(\wdat~61_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~61 .lut_mask = 16'hD8AA;
defparam \wdat~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N14
cycloneive_lcell_comb \rdat1[18]~58 (
// Equation(s):
// \rdat1[18]~58_combout  = (!always03 & ((always02 & (\wdat~61_combout )) # (!always02 & ((idex_ifrdat1_o_18)))))

	.dataa(\FU|always0~11_combout ),
	.datab(\FU|always0~15_combout ),
	.datac(\wdat~61_combout ),
	.datad(\IDEX|idex_if.rdat1_o [18]),
	.cin(gnd),
	.combout(\rdat1[18]~58_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[18]~58 .lut_mask = 16'h3120;
defparam \rdat1[18]~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N4
cycloneive_lcell_comb \mem_data~63 (
// Equation(s):
// \mem_data~63_combout  = (\mem_data~21_combout  & (((\mem_data~22_combout )))) # (!\mem_data~21_combout  & ((\mem_data~22_combout  & (exmem_ifout_o_18)) # (!\mem_data~22_combout  & ((exmem_ifnext_pc_o_18)))))

	.dataa(\mem_data~21_combout ),
	.datab(exmem_ifout_o_18),
	.datac(\mem_data~22_combout ),
	.datad(\EXMEM|exmem_if.next_pc_o [18]),
	.cin(gnd),
	.combout(\mem_data~63_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~63 .lut_mask = 16'hE5E0;
defparam \mem_data~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N20
cycloneive_lcell_comb \mem_data~64 (
// Equation(s):
// \mem_data~64_combout  = (\mem_data~63_combout  & (((ramiframload_18)) # (!\mem_data~21_combout ))) # (!\mem_data~63_combout  & (\mem_data~21_combout  & (exmem_ifimm_o_2)))

	.dataa(\mem_data~63_combout ),
	.datab(\mem_data~21_combout ),
	.datac(\EXMEM|exmem_if.imm_o [2]),
	.datad(ramiframload_18),
	.cin(gnd),
	.combout(\mem_data~64_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~64 .lut_mask = 16'hEA62;
defparam \mem_data~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N2
cycloneive_lcell_comb \rdat1[18]~59 (
// Equation(s):
// \rdat1[18]~59_combout  = (\rdat1[18]~58_combout ) # ((always03 & \mem_data~64_combout ))

	.dataa(gnd),
	.datab(\FU|always0~15_combout ),
	.datac(\rdat1[18]~58_combout ),
	.datad(\mem_data~64_combout ),
	.cin(gnd),
	.combout(\rdat1[18]~59_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[18]~59 .lut_mask = 16'hFCF0;
defparam \rdat1[18]~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N12
cycloneive_lcell_comb \wdat~62 (
// Equation(s):
// \wdat~62_combout  = (\wdat~18_combout  & ((memwb_ifdmemload_o_19) # ((\wdat~19_combout )))) # (!\wdat~18_combout  & (((memwb_ifout_o_19 & !\wdat~19_combout ))))

	.dataa(\MEMWB|memwb_if.dmemload_o [19]),
	.datab(\wdat~18_combout ),
	.datac(\MEMWB|memwb_if.out_o [19]),
	.datad(\wdat~19_combout ),
	.cin(gnd),
	.combout(\wdat~62_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~62 .lut_mask = 16'hCCB8;
defparam \wdat~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N4
cycloneive_lcell_comb \wdat~63 (
// Equation(s):
// \wdat~63_combout  = (\wdat~19_combout  & ((\wdat~62_combout  & ((memwb_ifimm_o_3))) # (!\wdat~62_combout  & (memwb_ifnext_pc_o_19)))) # (!\wdat~19_combout  & (((\wdat~62_combout ))))

	.dataa(\MEMWB|memwb_if.next_pc_o [19]),
	.datab(\MEMWB|memwb_if.imm_o [3]),
	.datac(\wdat~19_combout ),
	.datad(\wdat~62_combout ),
	.cin(gnd),
	.combout(\wdat~63_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~63 .lut_mask = 16'hCFA0;
defparam \wdat~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N26
cycloneive_lcell_comb \rdat1[19]~60 (
// Equation(s):
// \rdat1[19]~60_combout  = (!always03 & ((always02 & (\wdat~63_combout )) # (!always02 & ((idex_ifrdat1_o_19)))))

	.dataa(\FU|always0~15_combout ),
	.datab(\wdat~63_combout ),
	.datac(\IDEX|idex_if.rdat1_o [19]),
	.datad(\FU|always0~11_combout ),
	.cin(gnd),
	.combout(\rdat1[19]~60_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[19]~60 .lut_mask = 16'h4450;
defparam \rdat1[19]~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N30
cycloneive_lcell_comb \mem_data~65 (
// Equation(s):
// \mem_data~65_combout  = (\mem_data~22_combout  & (exmem_ifout_o_19 & (!\mem_data~21_combout ))) # (!\mem_data~22_combout  & (((\mem_data~21_combout ) # (exmem_ifnext_pc_o_19))))

	.dataa(\mem_data~22_combout ),
	.datab(exmem_ifout_o_19),
	.datac(\mem_data~21_combout ),
	.datad(\EXMEM|exmem_if.next_pc_o [19]),
	.cin(gnd),
	.combout(\mem_data~65_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~65 .lut_mask = 16'h5D58;
defparam \mem_data~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N12
cycloneive_lcell_comb \mem_data~66 (
// Equation(s):
// \mem_data~66_combout  = (\mem_data~65_combout  & ((exmem_ifimm_o_3) # ((!\mem_data~21_combout )))) # (!\mem_data~65_combout  & (((ramiframload_19 & \mem_data~21_combout ))))

	.dataa(\EXMEM|exmem_if.imm_o [3]),
	.datab(\mem_data~65_combout ),
	.datac(ramiframload_19),
	.datad(\mem_data~21_combout ),
	.cin(gnd),
	.combout(\mem_data~66_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~66 .lut_mask = 16'hB8CC;
defparam \mem_data~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N2
cycloneive_lcell_comb \rdat1[19]~61 (
// Equation(s):
// \rdat1[19]~61_combout  = (\rdat1[19]~60_combout ) # ((always03 & \mem_data~66_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(gnd),
	.datac(\rdat1[19]~60_combout ),
	.datad(\mem_data~66_combout ),
	.cin(gnd),
	.combout(\rdat1[19]~61_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[19]~61 .lut_mask = 16'hFAF0;
defparam \rdat1[19]~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N30
cycloneive_lcell_comb \wdat~64 (
// Equation(s):
// \wdat~64_combout  = (\wdat~19_combout  & (((\wdat~18_combout )))) # (!\wdat~19_combout  & ((\wdat~18_combout  & (memwb_ifdmemload_o_17)) # (!\wdat~18_combout  & ((memwb_ifout_o_17)))))

	.dataa(\wdat~19_combout ),
	.datab(\MEMWB|memwb_if.dmemload_o [17]),
	.datac(\MEMWB|memwb_if.out_o [17]),
	.datad(\wdat~18_combout ),
	.cin(gnd),
	.combout(\wdat~64_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~64 .lut_mask = 16'hEE50;
defparam \wdat~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N22
cycloneive_lcell_comb \wdat~65 (
// Equation(s):
// \wdat~65_combout  = (\wdat~19_combout  & ((\wdat~64_combout  & ((memwb_ifimm_o_1))) # (!\wdat~64_combout  & (memwb_ifnext_pc_o_17)))) # (!\wdat~19_combout  & (((\wdat~64_combout ))))

	.dataa(\MEMWB|memwb_if.next_pc_o [17]),
	.datab(\wdat~19_combout ),
	.datac(\wdat~64_combout ),
	.datad(\MEMWB|memwb_if.imm_o [1]),
	.cin(gnd),
	.combout(\wdat~65_combout ),
	.cout());
// synopsys translate_off
defparam \wdat~65 .lut_mask = 16'hF838;
defparam \wdat~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N14
cycloneive_lcell_comb \rdat1[17]~62 (
// Equation(s):
// \rdat1[17]~62_combout  = (!always03 & ((always02 & (\wdat~65_combout )) # (!always02 & ((idex_ifrdat1_o_17)))))

	.dataa(\FU|always0~15_combout ),
	.datab(\wdat~65_combout ),
	.datac(\FU|always0~11_combout ),
	.datad(\IDEX|idex_if.rdat1_o [17]),
	.cin(gnd),
	.combout(\rdat1[17]~62_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[17]~62 .lut_mask = 16'h4540;
defparam \rdat1[17]~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N8
cycloneive_lcell_comb \mem_data~67 (
// Equation(s):
// \mem_data~67_combout  = (\mem_data~22_combout  & (((!\mem_data~21_combout  & exmem_ifout_o_17)))) # (!\mem_data~22_combout  & ((exmem_ifnext_pc_o_17) # ((\mem_data~21_combout ))))

	.dataa(\EXMEM|exmem_if.next_pc_o [17]),
	.datab(\mem_data~22_combout ),
	.datac(\mem_data~21_combout ),
	.datad(exmem_ifout_o_17),
	.cin(gnd),
	.combout(\mem_data~67_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~67 .lut_mask = 16'h3E32;
defparam \mem_data~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N2
cycloneive_lcell_comb \mem_data~68 (
// Equation(s):
// \mem_data~68_combout  = (\mem_data~67_combout  & (((exmem_ifimm_o_1)) # (!\mem_data~21_combout ))) # (!\mem_data~67_combout  & (\mem_data~21_combout  & ((ramiframload_17))))

	.dataa(\mem_data~67_combout ),
	.datab(\mem_data~21_combout ),
	.datac(\EXMEM|exmem_if.imm_o [1]),
	.datad(ramiframload_17),
	.cin(gnd),
	.combout(\mem_data~68_combout ),
	.cout());
// synopsys translate_off
defparam \mem_data~68 .lut_mask = 16'hE6A2;
defparam \mem_data~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N0
cycloneive_lcell_comb \rdat1[17]~63 (
// Equation(s):
// \rdat1[17]~63_combout  = (\rdat1[17]~62_combout ) # ((always03 & \mem_data~68_combout ))

	.dataa(\FU|always0~15_combout ),
	.datab(\rdat1[17]~62_combout ),
	.datac(gnd),
	.datad(\mem_data~68_combout ),
	.cin(gnd),
	.combout(\rdat1[17]~63_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1[17]~63 .lut_mask = 16'hEECC;
defparam \rdat1[17]~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N2
cycloneive_lcell_comb \port_b~18 (
// Equation(s):
// \port_b~18_combout  = (idex_ifALUSel_o_1 & (!idex_ifALUSel_o_0 & idex_ifimm_o_15))

	.dataa(\IDEX|idex_if.ALUSel_o [1]),
	.datab(\IDEX|idex_if.ALUSel_o [0]),
	.datac(gnd),
	.datad(\IDEX|idex_if.imm_o [15]),
	.cin(gnd),
	.combout(\port_b~18_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~18 .lut_mask = 16'h2200;
defparam \port_b~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N4
cycloneive_lcell_comb \port_b~19 (
// Equation(s):
// \port_b~19_combout  = (\port_b~18_combout ) # ((\port_b~2_combout  & idex_ifrdat2_o_31))

	.dataa(\port_b~2_combout ),
	.datab(gnd),
	.datac(\IDEX|idex_if.rdat2_o [31]),
	.datad(\port_b~18_combout ),
	.cin(gnd),
	.combout(\port_b~19_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~19 .lut_mask = 16'hFFA0;
defparam \port_b~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N6
cycloneive_lcell_comb \port_b~20 (
// Equation(s):
// \port_b~20_combout  = (\port_b~19_combout ) # ((\port_b~0_combout  & fuifrtReplace_31))

	.dataa(\port_b~0_combout ),
	.datab(\port_b~19_combout ),
	.datac(gnd),
	.datad(\FU|fuif.rtReplace[31]~9_combout ),
	.cin(gnd),
	.combout(\port_b~20_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~20 .lut_mask = 16'hEECC;
defparam \port_b~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N22
cycloneive_lcell_comb \port_b~21 (
// Equation(s):
// \port_b~21_combout  = (\port_b~18_combout ) # ((idex_ifrdat2_o_16 & \port_b~2_combout ))

	.dataa(\IDEX|idex_if.rdat2_o [16]),
	.datab(gnd),
	.datac(\port_b~18_combout ),
	.datad(\port_b~2_combout ),
	.cin(gnd),
	.combout(\port_b~21_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~21 .lut_mask = 16'hFAF0;
defparam \port_b~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N10
cycloneive_lcell_comb \port_b~22 (
// Equation(s):
// \port_b~22_combout  = (\port_b~21_combout ) # ((\port_b~0_combout  & fuifrtReplace_16))

	.dataa(gnd),
	.datab(\port_b~0_combout ),
	.datac(\port_b~21_combout ),
	.datad(\FU|fuif.rtReplace[16]~10_combout ),
	.cin(gnd),
	.combout(\port_b~22_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~22 .lut_mask = 16'hFCF0;
defparam \port_b~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N26
cycloneive_lcell_comb \port_b~23 (
// Equation(s):
// \port_b~23_combout  = (\port_b~18_combout ) # ((idex_ifrdat2_o_17 & \port_b~2_combout ))

	.dataa(gnd),
	.datab(\IDEX|idex_if.rdat2_o [17]),
	.datac(\port_b~18_combout ),
	.datad(\port_b~2_combout ),
	.cin(gnd),
	.combout(\port_b~23_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~23 .lut_mask = 16'hFCF0;
defparam \port_b~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N30
cycloneive_lcell_comb \port_b~24 (
// Equation(s):
// \port_b~24_combout  = (\port_b~23_combout ) # ((\port_b~0_combout  & fuifrtReplace_17))

	.dataa(\port_b~0_combout ),
	.datab(gnd),
	.datac(\port_b~23_combout ),
	.datad(\FU|fuif.rtReplace[17]~11_combout ),
	.cin(gnd),
	.combout(\port_b~24_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~24 .lut_mask = 16'hFAF0;
defparam \port_b~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N14
cycloneive_lcell_comb \port_b~25 (
// Equation(s):
// \port_b~25_combout  = (\port_b~18_combout ) # ((idex_ifrdat2_o_18 & \port_b~2_combout ))

	.dataa(gnd),
	.datab(\IDEX|idex_if.rdat2_o [18]),
	.datac(\port_b~18_combout ),
	.datad(\port_b~2_combout ),
	.cin(gnd),
	.combout(\port_b~25_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~25 .lut_mask = 16'hFCF0;
defparam \port_b~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N18
cycloneive_lcell_comb \port_b~26 (
// Equation(s):
// \port_b~26_combout  = (\port_b~25_combout ) # ((\port_b~0_combout  & fuifrtReplace_18))

	.dataa(\port_b~0_combout ),
	.datab(gnd),
	.datac(\port_b~25_combout ),
	.datad(\FU|fuif.rtReplace[18]~12_combout ),
	.cin(gnd),
	.combout(\port_b~26_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~26 .lut_mask = 16'hFAF0;
defparam \port_b~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N28
cycloneive_lcell_comb \port_b~27 (
// Equation(s):
// \port_b~27_combout  = (\port_b~18_combout ) # ((idex_ifrdat2_o_19 & \port_b~2_combout ))

	.dataa(\IDEX|idex_if.rdat2_o [19]),
	.datab(gnd),
	.datac(\port_b~2_combout ),
	.datad(\port_b~18_combout ),
	.cin(gnd),
	.combout(\port_b~27_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~27 .lut_mask = 16'hFFA0;
defparam \port_b~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N10
cycloneive_lcell_comb \port_b~28 (
// Equation(s):
// \port_b~28_combout  = (\port_b~27_combout ) # ((\port_b~0_combout  & fuifrtReplace_19))

	.dataa(\port_b~0_combout ),
	.datab(gnd),
	.datac(\port_b~27_combout ),
	.datad(\FU|fuif.rtReplace[19]~13_combout ),
	.cin(gnd),
	.combout(\port_b~28_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~28 .lut_mask = 16'hFAF0;
defparam \port_b~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N26
cycloneive_lcell_comb \port_b~29 (
// Equation(s):
// \port_b~29_combout  = (\port_b~18_combout ) # ((idex_ifrdat2_o_20 & \port_b~2_combout ))

	.dataa(\IDEX|idex_if.rdat2_o [20]),
	.datab(\port_b~18_combout ),
	.datac(\port_b~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\port_b~29_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~29 .lut_mask = 16'hECEC;
defparam \port_b~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N2
cycloneive_lcell_comb \port_b~30 (
// Equation(s):
// \port_b~30_combout  = (\port_b~29_combout ) # ((\port_b~0_combout  & fuifrtReplace_20))

	.dataa(gnd),
	.datab(\port_b~0_combout ),
	.datac(\port_b~29_combout ),
	.datad(\FU|fuif.rtReplace[20]~14_combout ),
	.cin(gnd),
	.combout(\port_b~30_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~30 .lut_mask = 16'hFCF0;
defparam \port_b~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N6
cycloneive_lcell_comb \port_b~31 (
// Equation(s):
// \port_b~31_combout  = (\port_b~18_combout ) # ((idex_ifrdat2_o_21 & \port_b~2_combout ))

	.dataa(gnd),
	.datab(\IDEX|idex_if.rdat2_o [21]),
	.datac(\port_b~2_combout ),
	.datad(\port_b~18_combout ),
	.cin(gnd),
	.combout(\port_b~31_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~31 .lut_mask = 16'hFFC0;
defparam \port_b~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N18
cycloneive_lcell_comb \port_b~32 (
// Equation(s):
// \port_b~32_combout  = (\port_b~31_combout ) # ((\port_b~0_combout  & fuifrtReplace_21))

	.dataa(\port_b~0_combout ),
	.datab(gnd),
	.datac(\port_b~31_combout ),
	.datad(\FU|fuif.rtReplace[21]~15_combout ),
	.cin(gnd),
	.combout(\port_b~32_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~32 .lut_mask = 16'hFAF0;
defparam \port_b~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N8
cycloneive_lcell_comb \port_b~33 (
// Equation(s):
// \port_b~33_combout  = (\port_b~18_combout ) # ((\port_b~2_combout  & idex_ifrdat2_o_22))

	.dataa(\port_b~18_combout ),
	.datab(\port_b~2_combout ),
	.datac(gnd),
	.datad(\IDEX|idex_if.rdat2_o [22]),
	.cin(gnd),
	.combout(\port_b~33_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~33 .lut_mask = 16'hEEAA;
defparam \port_b~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N12
cycloneive_lcell_comb \port_b~34 (
// Equation(s):
// \port_b~34_combout  = (\port_b~33_combout ) # ((\port_b~0_combout  & fuifrtReplace_22))

	.dataa(gnd),
	.datab(\port_b~0_combout ),
	.datac(\port_b~33_combout ),
	.datad(\FU|fuif.rtReplace[22]~16_combout ),
	.cin(gnd),
	.combout(\port_b~34_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~34 .lut_mask = 16'hFCF0;
defparam \port_b~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N4
cycloneive_lcell_comb \port_b~35 (
// Equation(s):
// \port_b~35_combout  = (\port_b~18_combout ) # ((idex_ifrdat2_o_23 & \port_b~2_combout ))

	.dataa(\IDEX|idex_if.rdat2_o [23]),
	.datab(gnd),
	.datac(\port_b~2_combout ),
	.datad(\port_b~18_combout ),
	.cin(gnd),
	.combout(\port_b~35_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~35 .lut_mask = 16'hFFA0;
defparam \port_b~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N4
cycloneive_lcell_comb \port_b~36 (
// Equation(s):
// \port_b~36_combout  = (\port_b~35_combout ) # ((\port_b~0_combout  & fuifrtReplace_23))

	.dataa(gnd),
	.datab(\port_b~0_combout ),
	.datac(\port_b~35_combout ),
	.datad(\FU|fuif.rtReplace[23]~17_combout ),
	.cin(gnd),
	.combout(\port_b~36_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~36 .lut_mask = 16'hFCF0;
defparam \port_b~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N18
cycloneive_lcell_comb \port_b~37 (
// Equation(s):
// \port_b~37_combout  = (\port_b~18_combout ) # ((\port_b~2_combout  & idex_ifrdat2_o_24))

	.dataa(gnd),
	.datab(\port_b~2_combout ),
	.datac(\port_b~18_combout ),
	.datad(\IDEX|idex_if.rdat2_o [24]),
	.cin(gnd),
	.combout(\port_b~37_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~37 .lut_mask = 16'hFCF0;
defparam \port_b~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N30
cycloneive_lcell_comb \port_b~38 (
// Equation(s):
// \port_b~38_combout  = (\port_b~37_combout ) # ((\port_b~0_combout  & fuifrtReplace_24))

	.dataa(\port_b~0_combout ),
	.datab(\port_b~37_combout ),
	.datac(gnd),
	.datad(\FU|fuif.rtReplace[24]~18_combout ),
	.cin(gnd),
	.combout(\port_b~38_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~38 .lut_mask = 16'hEECC;
defparam \port_b~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N30
cycloneive_lcell_comb \port_b~39 (
// Equation(s):
// \port_b~39_combout  = (\port_b~18_combout ) # ((\port_b~2_combout  & idex_ifrdat2_o_25))

	.dataa(gnd),
	.datab(\port_b~18_combout ),
	.datac(\port_b~2_combout ),
	.datad(\IDEX|idex_if.rdat2_o [25]),
	.cin(gnd),
	.combout(\port_b~39_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~39 .lut_mask = 16'hFCCC;
defparam \port_b~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N8
cycloneive_lcell_comb \port_b~40 (
// Equation(s):
// \port_b~40_combout  = (\port_b~39_combout ) # ((\port_b~0_combout  & fuifrtReplace_25))

	.dataa(gnd),
	.datab(\port_b~0_combout ),
	.datac(\port_b~39_combout ),
	.datad(\FU|fuif.rtReplace[25]~19_combout ),
	.cin(gnd),
	.combout(\port_b~40_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~40 .lut_mask = 16'hFCF0;
defparam \port_b~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N10
cycloneive_lcell_comb \port_b~41 (
// Equation(s):
// \port_b~41_combout  = (\port_b~18_combout ) # ((idex_ifrdat2_o_26 & \port_b~2_combout ))

	.dataa(\IDEX|idex_if.rdat2_o [26]),
	.datab(\port_b~18_combout ),
	.datac(\port_b~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\port_b~41_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~41 .lut_mask = 16'hECEC;
defparam \port_b~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N20
cycloneive_lcell_comb \port_b~42 (
// Equation(s):
// \port_b~42_combout  = (\port_b~41_combout ) # ((\port_b~0_combout  & fuifrtReplace_26))

	.dataa(\port_b~0_combout ),
	.datab(gnd),
	.datac(\port_b~41_combout ),
	.datad(\FU|fuif.rtReplace[26]~20_combout ),
	.cin(gnd),
	.combout(\port_b~42_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~42 .lut_mask = 16'hFAF0;
defparam \port_b~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N26
cycloneive_lcell_comb \port_b~43 (
// Equation(s):
// \port_b~43_combout  = (idex_ifALUSel_o_1 & ((idex_ifimm_o_5) # ((idex_ifrdat2_o_5 & \port_b~2_combout )))) # (!idex_ifALUSel_o_1 & (idex_ifrdat2_o_5 & ((\port_b~2_combout ))))

	.dataa(\IDEX|idex_if.ALUSel_o [1]),
	.datab(\IDEX|idex_if.rdat2_o [5]),
	.datac(\IDEX|idex_if.imm_o [5]),
	.datad(\port_b~2_combout ),
	.cin(gnd),
	.combout(\port_b~43_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~43 .lut_mask = 16'hECA0;
defparam \port_b~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N18
cycloneive_lcell_comb \port_b~44 (
// Equation(s):
// \port_b~44_combout  = (\port_b~43_combout ) # ((\port_b~0_combout  & fuifrtReplace_5))

	.dataa(gnd),
	.datab(\port_b~0_combout ),
	.datac(\port_b~43_combout ),
	.datad(\FU|fuif.rtReplace[5]~21_combout ),
	.cin(gnd),
	.combout(\port_b~44_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~44 .lut_mask = 16'hFCF0;
defparam \port_b~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N28
cycloneive_lcell_comb \port_b~45 (
// Equation(s):
// \port_b~45_combout  = (idex_ifrdat2_o_6 & ((\port_b~2_combout ) # ((idex_ifALUSel_o_1 & idex_ifimm_o_6)))) # (!idex_ifrdat2_o_6 & (idex_ifALUSel_o_1 & (idex_ifimm_o_6)))

	.dataa(\IDEX|idex_if.rdat2_o [6]),
	.datab(\IDEX|idex_if.ALUSel_o [1]),
	.datac(\IDEX|idex_if.imm_o [6]),
	.datad(\port_b~2_combout ),
	.cin(gnd),
	.combout(\port_b~45_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~45 .lut_mask = 16'hEAC0;
defparam \port_b~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N30
cycloneive_lcell_comb \port_b~46 (
// Equation(s):
// \port_b~46_combout  = (\port_b~45_combout ) # ((\port_b~0_combout  & fuifrtReplace_6))

	.dataa(\port_b~0_combout ),
	.datab(gnd),
	.datac(\port_b~45_combout ),
	.datad(\FU|fuif.rtReplace[6]~22_combout ),
	.cin(gnd),
	.combout(\port_b~46_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~46 .lut_mask = 16'hFAF0;
defparam \port_b~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N14
cycloneive_lcell_comb \port_b~47 (
// Equation(s):
// \port_b~47_combout  = (idex_ifALUSel_o_1 & ((idex_ifimm_o_7) # ((idex_ifrdat2_o_7 & \port_b~2_combout )))) # (!idex_ifALUSel_o_1 & (idex_ifrdat2_o_7 & ((\port_b~2_combout ))))

	.dataa(\IDEX|idex_if.ALUSel_o [1]),
	.datab(\IDEX|idex_if.rdat2_o [7]),
	.datac(\IDEX|idex_if.imm_o [7]),
	.datad(\port_b~2_combout ),
	.cin(gnd),
	.combout(\port_b~47_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~47 .lut_mask = 16'hECA0;
defparam \port_b~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N26
cycloneive_lcell_comb \port_b~48 (
// Equation(s):
// \port_b~48_combout  = (\port_b~47_combout ) # ((\port_b~0_combout  & fuifrtReplace_7))

	.dataa(\port_b~0_combout ),
	.datab(gnd),
	.datac(\port_b~47_combout ),
	.datad(\FU|fuif.rtReplace[7]~23_combout ),
	.cin(gnd),
	.combout(\port_b~48_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~48 .lut_mask = 16'hFAF0;
defparam \port_b~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N0
cycloneive_lcell_comb \port_b~49 (
// Equation(s):
// \port_b~49_combout  = (idex_ifimm_o_8 & ((idex_ifALUSel_o_1) # ((idex_ifrdat2_o_8 & \port_b~2_combout )))) # (!idex_ifimm_o_8 & (idex_ifrdat2_o_8 & ((\port_b~2_combout ))))

	.dataa(\IDEX|idex_if.imm_o [8]),
	.datab(\IDEX|idex_if.rdat2_o [8]),
	.datac(\IDEX|idex_if.ALUSel_o [1]),
	.datad(\port_b~2_combout ),
	.cin(gnd),
	.combout(\port_b~49_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~49 .lut_mask = 16'hECA0;
defparam \port_b~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N2
cycloneive_lcell_comb \port_b~50 (
// Equation(s):
// \port_b~50_combout  = (\port_b~49_combout ) # ((\port_b~0_combout  & fuifrtReplace_8))

	.dataa(\port_b~0_combout ),
	.datab(gnd),
	.datac(\port_b~49_combout ),
	.datad(\FU|fuif.rtReplace[8]~24_combout ),
	.cin(gnd),
	.combout(\port_b~50_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~50 .lut_mask = 16'hFAF0;
defparam \port_b~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N16
cycloneive_lcell_comb \port_b~51 (
// Equation(s):
// \port_b~51_combout  = (\port_b~18_combout ) # ((idex_ifrdat2_o_27 & \port_b~2_combout ))

	.dataa(\IDEX|idex_if.rdat2_o [27]),
	.datab(gnd),
	.datac(\port_b~18_combout ),
	.datad(\port_b~2_combout ),
	.cin(gnd),
	.combout(\port_b~51_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~51 .lut_mask = 16'hFAF0;
defparam \port_b~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N24
cycloneive_lcell_comb \port_b~52 (
// Equation(s):
// \port_b~52_combout  = (\port_b~51_combout ) # ((\port_b~0_combout  & fuifrtReplace_27))

	.dataa(gnd),
	.datab(\port_b~0_combout ),
	.datac(\port_b~51_combout ),
	.datad(\FU|fuif.rtReplace[27]~25_combout ),
	.cin(gnd),
	.combout(\port_b~52_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~52 .lut_mask = 16'hFCF0;
defparam \port_b~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N14
cycloneive_lcell_comb \port_b~53 (
// Equation(s):
// \port_b~53_combout  = (\port_b~18_combout ) # ((\port_b~2_combout  & idex_ifrdat2_o_28))

	.dataa(\port_b~18_combout ),
	.datab(gnd),
	.datac(\port_b~2_combout ),
	.datad(\IDEX|idex_if.rdat2_o [28]),
	.cin(gnd),
	.combout(\port_b~53_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~53 .lut_mask = 16'hFAAA;
defparam \port_b~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N10
cycloneive_lcell_comb \port_b~54 (
// Equation(s):
// \port_b~54_combout  = (\port_b~53_combout ) # ((\port_b~0_combout  & fuifrtReplace_28))

	.dataa(\port_b~0_combout ),
	.datab(gnd),
	.datac(\port_b~53_combout ),
	.datad(\FU|fuif.rtReplace[28]~26_combout ),
	.cin(gnd),
	.combout(\port_b~54_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~54 .lut_mask = 16'hFAF0;
defparam \port_b~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N22
cycloneive_lcell_comb \port_b~55 (
// Equation(s):
// \port_b~55_combout  = (\port_b~18_combout ) # ((idex_ifrdat2_o_29 & \port_b~2_combout ))

	.dataa(gnd),
	.datab(\IDEX|idex_if.rdat2_o [29]),
	.datac(\port_b~2_combout ),
	.datad(\port_b~18_combout ),
	.cin(gnd),
	.combout(\port_b~55_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~55 .lut_mask = 16'hFFC0;
defparam \port_b~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N14
cycloneive_lcell_comb \port_b~56 (
// Equation(s):
// \port_b~56_combout  = (\port_b~55_combout ) # ((\port_b~0_combout  & fuifrtReplace_29))

	.dataa(gnd),
	.datab(\port_b~0_combout ),
	.datac(\port_b~55_combout ),
	.datad(\FU|fuif.rtReplace[29]~27_combout ),
	.cin(gnd),
	.combout(\port_b~56_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~56 .lut_mask = 16'hFCF0;
defparam \port_b~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N8
cycloneive_lcell_comb \port_b~57 (
// Equation(s):
// \port_b~57_combout  = (\port_b~18_combout ) # ((idex_ifrdat2_o_30 & \port_b~2_combout ))

	.dataa(\IDEX|idex_if.rdat2_o [30]),
	.datab(gnd),
	.datac(\port_b~2_combout ),
	.datad(\port_b~18_combout ),
	.cin(gnd),
	.combout(\port_b~57_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~57 .lut_mask = 16'hFFA0;
defparam \port_b~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N26
cycloneive_lcell_comb \port_b~58 (
// Equation(s):
// \port_b~58_combout  = (\port_b~57_combout ) # ((\port_b~0_combout  & fuifrtReplace_30))

	.dataa(\port_b~0_combout ),
	.datab(gnd),
	.datac(\port_b~57_combout ),
	.datad(\FU|fuif.rtReplace[30]~28_combout ),
	.cin(gnd),
	.combout(\port_b~58_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~58 .lut_mask = 16'hFAF0;
defparam \port_b~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N10
cycloneive_lcell_comb \port_b~59 (
// Equation(s):
// \port_b~59_combout  = (idex_ifALUSel_o_1 & ((idex_ifimm_o_9) # ((idex_ifrdat2_o_9 & \port_b~2_combout )))) # (!idex_ifALUSel_o_1 & (idex_ifrdat2_o_9 & ((\port_b~2_combout ))))

	.dataa(\IDEX|idex_if.ALUSel_o [1]),
	.datab(\IDEX|idex_if.rdat2_o [9]),
	.datac(\IDEX|idex_if.imm_o [9]),
	.datad(\port_b~2_combout ),
	.cin(gnd),
	.combout(\port_b~59_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~59 .lut_mask = 16'hECA0;
defparam \port_b~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N2
cycloneive_lcell_comb \port_b~60 (
// Equation(s):
// \port_b~60_combout  = (\port_b~59_combout ) # ((\port_b~0_combout  & fuifrtReplace_9))

	.dataa(\port_b~59_combout ),
	.datab(gnd),
	.datac(\port_b~0_combout ),
	.datad(\FU|fuif.rtReplace[9]~29_combout ),
	.cin(gnd),
	.combout(\port_b~60_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~60 .lut_mask = 16'hFAAA;
defparam \port_b~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N18
cycloneive_lcell_comb \port_b~61 (
// Equation(s):
// \port_b~61_combout  = (idex_ifrdat2_o_14 & ((\port_b~2_combout ) # ((idex_ifimm_o_14 & idex_ifALUSel_o_1)))) # (!idex_ifrdat2_o_14 & (idex_ifimm_o_14 & ((idex_ifALUSel_o_1))))

	.dataa(\IDEX|idex_if.rdat2_o [14]),
	.datab(\IDEX|idex_if.imm_o [14]),
	.datac(\port_b~2_combout ),
	.datad(\IDEX|idex_if.ALUSel_o [1]),
	.cin(gnd),
	.combout(\port_b~61_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~61 .lut_mask = 16'hECA0;
defparam \port_b~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N26
cycloneive_lcell_comb \port_b~62 (
// Equation(s):
// \port_b~62_combout  = (idex_ifrdat2_o_15 & ((\port_b~2_combout ) # ((idex_ifimm_o_15 & idex_ifALUSel_o_1)))) # (!idex_ifrdat2_o_15 & (((idex_ifimm_o_15 & idex_ifALUSel_o_1))))

	.dataa(\IDEX|idex_if.rdat2_o [15]),
	.datab(\port_b~2_combout ),
	.datac(\IDEX|idex_if.imm_o [15]),
	.datad(\IDEX|idex_if.ALUSel_o [1]),
	.cin(gnd),
	.combout(\port_b~62_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~62 .lut_mask = 16'hF888;
defparam \port_b~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N16
cycloneive_lcell_comb \port_b~63 (
// Equation(s):
// \port_b~63_combout  = (\port_b~62_combout ) # ((\port_b~0_combout  & fuifrtReplace_15))

	.dataa(gnd),
	.datab(\port_b~0_combout ),
	.datac(\port_b~62_combout ),
	.datad(\FU|fuif.rtReplace[15]~31_combout ),
	.cin(gnd),
	.combout(\port_b~63_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~63 .lut_mask = 16'hFCF0;
defparam \port_b~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N22
cycloneive_lcell_comb \port_b~64 (
// Equation(s):
// \port_b~64_combout  = (idex_ifrdat2_o_10 & ((\port_b~2_combout ) # ((idex_ifimm_o_10 & idex_ifALUSel_o_1)))) # (!idex_ifrdat2_o_10 & (idex_ifimm_o_10 & ((idex_ifALUSel_o_1))))

	.dataa(\IDEX|idex_if.rdat2_o [10]),
	.datab(\IDEX|idex_if.imm_o [10]),
	.datac(\port_b~2_combout ),
	.datad(\IDEX|idex_if.ALUSel_o [1]),
	.cin(gnd),
	.combout(\port_b~64_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~64 .lut_mask = 16'hECA0;
defparam \port_b~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N2
cycloneive_lcell_comb \port_b~65 (
// Equation(s):
// \port_b~65_combout  = (\port_b~64_combout ) # ((\port_b~0_combout  & fuifrtReplace_10))

	.dataa(\port_b~64_combout ),
	.datab(\port_b~0_combout ),
	.datac(gnd),
	.datad(\FU|fuif.rtReplace[10]~32_combout ),
	.cin(gnd),
	.combout(\port_b~65_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~65 .lut_mask = 16'hEEAA;
defparam \port_b~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N0
cycloneive_lcell_comb \port_b~66 (
// Equation(s):
// \port_b~66_combout  = (idex_ifrdat2_o_11 & ((\port_b~2_combout ) # ((idex_ifALUSel_o_1 & idex_ifimm_o_11)))) # (!idex_ifrdat2_o_11 & (idex_ifALUSel_o_1 & ((idex_ifimm_o_11))))

	.dataa(\IDEX|idex_if.rdat2_o [11]),
	.datab(\IDEX|idex_if.ALUSel_o [1]),
	.datac(\port_b~2_combout ),
	.datad(\IDEX|idex_if.imm_o [11]),
	.cin(gnd),
	.combout(\port_b~66_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~66 .lut_mask = 16'hECA0;
defparam \port_b~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N30
cycloneive_lcell_comb \port_b~67 (
// Equation(s):
// \port_b~67_combout  = (\port_b~66_combout ) # ((\port_b~0_combout  & fuifrtReplace_11))

	.dataa(\port_b~0_combout ),
	.datab(gnd),
	.datac(\port_b~66_combout ),
	.datad(\FU|fuif.rtReplace[11]~33_combout ),
	.cin(gnd),
	.combout(\port_b~67_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~67 .lut_mask = 16'hFAF0;
defparam \port_b~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N2
cycloneive_lcell_comb \port_b~68 (
// Equation(s):
// \port_b~68_combout  = (idex_ifrdat2_o_12 & ((\port_b~2_combout ) # ((idex_ifALUSel_o_1 & idex_ifimm_o_12)))) # (!idex_ifrdat2_o_12 & (idex_ifALUSel_o_1 & ((idex_ifimm_o_12))))

	.dataa(\IDEX|idex_if.rdat2_o [12]),
	.datab(\IDEX|idex_if.ALUSel_o [1]),
	.datac(\port_b~2_combout ),
	.datad(\IDEX|idex_if.imm_o [12]),
	.cin(gnd),
	.combout(\port_b~68_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~68 .lut_mask = 16'hECA0;
defparam \port_b~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N26
cycloneive_lcell_comb \port_b~69 (
// Equation(s):
// \port_b~69_combout  = (\port_b~2_combout  & ((idex_ifrdat2_o_13) # ((idex_ifALUSel_o_1 & idex_ifimm_o_13)))) # (!\port_b~2_combout  & (((idex_ifALUSel_o_1 & idex_ifimm_o_13))))

	.dataa(\port_b~2_combout ),
	.datab(\IDEX|idex_if.rdat2_o [13]),
	.datac(\IDEX|idex_if.ALUSel_o [1]),
	.datad(\IDEX|idex_if.imm_o [13]),
	.cin(gnd),
	.combout(\port_b~69_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~69 .lut_mask = 16'hF888;
defparam \port_b~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N20
cycloneive_lcell_comb \port_b~70 (
// Equation(s):
// \port_b~70_combout  = (\port_b~69_combout ) # ((\port_b~0_combout  & fuifrtReplace_13))

	.dataa(gnd),
	.datab(\port_b~0_combout ),
	.datac(\port_b~69_combout ),
	.datad(\FU|fuif.rtReplace[13]~35_combout ),
	.cin(gnd),
	.combout(\port_b~70_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~70 .lut_mask = 16'hFCF0;
defparam \port_b~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N16
cycloneive_lcell_comb \port_b~71 (
// Equation(s):
// \port_b~71_combout  = (\port_b~61_combout ) # ((\port_b~0_combout  & fuifrtReplace_14))

	.dataa(\port_b~0_combout ),
	.datab(gnd),
	.datac(\port_b~61_combout ),
	.datad(\FU|fuif.rtReplace[14]~30_combout ),
	.cin(gnd),
	.combout(\port_b~71_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~71 .lut_mask = 16'hFAF0;
defparam \port_b~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N12
cycloneive_lcell_comb \port_b~72 (
// Equation(s):
// \port_b~72_combout  = (\port_b~68_combout ) # ((\port_b~0_combout  & fuifrtReplace_12))

	.dataa(\port_b~0_combout ),
	.datab(gnd),
	.datac(\FU|fuif.rtReplace[12]~34_combout ),
	.datad(\port_b~68_combout ),
	.cin(gnd),
	.combout(\port_b~72_combout ),
	.cout());
// synopsys translate_off
defparam \port_b~72 .lut_mask = 16'hFFA0;
defparam \port_b~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N29
dffeas \pc[1] (
	.clk(CLK),
	.d(\pc[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pc[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_1),
	.prn(vcc));
// synopsys translate_off
defparam \pc[1] .is_wysiwyg = "true";
defparam \pc[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N31
dffeas \pc[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\new_pc~1_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\pc[1]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_0),
	.prn(vcc));
// synopsys translate_off
defparam \pc[0] .is_wysiwyg = "true";
defparam \pc[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N5
dffeas \pc[3] (
	.clk(CLK),
	.d(\new_pc[3]~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_3),
	.prn(vcc));
// synopsys translate_off
defparam \pc[3] .is_wysiwyg = "true";
defparam \pc[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N27
dffeas \pc[2] (
	.clk(CLK),
	.d(\new_pc[2]~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_2),
	.prn(vcc));
// synopsys translate_off
defparam \pc[2] .is_wysiwyg = "true";
defparam \pc[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y28_N21
dffeas \pc[5] (
	.clk(CLK),
	.d(\new_pc[5]~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_5),
	.prn(vcc));
// synopsys translate_off
defparam \pc[5] .is_wysiwyg = "true";
defparam \pc[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y28_N31
dffeas \pc[4] (
	.clk(CLK),
	.d(\new_pc[4]~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_4),
	.prn(vcc));
// synopsys translate_off
defparam \pc[4] .is_wysiwyg = "true";
defparam \pc[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y29_N29
dffeas \pc[7] (
	.clk(CLK),
	.d(\new_pc[7]~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_7),
	.prn(vcc));
// synopsys translate_off
defparam \pc[7] .is_wysiwyg = "true";
defparam \pc[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y29_N3
dffeas \pc[6] (
	.clk(CLK),
	.d(\new_pc[6]~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_6),
	.prn(vcc));
// synopsys translate_off
defparam \pc[6] .is_wysiwyg = "true";
defparam \pc[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y28_N25
dffeas \pc[9] (
	.clk(CLK),
	.d(\new_pc[9]~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_9),
	.prn(vcc));
// synopsys translate_off
defparam \pc[9] .is_wysiwyg = "true";
defparam \pc[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y28_N3
dffeas \pc[8] (
	.clk(CLK),
	.d(\new_pc[8]~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_8),
	.prn(vcc));
// synopsys translate_off
defparam \pc[8] .is_wysiwyg = "true";
defparam \pc[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N9
dffeas \pc[11] (
	.clk(CLK),
	.d(\new_pc[11]~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_11),
	.prn(vcc));
// synopsys translate_off
defparam \pc[11] .is_wysiwyg = "true";
defparam \pc[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N27
dffeas \pc[10] (
	.clk(CLK),
	.d(\new_pc[10]~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_10),
	.prn(vcc));
// synopsys translate_off
defparam \pc[10] .is_wysiwyg = "true";
defparam \pc[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N17
dffeas \pc[13] (
	.clk(CLK),
	.d(\new_pc[13]~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_13),
	.prn(vcc));
// synopsys translate_off
defparam \pc[13] .is_wysiwyg = "true";
defparam \pc[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N27
dffeas \pc[12] (
	.clk(CLK),
	.d(\new_pc[12]~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_12),
	.prn(vcc));
// synopsys translate_off
defparam \pc[12] .is_wysiwyg = "true";
defparam \pc[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N3
dffeas \pc[15] (
	.clk(CLK),
	.d(\new_pc[15]~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_15),
	.prn(vcc));
// synopsys translate_off
defparam \pc[15] .is_wysiwyg = "true";
defparam \pc[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y28_N13
dffeas \pc[14] (
	.clk(CLK),
	.d(\new_pc[14]~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_14),
	.prn(vcc));
// synopsys translate_off
defparam \pc[14] .is_wysiwyg = "true";
defparam \pc[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N5
dffeas \pc[17] (
	.clk(CLK),
	.d(\new_pc[17]~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_17),
	.prn(vcc));
// synopsys translate_off
defparam \pc[17] .is_wysiwyg = "true";
defparam \pc[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N9
dffeas \pc[16] (
	.clk(CLK),
	.d(\new_pc[16]~33_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_16),
	.prn(vcc));
// synopsys translate_off
defparam \pc[16] .is_wysiwyg = "true";
defparam \pc[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N15
dffeas \pc[19] (
	.clk(CLK),
	.d(\new_pc[19]~35_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_19),
	.prn(vcc));
// synopsys translate_off
defparam \pc[19] .is_wysiwyg = "true";
defparam \pc[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N5
dffeas \pc[18] (
	.clk(CLK),
	.d(\new_pc[18]~37_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_18),
	.prn(vcc));
// synopsys translate_off
defparam \pc[18] .is_wysiwyg = "true";
defparam \pc[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N5
dffeas \pc[21] (
	.clk(CLK),
	.d(\new_pc[21]~39_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_21),
	.prn(vcc));
// synopsys translate_off
defparam \pc[21] .is_wysiwyg = "true";
defparam \pc[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N1
dffeas \pc[20] (
	.clk(CLK),
	.d(\new_pc[20]~41_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_20),
	.prn(vcc));
// synopsys translate_off
defparam \pc[20] .is_wysiwyg = "true";
defparam \pc[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N23
dffeas \pc[23] (
	.clk(CLK),
	.d(\new_pc[23]~43_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_23),
	.prn(vcc));
// synopsys translate_off
defparam \pc[23] .is_wysiwyg = "true";
defparam \pc[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N29
dffeas \pc[22] (
	.clk(CLK),
	.d(\new_pc[22]~45_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_22),
	.prn(vcc));
// synopsys translate_off
defparam \pc[22] .is_wysiwyg = "true";
defparam \pc[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N25
dffeas \pc[25] (
	.clk(CLK),
	.d(\new_pc[25]~47_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_25),
	.prn(vcc));
// synopsys translate_off
defparam \pc[25] .is_wysiwyg = "true";
defparam \pc[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y32_N27
dffeas \pc[24] (
	.clk(CLK),
	.d(\new_pc[24]~49_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_24),
	.prn(vcc));
// synopsys translate_off
defparam \pc[24] .is_wysiwyg = "true";
defparam \pc[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y32_N13
dffeas \pc[27] (
	.clk(CLK),
	.d(\new_pc[27]~51_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_27),
	.prn(vcc));
// synopsys translate_off
defparam \pc[27] .is_wysiwyg = "true";
defparam \pc[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y32_N9
dffeas \pc[26] (
	.clk(CLK),
	.d(\new_pc[26]~53_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_26),
	.prn(vcc));
// synopsys translate_off
defparam \pc[26] .is_wysiwyg = "true";
defparam \pc[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N5
dffeas \pc[29] (
	.clk(CLK),
	.d(\new_pc[29]~55_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_29),
	.prn(vcc));
// synopsys translate_off
defparam \pc[29] .is_wysiwyg = "true";
defparam \pc[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N29
dffeas \pc[28] (
	.clk(CLK),
	.d(\new_pc[28]~57_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_28),
	.prn(vcc));
// synopsys translate_off
defparam \pc[28] .is_wysiwyg = "true";
defparam \pc[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y28_N19
dffeas \pc[31] (
	.clk(CLK),
	.d(\new_pc[31]~59_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_31),
	.prn(vcc));
// synopsys translate_off
defparam \pc[31] .is_wysiwyg = "true";
defparam \pc[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y29_N9
dffeas \pc[30] (
	.clk(CLK),
	.d(\new_pc[30]~61_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_30),
	.prn(vcc));
// synopsys translate_off
defparam \pc[30] .is_wysiwyg = "true";
defparam \pc[30] .power_up = "low";
// synopsys translate_on

// Location: DDIOOUTCELL_X47_Y0_N4
dffeas \dpif.halt (
	.clk(CLK),
	.d(\dpif.halt~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dpifhalt),
	.prn(vcc));
// synopsys translate_off
defparam \dpif.halt .is_wysiwyg = "true";
defparam \dpif.halt .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N4
cycloneive_lcell_comb \new_pc~0 (
// Equation(s):
// \new_pc~0_combout  = (idex_ifjumpSel_o_1 & ((idex_ifjumpSel_o_0 & ((idex_ifnext_pc_o_1))) # (!idex_ifjumpSel_o_0 & (idex_ifrdat1_o_1)))) # (!idex_ifjumpSel_o_1 & (!idex_ifjumpSel_o_0 & ((idex_ifnext_pc_o_1))))

	.dataa(\IDEX|idex_if.jumpSel_o [1]),
	.datab(\IDEX|idex_if.jumpSel_o [0]),
	.datac(\IDEX|idex_if.rdat1_o [1]),
	.datad(\IDEX|idex_if.next_pc_o [1]),
	.cin(gnd),
	.combout(\new_pc~0_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc~0 .lut_mask = 16'hB920;
defparam \new_pc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N28
cycloneive_lcell_comb \pc[1]~feeder (
// Equation(s):
// \pc[1]~feeder_combout  = \new_pc~0_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\new_pc~0_combout ),
	.cin(gnd),
	.combout(\pc[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \pc[1]~feeder .lut_mask = 16'hFF00;
defparam \pc[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N20
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// \always0~0_combout  = (!huiffreeze & always13)

	.dataa(gnd),
	.datab(\HU|huif.freeze~2_combout ),
	.datac(gnd),
	.datad(always13),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'h3300;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N22
cycloneive_lcell_comb \pc[1]~0 (
// Equation(s):
// \pc[1]~0_combout  = (\always0~0_combout  & ((idex_ifjumpSel_o_0 & ((huifflush) # (!idex_ifjumpSel_o_1))) # (!idex_ifjumpSel_o_0 & (idex_ifjumpSel_o_1))))

	.dataa(\IDEX|idex_if.jumpSel_o [0]),
	.datab(\always0~0_combout ),
	.datac(\IDEX|idex_if.jumpSel_o [1]),
	.datad(\HU|huif.flush~0_combout ),
	.cin(gnd),
	.combout(\pc[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \pc[1]~0 .lut_mask = 16'hC848;
defparam \pc[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N20
cycloneive_lcell_comb \new_pc~1 (
// Equation(s):
// \new_pc~1_combout  = (idex_ifjumpSel_o_1 & ((idex_ifjumpSel_o_0 & (idex_ifnext_pc_o_0)) # (!idex_ifjumpSel_o_0 & ((idex_ifrdat1_o_0))))) # (!idex_ifjumpSel_o_1 & (idex_ifnext_pc_o_0 & ((!idex_ifjumpSel_o_0))))

	.dataa(\IDEX|idex_if.jumpSel_o [1]),
	.datab(\IDEX|idex_if.next_pc_o [0]),
	.datac(\IDEX|idex_if.rdat1_o [0]),
	.datad(\IDEX|idex_if.jumpSel_o [0]),
	.cin(gnd),
	.combout(\new_pc~1_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc~1 .lut_mask = 16'h88E4;
defparam \new_pc~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N28
cycloneive_lcell_comb \pc[31]~1 (
// Equation(s):
// \pc[31]~1_combout  = idex_ifjumpSel_o_0 $ (idex_ifjumpSel_o_1)

	.dataa(\IDEX|idex_if.jumpSel_o [0]),
	.datab(gnd),
	.datac(gnd),
	.datad(\IDEX|idex_if.jumpSel_o [1]),
	.cin(gnd),
	.combout(\pc[31]~1_combout ),
	.cout());
// synopsys translate_off
defparam \pc[31]~1 .lut_mask = 16'h55AA;
defparam \pc[31]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N2
cycloneive_lcell_comb \Add1~0 (
// Equation(s):
// \Add1~0_combout  = (idex_ifnext_pc_o_2 & (idex_ifimm_o_0 $ (VCC))) # (!idex_ifnext_pc_o_2 & (idex_ifimm_o_0 & VCC))
// \Add1~1  = CARRY((idex_ifnext_pc_o_2 & idex_ifimm_o_0))

	.dataa(\IDEX|idex_if.next_pc_o [2]),
	.datab(\IDEX|idex_if.imm_o [0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h6688;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N4
cycloneive_lcell_comb \Add1~2 (
// Equation(s):
// \Add1~2_combout  = (idex_ifnext_pc_o_3 & ((idex_ifimm_o_1 & (\Add1~1  & VCC)) # (!idex_ifimm_o_1 & (!\Add1~1 )))) # (!idex_ifnext_pc_o_3 & ((idex_ifimm_o_1 & (!\Add1~1 )) # (!idex_ifimm_o_1 & ((\Add1~1 ) # (GND)))))
// \Add1~3  = CARRY((idex_ifnext_pc_o_3 & (!idex_ifimm_o_1 & !\Add1~1 )) # (!idex_ifnext_pc_o_3 & ((!\Add1~1 ) # (!idex_ifimm_o_1))))

	.dataa(\IDEX|idex_if.next_pc_o [3]),
	.datab(\IDEX|idex_if.imm_o [1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h9617;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N2
cycloneive_lcell_comb \nextpc[2]~0 (
// Equation(s):
// \nextpc[2]~0_combout  = pc_2 $ (VCC)
// \nextpc[2]~1  = CARRY(pc_2)

	.dataa(gnd),
	.datab(pc_2),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\nextpc[2]~0_combout ),
	.cout(\nextpc[2]~1 ));
// synopsys translate_off
defparam \nextpc[2]~0 .lut_mask = 16'h33CC;
defparam \nextpc[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N4
cycloneive_lcell_comb \nextpc[3]~2 (
// Equation(s):
// \nextpc[3]~2_combout  = (pc_3 & (!\nextpc[2]~1 )) # (!pc_3 & ((\nextpc[2]~1 ) # (GND)))
// \nextpc[3]~3  = CARRY((!\nextpc[2]~1 ) # (!pc_3))

	.dataa(gnd),
	.datab(pc_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[2]~1 ),
	.combout(\nextpc[3]~2_combout ),
	.cout(\nextpc[3]~3 ));
// synopsys translate_off
defparam \nextpc[3]~2 .lut_mask = 16'h3C3F;
defparam \nextpc[3]~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N2
cycloneive_lcell_comb \pc[31]~2 (
// Equation(s):
// \pc[31]~2_combout  = (idex_ifjumpSel_o_0 & (((idex_ifPCSel_o & flush)) # (!idex_ifjumpSel_o_1)))

	.dataa(\IDEX|idex_if.jumpSel_o [0]),
	.datab(\IDEX|idex_if.PCSel_o~q ),
	.datac(\IDEX|idex_if.jumpSel_o [1]),
	.datad(\HU|flush~0_combout ),
	.cin(gnd),
	.combout(\pc[31]~2_combout ),
	.cout());
// synopsys translate_off
defparam \pc[31]~2 .lut_mask = 16'h8A0A;
defparam \pc[31]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N20
cycloneive_lcell_comb \new_pc[3]~2 (
// Equation(s):
// \new_pc[3]~2_combout  = (\pc[31]~1_combout  & ((\pc[31]~2_combout  & ((idex_ifimm_26_o_1))) # (!\pc[31]~2_combout  & (idex_ifrdat1_o_3)))) # (!\pc[31]~1_combout  & (((\pc[31]~2_combout ))))

	.dataa(\pc[31]~1_combout ),
	.datab(\IDEX|idex_if.rdat1_o [3]),
	.datac(\IDEX|idex_if.imm_26_o [1]),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[3]~2_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[3]~2 .lut_mask = 16'hF588;
defparam \new_pc[3]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N4
cycloneive_lcell_comb \new_pc[3]~3 (
// Equation(s):
// \new_pc[3]~3_combout  = (\pc[31]~1_combout  & (((\new_pc[3]~2_combout )))) # (!\pc[31]~1_combout  & ((\new_pc[3]~2_combout  & (\Add1~2_combout )) # (!\new_pc[3]~2_combout  & ((\nextpc[3]~2_combout )))))

	.dataa(\pc[31]~1_combout ),
	.datab(\Add1~2_combout ),
	.datac(\nextpc[3]~2_combout ),
	.datad(\new_pc[3]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[3]~3 .lut_mask = 16'hEE50;
defparam \new_pc[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N16
cycloneive_lcell_comb \new_pc[2]~4 (
// Equation(s):
// \new_pc[2]~4_combout  = (\pc[31]~1_combout  & ((idex_ifrdat1_o_2) # ((\pc[31]~2_combout )))) # (!\pc[31]~1_combout  & (((\nextpc[2]~0_combout  & !\pc[31]~2_combout ))))

	.dataa(\pc[31]~1_combout ),
	.datab(\IDEX|idex_if.rdat1_o [2]),
	.datac(\nextpc[2]~0_combout ),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[2]~4_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[2]~4 .lut_mask = 16'hAAD8;
defparam \new_pc[2]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N26
cycloneive_lcell_comb \new_pc[2]~5 (
// Equation(s):
// \new_pc[2]~5_combout  = (\pc[31]~2_combout  & ((\new_pc[2]~4_combout  & (idex_ifimm_26_o_0)) # (!\new_pc[2]~4_combout  & ((\Add1~0_combout ))))) # (!\pc[31]~2_combout  & (((\new_pc[2]~4_combout ))))

	.dataa(\IDEX|idex_if.imm_26_o [0]),
	.datab(\pc[31]~2_combout ),
	.datac(\Add1~0_combout ),
	.datad(\new_pc[2]~4_combout ),
	.cin(gnd),
	.combout(\new_pc[2]~5_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[2]~5 .lut_mask = 16'hBBC0;
defparam \new_pc[2]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N6
cycloneive_lcell_comb \nextpc[4]~4 (
// Equation(s):
// \nextpc[4]~4_combout  = (pc_4 & (\nextpc[3]~3  $ (GND))) # (!pc_4 & (!\nextpc[3]~3  & VCC))
// \nextpc[4]~5  = CARRY((pc_4 & !\nextpc[3]~3 ))

	.dataa(pc_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[3]~3 ),
	.combout(\nextpc[4]~4_combout ),
	.cout(\nextpc[4]~5 ));
// synopsys translate_off
defparam \nextpc[4]~4 .lut_mask = 16'hA50A;
defparam \nextpc[4]~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N8
cycloneive_lcell_comb \nextpc[5]~6 (
// Equation(s):
// \nextpc[5]~6_combout  = (pc_5 & (!\nextpc[4]~5 )) # (!pc_5 & ((\nextpc[4]~5 ) # (GND)))
// \nextpc[5]~7  = CARRY((!\nextpc[4]~5 ) # (!pc_5))

	.dataa(pc_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[4]~5 ),
	.combout(\nextpc[5]~6_combout ),
	.cout(\nextpc[5]~7 ));
// synopsys translate_off
defparam \nextpc[5]~6 .lut_mask = 16'h5A5F;
defparam \nextpc[5]~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N6
cycloneive_lcell_comb \Add1~4 (
// Equation(s):
// \Add1~4_combout  = ((idex_ifnext_pc_o_4 $ (idex_ifimm_o_2 $ (!\Add1~3 )))) # (GND)
// \Add1~5  = CARRY((idex_ifnext_pc_o_4 & ((idex_ifimm_o_2) # (!\Add1~3 ))) # (!idex_ifnext_pc_o_4 & (idex_ifimm_o_2 & !\Add1~3 )))

	.dataa(\IDEX|idex_if.next_pc_o [4]),
	.datab(\IDEX|idex_if.imm_o [2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'h698E;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N8
cycloneive_lcell_comb \Add1~6 (
// Equation(s):
// \Add1~6_combout  = (idex_ifimm_o_3 & ((idex_ifnext_pc_o_5 & (\Add1~5  & VCC)) # (!idex_ifnext_pc_o_5 & (!\Add1~5 )))) # (!idex_ifimm_o_3 & ((idex_ifnext_pc_o_5 & (!\Add1~5 )) # (!idex_ifnext_pc_o_5 & ((\Add1~5 ) # (GND)))))
// \Add1~7  = CARRY((idex_ifimm_o_3 & (!idex_ifnext_pc_o_5 & !\Add1~5 )) # (!idex_ifimm_o_3 & ((!\Add1~5 ) # (!idex_ifnext_pc_o_5))))

	.dataa(\IDEX|idex_if.imm_o [3]),
	.datab(\IDEX|idex_if.next_pc_o [5]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h9617;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N0
cycloneive_lcell_comb \new_pc[5]~6 (
// Equation(s):
// \new_pc[5]~6_combout  = (\pc[31]~1_combout  & ((\pc[31]~2_combout  & (idex_ifimm_26_o_3)) # (!\pc[31]~2_combout  & ((idex_ifrdat1_o_5))))) # (!\pc[31]~1_combout  & (((\pc[31]~2_combout ))))

	.dataa(\IDEX|idex_if.imm_26_o [3]),
	.datab(\pc[31]~1_combout ),
	.datac(\IDEX|idex_if.rdat1_o [5]),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[5]~6_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[5]~6 .lut_mask = 16'hBBC0;
defparam \new_pc[5]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N20
cycloneive_lcell_comb \new_pc[5]~7 (
// Equation(s):
// \new_pc[5]~7_combout  = (\pc[31]~1_combout  & (((\new_pc[5]~6_combout )))) # (!\pc[31]~1_combout  & ((\new_pc[5]~6_combout  & ((\Add1~6_combout ))) # (!\new_pc[5]~6_combout  & (\nextpc[5]~6_combout ))))

	.dataa(\nextpc[5]~6_combout ),
	.datab(\pc[31]~1_combout ),
	.datac(\Add1~6_combout ),
	.datad(\new_pc[5]~6_combout ),
	.cin(gnd),
	.combout(\new_pc[5]~7_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[5]~7 .lut_mask = 16'hFC22;
defparam \new_pc[5]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N6
cycloneive_lcell_comb \new_pc[4]~8 (
// Equation(s):
// \new_pc[4]~8_combout  = (\pc[31]~1_combout  & ((idex_ifrdat1_o_4) # ((\pc[31]~2_combout )))) # (!\pc[31]~1_combout  & (((\nextpc[4]~4_combout  & !\pc[31]~2_combout ))))

	.dataa(\IDEX|idex_if.rdat1_o [4]),
	.datab(\pc[31]~1_combout ),
	.datac(\nextpc[4]~4_combout ),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[4]~8_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[4]~8 .lut_mask = 16'hCCB8;
defparam \new_pc[4]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N30
cycloneive_lcell_comb \new_pc[4]~9 (
// Equation(s):
// \new_pc[4]~9_combout  = (\pc[31]~2_combout  & ((\new_pc[4]~8_combout  & ((idex_ifimm_26_o_2))) # (!\new_pc[4]~8_combout  & (\Add1~4_combout )))) # (!\pc[31]~2_combout  & (((\new_pc[4]~8_combout ))))

	.dataa(\Add1~4_combout ),
	.datab(\IDEX|idex_if.imm_26_o [2]),
	.datac(\pc[31]~2_combout ),
	.datad(\new_pc[4]~8_combout ),
	.cin(gnd),
	.combout(\new_pc[4]~9_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[4]~9 .lut_mask = 16'hCFA0;
defparam \new_pc[4]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N10
cycloneive_lcell_comb \Add1~8 (
// Equation(s):
// \Add1~8_combout  = ((idex_ifnext_pc_o_6 $ (idex_ifimm_o_4 $ (!\Add1~7 )))) # (GND)
// \Add1~9  = CARRY((idex_ifnext_pc_o_6 & ((idex_ifimm_o_4) # (!\Add1~7 ))) # (!idex_ifnext_pc_o_6 & (idex_ifimm_o_4 & !\Add1~7 )))

	.dataa(\IDEX|idex_if.next_pc_o [6]),
	.datab(\IDEX|idex_if.imm_o [4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'h698E;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N12
cycloneive_lcell_comb \Add1~10 (
// Equation(s):
// \Add1~10_combout  = (idex_ifnext_pc_o_7 & ((idex_ifimm_o_5 & (\Add1~9  & VCC)) # (!idex_ifimm_o_5 & (!\Add1~9 )))) # (!idex_ifnext_pc_o_7 & ((idex_ifimm_o_5 & (!\Add1~9 )) # (!idex_ifimm_o_5 & ((\Add1~9 ) # (GND)))))
// \Add1~11  = CARRY((idex_ifnext_pc_o_7 & (!idex_ifimm_o_5 & !\Add1~9 )) # (!idex_ifnext_pc_o_7 & ((!\Add1~9 ) # (!idex_ifimm_o_5))))

	.dataa(\IDEX|idex_if.next_pc_o [7]),
	.datab(\IDEX|idex_if.imm_o [5]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h9617;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N10
cycloneive_lcell_comb \nextpc[6]~8 (
// Equation(s):
// \nextpc[6]~8_combout  = (pc_6 & (\nextpc[5]~7  $ (GND))) # (!pc_6 & (!\nextpc[5]~7  & VCC))
// \nextpc[6]~9  = CARRY((pc_6 & !\nextpc[5]~7 ))

	.dataa(gnd),
	.datab(pc_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[5]~7 ),
	.combout(\nextpc[6]~8_combout ),
	.cout(\nextpc[6]~9 ));
// synopsys translate_off
defparam \nextpc[6]~8 .lut_mask = 16'hC30C;
defparam \nextpc[6]~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N12
cycloneive_lcell_comb \nextpc[7]~10 (
// Equation(s):
// \nextpc[7]~10_combout  = (pc_7 & (!\nextpc[6]~9 )) # (!pc_7 & ((\nextpc[6]~9 ) # (GND)))
// \nextpc[7]~11  = CARRY((!\nextpc[6]~9 ) # (!pc_7))

	.dataa(gnd),
	.datab(pc_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[6]~9 ),
	.combout(\nextpc[7]~10_combout ),
	.cout(\nextpc[7]~11 ));
// synopsys translate_off
defparam \nextpc[7]~10 .lut_mask = 16'h3C3F;
defparam \nextpc[7]~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N12
cycloneive_lcell_comb \new_pc[7]~10 (
// Equation(s):
// \new_pc[7]~10_combout  = (\pc[31]~1_combout  & ((\pc[31]~2_combout  & ((idex_ifimm_26_o_5))) # (!\pc[31]~2_combout  & (idex_ifrdat1_o_7)))) # (!\pc[31]~1_combout  & (((\pc[31]~2_combout ))))

	.dataa(\IDEX|idex_if.rdat1_o [7]),
	.datab(\pc[31]~1_combout ),
	.datac(\IDEX|idex_if.imm_26_o [5]),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[7]~10_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[7]~10 .lut_mask = 16'hF388;
defparam \new_pc[7]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N28
cycloneive_lcell_comb \new_pc[7]~11 (
// Equation(s):
// \new_pc[7]~11_combout  = (\pc[31]~1_combout  & (((\new_pc[7]~10_combout )))) # (!\pc[31]~1_combout  & ((\new_pc[7]~10_combout  & (\Add1~10_combout )) # (!\new_pc[7]~10_combout  & ((\nextpc[7]~10_combout )))))

	.dataa(\Add1~10_combout ),
	.datab(\pc[31]~1_combout ),
	.datac(\nextpc[7]~10_combout ),
	.datad(\new_pc[7]~10_combout ),
	.cin(gnd),
	.combout(\new_pc[7]~11_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[7]~11 .lut_mask = 16'hEE30;
defparam \new_pc[7]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N10
cycloneive_lcell_comb \new_pc[6]~12 (
// Equation(s):
// \new_pc[6]~12_combout  = (\pc[31]~1_combout  & ((idex_ifrdat1_o_6) # ((\pc[31]~2_combout )))) # (!\pc[31]~1_combout  & (((\nextpc[6]~8_combout  & !\pc[31]~2_combout ))))

	.dataa(\IDEX|idex_if.rdat1_o [6]),
	.datab(\pc[31]~1_combout ),
	.datac(\nextpc[6]~8_combout ),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[6]~12_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[6]~12 .lut_mask = 16'hCCB8;
defparam \new_pc[6]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N2
cycloneive_lcell_comb \new_pc[6]~13 (
// Equation(s):
// \new_pc[6]~13_combout  = (\pc[31]~2_combout  & ((\new_pc[6]~12_combout  & (idex_ifimm_26_o_4)) # (!\new_pc[6]~12_combout  & ((\Add1~8_combout ))))) # (!\pc[31]~2_combout  & (((\new_pc[6]~12_combout ))))

	.dataa(\IDEX|idex_if.imm_26_o [4]),
	.datab(\Add1~8_combout ),
	.datac(\pc[31]~2_combout ),
	.datad(\new_pc[6]~12_combout ),
	.cin(gnd),
	.combout(\new_pc[6]~13_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[6]~13 .lut_mask = 16'hAFC0;
defparam \new_pc[6]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N14
cycloneive_lcell_comb \nextpc[8]~12 (
// Equation(s):
// \nextpc[8]~12_combout  = (pc_8 & (\nextpc[7]~11  $ (GND))) # (!pc_8 & (!\nextpc[7]~11  & VCC))
// \nextpc[8]~13  = CARRY((pc_8 & !\nextpc[7]~11 ))

	.dataa(gnd),
	.datab(pc_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[7]~11 ),
	.combout(\nextpc[8]~12_combout ),
	.cout(\nextpc[8]~13 ));
// synopsys translate_off
defparam \nextpc[8]~12 .lut_mask = 16'hC30C;
defparam \nextpc[8]~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N16
cycloneive_lcell_comb \nextpc[9]~14 (
// Equation(s):
// \nextpc[9]~14_combout  = (pc_9 & (!\nextpc[8]~13 )) # (!pc_9 & ((\nextpc[8]~13 ) # (GND)))
// \nextpc[9]~15  = CARRY((!\nextpc[8]~13 ) # (!pc_9))

	.dataa(pc_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[8]~13 ),
	.combout(\nextpc[9]~14_combout ),
	.cout(\nextpc[9]~15 ));
// synopsys translate_off
defparam \nextpc[9]~14 .lut_mask = 16'h5A5F;
defparam \nextpc[9]~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N14
cycloneive_lcell_comb \Add1~12 (
// Equation(s):
// \Add1~12_combout  = ((idex_ifimm_o_6 $ (idex_ifnext_pc_o_8 $ (!\Add1~11 )))) # (GND)
// \Add1~13  = CARRY((idex_ifimm_o_6 & ((idex_ifnext_pc_o_8) # (!\Add1~11 ))) # (!idex_ifimm_o_6 & (idex_ifnext_pc_o_8 & !\Add1~11 )))

	.dataa(\IDEX|idex_if.imm_o [6]),
	.datab(\IDEX|idex_if.next_pc_o [8]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout(\Add1~13 ));
// synopsys translate_off
defparam \Add1~12 .lut_mask = 16'h698E;
defparam \Add1~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N16
cycloneive_lcell_comb \Add1~14 (
// Equation(s):
// \Add1~14_combout  = (idex_ifimm_o_7 & ((idex_ifnext_pc_o_9 & (\Add1~13  & VCC)) # (!idex_ifnext_pc_o_9 & (!\Add1~13 )))) # (!idex_ifimm_o_7 & ((idex_ifnext_pc_o_9 & (!\Add1~13 )) # (!idex_ifnext_pc_o_9 & ((\Add1~13 ) # (GND)))))
// \Add1~15  = CARRY((idex_ifimm_o_7 & (!idex_ifnext_pc_o_9 & !\Add1~13 )) # (!idex_ifimm_o_7 & ((!\Add1~13 ) # (!idex_ifnext_pc_o_9))))

	.dataa(\IDEX|idex_if.imm_o [7]),
	.datab(\IDEX|idex_if.next_pc_o [9]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~13 ),
	.combout(\Add1~14_combout ),
	.cout(\Add1~15 ));
// synopsys translate_off
defparam \Add1~14 .lut_mask = 16'h9617;
defparam \Add1~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N16
cycloneive_lcell_comb \new_pc[9]~14 (
// Equation(s):
// \new_pc[9]~14_combout  = (\pc[31]~1_combout  & ((\pc[31]~2_combout  & (idex_ifimm_26_o_7)) # (!\pc[31]~2_combout  & ((idex_ifrdat1_o_9))))) # (!\pc[31]~1_combout  & (((\pc[31]~2_combout ))))

	.dataa(\pc[31]~1_combout ),
	.datab(\IDEX|idex_if.imm_26_o [7]),
	.datac(\pc[31]~2_combout ),
	.datad(\IDEX|idex_if.rdat1_o [9]),
	.cin(gnd),
	.combout(\new_pc[9]~14_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[9]~14 .lut_mask = 16'hDAD0;
defparam \new_pc[9]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N24
cycloneive_lcell_comb \new_pc[9]~15 (
// Equation(s):
// \new_pc[9]~15_combout  = (\pc[31]~1_combout  & (((\new_pc[9]~14_combout )))) # (!\pc[31]~1_combout  & ((\new_pc[9]~14_combout  & ((\Add1~14_combout ))) # (!\new_pc[9]~14_combout  & (\nextpc[9]~14_combout ))))

	.dataa(\pc[31]~1_combout ),
	.datab(\nextpc[9]~14_combout ),
	.datac(\Add1~14_combout ),
	.datad(\new_pc[9]~14_combout ),
	.cin(gnd),
	.combout(\new_pc[9]~15_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[9]~15 .lut_mask = 16'hFA44;
defparam \new_pc[9]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N22
cycloneive_lcell_comb \new_pc[8]~16 (
// Equation(s):
// \new_pc[8]~16_combout  = (\pc[31]~1_combout  & (((\pc[31]~2_combout ) # (idex_ifrdat1_o_8)))) # (!\pc[31]~1_combout  & (\nextpc[8]~12_combout  & (!\pc[31]~2_combout )))

	.dataa(\pc[31]~1_combout ),
	.datab(\nextpc[8]~12_combout ),
	.datac(\pc[31]~2_combout ),
	.datad(\IDEX|idex_if.rdat1_o [8]),
	.cin(gnd),
	.combout(\new_pc[8]~16_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[8]~16 .lut_mask = 16'hAEA4;
defparam \new_pc[8]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N2
cycloneive_lcell_comb \new_pc[8]~17 (
// Equation(s):
// \new_pc[8]~17_combout  = (\pc[31]~2_combout  & ((\new_pc[8]~16_combout  & (idex_ifimm_26_o_6)) # (!\new_pc[8]~16_combout  & ((\Add1~12_combout ))))) # (!\pc[31]~2_combout  & (((\new_pc[8]~16_combout ))))

	.dataa(\IDEX|idex_if.imm_26_o [6]),
	.datab(\pc[31]~2_combout ),
	.datac(\new_pc[8]~16_combout ),
	.datad(\Add1~12_combout ),
	.cin(gnd),
	.combout(\new_pc[8]~17_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[8]~17 .lut_mask = 16'hBCB0;
defparam \new_pc[8]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N18
cycloneive_lcell_comb \nextpc[10]~16 (
// Equation(s):
// \nextpc[10]~16_combout  = (pc_10 & (\nextpc[9]~15  $ (GND))) # (!pc_10 & (!\nextpc[9]~15  & VCC))
// \nextpc[10]~17  = CARRY((pc_10 & !\nextpc[9]~15 ))

	.dataa(gnd),
	.datab(pc_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[9]~15 ),
	.combout(\nextpc[10]~16_combout ),
	.cout(\nextpc[10]~17 ));
// synopsys translate_off
defparam \nextpc[10]~16 .lut_mask = 16'hC30C;
defparam \nextpc[10]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N20
cycloneive_lcell_comb \nextpc[11]~18 (
// Equation(s):
// \nextpc[11]~18_combout  = (pc_11 & (!\nextpc[10]~17 )) # (!pc_11 & ((\nextpc[10]~17 ) # (GND)))
// \nextpc[11]~19  = CARRY((!\nextpc[10]~17 ) # (!pc_11))

	.dataa(pc_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[10]~17 ),
	.combout(\nextpc[11]~18_combout ),
	.cout(\nextpc[11]~19 ));
// synopsys translate_off
defparam \nextpc[11]~18 .lut_mask = 16'h5A5F;
defparam \nextpc[11]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N18
cycloneive_lcell_comb \Add1~16 (
// Equation(s):
// \Add1~16_combout  = ((idex_ifimm_o_8 $ (idex_ifnext_pc_o_10 $ (!\Add1~15 )))) # (GND)
// \Add1~17  = CARRY((idex_ifimm_o_8 & ((idex_ifnext_pc_o_10) # (!\Add1~15 ))) # (!idex_ifimm_o_8 & (idex_ifnext_pc_o_10 & !\Add1~15 )))

	.dataa(\IDEX|idex_if.imm_o [8]),
	.datab(\IDEX|idex_if.next_pc_o [10]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~15 ),
	.combout(\Add1~16_combout ),
	.cout(\Add1~17 ));
// synopsys translate_off
defparam \Add1~16 .lut_mask = 16'h698E;
defparam \Add1~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N20
cycloneive_lcell_comb \Add1~18 (
// Equation(s):
// \Add1~18_combout  = (idex_ifimm_o_9 & ((idex_ifnext_pc_o_11 & (\Add1~17  & VCC)) # (!idex_ifnext_pc_o_11 & (!\Add1~17 )))) # (!idex_ifimm_o_9 & ((idex_ifnext_pc_o_11 & (!\Add1~17 )) # (!idex_ifnext_pc_o_11 & ((\Add1~17 ) # (GND)))))
// \Add1~19  = CARRY((idex_ifimm_o_9 & (!idex_ifnext_pc_o_11 & !\Add1~17 )) # (!idex_ifimm_o_9 & ((!\Add1~17 ) # (!idex_ifnext_pc_o_11))))

	.dataa(\IDEX|idex_if.imm_o [9]),
	.datab(\IDEX|idex_if.next_pc_o [11]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~17 ),
	.combout(\Add1~18_combout ),
	.cout(\Add1~19 ));
// synopsys translate_off
defparam \Add1~18 .lut_mask = 16'h9617;
defparam \Add1~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N18
cycloneive_lcell_comb \new_pc[11]~18 (
// Equation(s):
// \new_pc[11]~18_combout  = (\pc[31]~1_combout  & ((\pc[31]~2_combout  & (idex_ifimm_26_o_9)) # (!\pc[31]~2_combout  & ((idex_ifrdat1_o_11))))) # (!\pc[31]~1_combout  & (((\pc[31]~2_combout ))))

	.dataa(\IDEX|idex_if.imm_26_o [9]),
	.datab(\pc[31]~1_combout ),
	.datac(\IDEX|idex_if.rdat1_o [11]),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[11]~18_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[11]~18 .lut_mask = 16'hBBC0;
defparam \new_pc[11]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N8
cycloneive_lcell_comb \new_pc[11]~19 (
// Equation(s):
// \new_pc[11]~19_combout  = (\pc[31]~1_combout  & (((\new_pc[11]~18_combout )))) # (!\pc[31]~1_combout  & ((\new_pc[11]~18_combout  & ((\Add1~18_combout ))) # (!\new_pc[11]~18_combout  & (\nextpc[11]~18_combout ))))

	.dataa(\nextpc[11]~18_combout ),
	.datab(\pc[31]~1_combout ),
	.datac(\Add1~18_combout ),
	.datad(\new_pc[11]~18_combout ),
	.cin(gnd),
	.combout(\new_pc[11]~19_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[11]~19 .lut_mask = 16'hFC22;
defparam \new_pc[11]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N4
cycloneive_lcell_comb \new_pc[10]~20 (
// Equation(s):
// \new_pc[10]~20_combout  = (\pc[31]~1_combout  & ((idex_ifrdat1_o_10) # ((\pc[31]~2_combout )))) # (!\pc[31]~1_combout  & (((\nextpc[10]~16_combout  & !\pc[31]~2_combout ))))

	.dataa(\IDEX|idex_if.rdat1_o [10]),
	.datab(\pc[31]~1_combout ),
	.datac(\nextpc[10]~16_combout ),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[10]~20_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[10]~20 .lut_mask = 16'hCCB8;
defparam \new_pc[10]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N26
cycloneive_lcell_comb \new_pc[10]~21 (
// Equation(s):
// \new_pc[10]~21_combout  = (\new_pc[10]~20_combout  & ((idex_ifimm_26_o_8) # ((!\pc[31]~2_combout )))) # (!\new_pc[10]~20_combout  & (((\Add1~16_combout  & \pc[31]~2_combout ))))

	.dataa(\IDEX|idex_if.imm_26_o [8]),
	.datab(\Add1~16_combout ),
	.datac(\new_pc[10]~20_combout ),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[10]~21_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[10]~21 .lut_mask = 16'hACF0;
defparam \new_pc[10]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N22
cycloneive_lcell_comb \Add1~20 (
// Equation(s):
// \Add1~20_combout  = ((idex_ifimm_o_10 $ (idex_ifnext_pc_o_12 $ (!\Add1~19 )))) # (GND)
// \Add1~21  = CARRY((idex_ifimm_o_10 & ((idex_ifnext_pc_o_12) # (!\Add1~19 ))) # (!idex_ifimm_o_10 & (idex_ifnext_pc_o_12 & !\Add1~19 )))

	.dataa(\IDEX|idex_if.imm_o [10]),
	.datab(\IDEX|idex_if.next_pc_o [12]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~19 ),
	.combout(\Add1~20_combout ),
	.cout(\Add1~21 ));
// synopsys translate_off
defparam \Add1~20 .lut_mask = 16'h698E;
defparam \Add1~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N24
cycloneive_lcell_comb \Add1~22 (
// Equation(s):
// \Add1~22_combout  = (idex_ifimm_o_11 & ((idex_ifnext_pc_o_13 & (\Add1~21  & VCC)) # (!idex_ifnext_pc_o_13 & (!\Add1~21 )))) # (!idex_ifimm_o_11 & ((idex_ifnext_pc_o_13 & (!\Add1~21 )) # (!idex_ifnext_pc_o_13 & ((\Add1~21 ) # (GND)))))
// \Add1~23  = CARRY((idex_ifimm_o_11 & (!idex_ifnext_pc_o_13 & !\Add1~21 )) # (!idex_ifimm_o_11 & ((!\Add1~21 ) # (!idex_ifnext_pc_o_13))))

	.dataa(\IDEX|idex_if.imm_o [11]),
	.datab(\IDEX|idex_if.next_pc_o [13]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~21 ),
	.combout(\Add1~22_combout ),
	.cout(\Add1~23 ));
// synopsys translate_off
defparam \Add1~22 .lut_mask = 16'h9617;
defparam \Add1~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N22
cycloneive_lcell_comb \nextpc[12]~20 (
// Equation(s):
// \nextpc[12]~20_combout  = (pc_12 & (\nextpc[11]~19  $ (GND))) # (!pc_12 & (!\nextpc[11]~19  & VCC))
// \nextpc[12]~21  = CARRY((pc_12 & !\nextpc[11]~19 ))

	.dataa(pc_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[11]~19 ),
	.combout(\nextpc[12]~20_combout ),
	.cout(\nextpc[12]~21 ));
// synopsys translate_off
defparam \nextpc[12]~20 .lut_mask = 16'hA50A;
defparam \nextpc[12]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N24
cycloneive_lcell_comb \nextpc[13]~22 (
// Equation(s):
// \nextpc[13]~22_combout  = (pc_13 & (!\nextpc[12]~21 )) # (!pc_13 & ((\nextpc[12]~21 ) # (GND)))
// \nextpc[13]~23  = CARRY((!\nextpc[12]~21 ) # (!pc_13))

	.dataa(pc_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[12]~21 ),
	.combout(\nextpc[13]~22_combout ),
	.cout(\nextpc[13]~23 ));
// synopsys translate_off
defparam \nextpc[13]~22 .lut_mask = 16'h5A5F;
defparam \nextpc[13]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N20
cycloneive_lcell_comb \new_pc[13]~22 (
// Equation(s):
// \new_pc[13]~22_combout  = (\pc[31]~1_combout  & ((\pc[31]~2_combout  & ((idex_ifimm_26_o_11))) # (!\pc[31]~2_combout  & (idex_ifrdat1_o_13)))) # (!\pc[31]~1_combout  & (((\pc[31]~2_combout ))))

	.dataa(\pc[31]~1_combout ),
	.datab(\IDEX|idex_if.rdat1_o [13]),
	.datac(\IDEX|idex_if.imm_26_o [11]),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[13]~22_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[13]~22 .lut_mask = 16'hF588;
defparam \new_pc[13]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N16
cycloneive_lcell_comb \new_pc[13]~23 (
// Equation(s):
// \new_pc[13]~23_combout  = (\pc[31]~1_combout  & (((\new_pc[13]~22_combout )))) # (!\pc[31]~1_combout  & ((\new_pc[13]~22_combout  & (\Add1~22_combout )) # (!\new_pc[13]~22_combout  & ((\nextpc[13]~22_combout )))))

	.dataa(\pc[31]~1_combout ),
	.datab(\Add1~22_combout ),
	.datac(\nextpc[13]~22_combout ),
	.datad(\new_pc[13]~22_combout ),
	.cin(gnd),
	.combout(\new_pc[13]~23_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[13]~23 .lut_mask = 16'hEE50;
defparam \new_pc[13]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N22
cycloneive_lcell_comb \new_pc[12]~24 (
// Equation(s):
// \new_pc[12]~24_combout  = (\pc[31]~1_combout  & ((idex_ifrdat1_o_12) # ((\pc[31]~2_combout )))) # (!\pc[31]~1_combout  & (((!\pc[31]~2_combout  & \nextpc[12]~20_combout ))))

	.dataa(\IDEX|idex_if.rdat1_o [12]),
	.datab(\pc[31]~1_combout ),
	.datac(\pc[31]~2_combout ),
	.datad(\nextpc[12]~20_combout ),
	.cin(gnd),
	.combout(\new_pc[12]~24_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[12]~24 .lut_mask = 16'hCBC8;
defparam \new_pc[12]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N26
cycloneive_lcell_comb \new_pc[12]~25 (
// Equation(s):
// \new_pc[12]~25_combout  = (\pc[31]~2_combout  & ((\new_pc[12]~24_combout  & ((idex_ifimm_26_o_10))) # (!\new_pc[12]~24_combout  & (\Add1~20_combout )))) # (!\pc[31]~2_combout  & (((\new_pc[12]~24_combout ))))

	.dataa(\Add1~20_combout ),
	.datab(\IDEX|idex_if.imm_26_o [10]),
	.datac(\pc[31]~2_combout ),
	.datad(\new_pc[12]~24_combout ),
	.cin(gnd),
	.combout(\new_pc[12]~25_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[12]~25 .lut_mask = 16'hCFA0;
defparam \new_pc[12]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N26
cycloneive_lcell_comb \nextpc[14]~24 (
// Equation(s):
// \nextpc[14]~24_combout  = (pc_14 & (\nextpc[13]~23  $ (GND))) # (!pc_14 & (!\nextpc[13]~23  & VCC))
// \nextpc[14]~25  = CARRY((pc_14 & !\nextpc[13]~23 ))

	.dataa(gnd),
	.datab(pc_14),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[13]~23 ),
	.combout(\nextpc[14]~24_combout ),
	.cout(\nextpc[14]~25 ));
// synopsys translate_off
defparam \nextpc[14]~24 .lut_mask = 16'hC30C;
defparam \nextpc[14]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N28
cycloneive_lcell_comb \nextpc[15]~26 (
// Equation(s):
// \nextpc[15]~26_combout  = (pc_15 & (!\nextpc[14]~25 )) # (!pc_15 & ((\nextpc[14]~25 ) # (GND)))
// \nextpc[15]~27  = CARRY((!\nextpc[14]~25 ) # (!pc_15))

	.dataa(pc_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[14]~25 ),
	.combout(\nextpc[15]~26_combout ),
	.cout(\nextpc[15]~27 ));
// synopsys translate_off
defparam \nextpc[15]~26 .lut_mask = 16'h5A5F;
defparam \nextpc[15]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N26
cycloneive_lcell_comb \Add1~24 (
// Equation(s):
// \Add1~24_combout  = ((idex_ifnext_pc_o_14 $ (idex_ifimm_o_12 $ (!\Add1~23 )))) # (GND)
// \Add1~25  = CARRY((idex_ifnext_pc_o_14 & ((idex_ifimm_o_12) # (!\Add1~23 ))) # (!idex_ifnext_pc_o_14 & (idex_ifimm_o_12 & !\Add1~23 )))

	.dataa(\IDEX|idex_if.next_pc_o [14]),
	.datab(\IDEX|idex_if.imm_o [12]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~23 ),
	.combout(\Add1~24_combout ),
	.cout(\Add1~25 ));
// synopsys translate_off
defparam \Add1~24 .lut_mask = 16'h698E;
defparam \Add1~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N28
cycloneive_lcell_comb \Add1~26 (
// Equation(s):
// \Add1~26_combout  = (idex_ifimm_o_13 & ((idex_ifnext_pc_o_15 & (\Add1~25  & VCC)) # (!idex_ifnext_pc_o_15 & (!\Add1~25 )))) # (!idex_ifimm_o_13 & ((idex_ifnext_pc_o_15 & (!\Add1~25 )) # (!idex_ifnext_pc_o_15 & ((\Add1~25 ) # (GND)))))
// \Add1~27  = CARRY((idex_ifimm_o_13 & (!idex_ifnext_pc_o_15 & !\Add1~25 )) # (!idex_ifimm_o_13 & ((!\Add1~25 ) # (!idex_ifnext_pc_o_15))))

	.dataa(\IDEX|idex_if.imm_o [13]),
	.datab(\IDEX|idex_if.next_pc_o [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~25 ),
	.combout(\Add1~26_combout ),
	.cout(\Add1~27 ));
// synopsys translate_off
defparam \Add1~26 .lut_mask = 16'h9617;
defparam \Add1~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N0
cycloneive_lcell_comb \new_pc[15]~26 (
// Equation(s):
// \new_pc[15]~26_combout  = (\pc[31]~1_combout  & ((\pc[31]~2_combout  & ((idex_ifimm_26_o_13))) # (!\pc[31]~2_combout  & (idex_ifrdat1_o_15)))) # (!\pc[31]~1_combout  & (((\pc[31]~2_combout ))))

	.dataa(\pc[31]~1_combout ),
	.datab(\IDEX|idex_if.rdat1_o [15]),
	.datac(\IDEX|idex_if.imm_26_o [13]),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[15]~26_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[15]~26 .lut_mask = 16'hF588;
defparam \new_pc[15]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N2
cycloneive_lcell_comb \new_pc[15]~27 (
// Equation(s):
// \new_pc[15]~27_combout  = (\pc[31]~1_combout  & (((\new_pc[15]~26_combout )))) # (!\pc[31]~1_combout  & ((\new_pc[15]~26_combout  & ((\Add1~26_combout ))) # (!\new_pc[15]~26_combout  & (\nextpc[15]~26_combout ))))

	.dataa(\pc[31]~1_combout ),
	.datab(\nextpc[15]~26_combout ),
	.datac(\Add1~26_combout ),
	.datad(\new_pc[15]~26_combout ),
	.cin(gnd),
	.combout(\new_pc[15]~27_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[15]~27 .lut_mask = 16'hFA44;
defparam \new_pc[15]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N0
cycloneive_lcell_comb \new_pc[14]~28 (
// Equation(s):
// \new_pc[14]~28_combout  = (\pc[31]~1_combout  & ((idex_ifrdat1_o_14) # ((\pc[31]~2_combout )))) # (!\pc[31]~1_combout  & (((!\pc[31]~2_combout  & \nextpc[14]~24_combout ))))

	.dataa(\pc[31]~1_combout ),
	.datab(\IDEX|idex_if.rdat1_o [14]),
	.datac(\pc[31]~2_combout ),
	.datad(\nextpc[14]~24_combout ),
	.cin(gnd),
	.combout(\new_pc[14]~28_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[14]~28 .lut_mask = 16'hADA8;
defparam \new_pc[14]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N12
cycloneive_lcell_comb \new_pc[14]~29 (
// Equation(s):
// \new_pc[14]~29_combout  = (\pc[31]~2_combout  & ((\new_pc[14]~28_combout  & (idex_ifimm_26_o_12)) # (!\new_pc[14]~28_combout  & ((\Add1~24_combout ))))) # (!\pc[31]~2_combout  & (((\new_pc[14]~28_combout ))))

	.dataa(\IDEX|idex_if.imm_26_o [12]),
	.datab(\Add1~24_combout ),
	.datac(\pc[31]~2_combout ),
	.datad(\new_pc[14]~28_combout ),
	.cin(gnd),
	.combout(\new_pc[14]~29_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[14]~29 .lut_mask = 16'hAFC0;
defparam \new_pc[14]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N30
cycloneive_lcell_comb \Add1~28 (
// Equation(s):
// \Add1~28_combout  = ((idex_ifnext_pc_o_16 $ (idex_ifimm_o_14 $ (!\Add1~27 )))) # (GND)
// \Add1~29  = CARRY((idex_ifnext_pc_o_16 & ((idex_ifimm_o_14) # (!\Add1~27 ))) # (!idex_ifnext_pc_o_16 & (idex_ifimm_o_14 & !\Add1~27 )))

	.dataa(\IDEX|idex_if.next_pc_o [16]),
	.datab(\IDEX|idex_if.imm_o [14]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~27 ),
	.combout(\Add1~28_combout ),
	.cout(\Add1~29 ));
// synopsys translate_off
defparam \Add1~28 .lut_mask = 16'h698E;
defparam \Add1~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N0
cycloneive_lcell_comb \Add1~30 (
// Equation(s):
// \Add1~30_combout  = (idex_ifnext_pc_o_17 & ((idex_ifimm_o_15 & (\Add1~29  & VCC)) # (!idex_ifimm_o_15 & (!\Add1~29 )))) # (!idex_ifnext_pc_o_17 & ((idex_ifimm_o_15 & (!\Add1~29 )) # (!idex_ifimm_o_15 & ((\Add1~29 ) # (GND)))))
// \Add1~31  = CARRY((idex_ifnext_pc_o_17 & (!idex_ifimm_o_15 & !\Add1~29 )) # (!idex_ifnext_pc_o_17 & ((!\Add1~29 ) # (!idex_ifimm_o_15))))

	.dataa(\IDEX|idex_if.next_pc_o [17]),
	.datab(\IDEX|idex_if.imm_o [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~29 ),
	.combout(\Add1~30_combout ),
	.cout(\Add1~31 ));
// synopsys translate_off
defparam \Add1~30 .lut_mask = 16'h9617;
defparam \Add1~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N0
cycloneive_lcell_comb \nextpc[17]~30 (
// Equation(s):
// \nextpc[17]~30_combout  = (pc_17 & (!\nextpc[16]~29 )) # (!pc_17 & ((\nextpc[16]~29 ) # (GND)))
// \nextpc[17]~31  = CARRY((!\nextpc[16]~29 ) # (!pc_17))

	.dataa(gnd),
	.datab(pc_17),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[16]~29 ),
	.combout(\nextpc[17]~30_combout ),
	.cout(\nextpc[17]~31 ));
// synopsys translate_off
defparam \nextpc[17]~30 .lut_mask = 16'h3C3F;
defparam \nextpc[17]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N12
cycloneive_lcell_comb \new_pc[17]~30 (
// Equation(s):
// \new_pc[17]~30_combout  = (\pc[31]~1_combout  & ((\pc[31]~2_combout  & (idex_ifimm_26_o_15)) # (!\pc[31]~2_combout  & ((idex_ifrdat1_o_17))))) # (!\pc[31]~1_combout  & (((\pc[31]~2_combout ))))

	.dataa(\IDEX|idex_if.imm_26_o [15]),
	.datab(\pc[31]~1_combout ),
	.datac(\pc[31]~2_combout ),
	.datad(\IDEX|idex_if.rdat1_o [17]),
	.cin(gnd),
	.combout(\new_pc[17]~30_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[17]~30 .lut_mask = 16'hBCB0;
defparam \new_pc[17]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N4
cycloneive_lcell_comb \new_pc[17]~31 (
// Equation(s):
// \new_pc[17]~31_combout  = (\pc[31]~1_combout  & (((\new_pc[17]~30_combout )))) # (!\pc[31]~1_combout  & ((\new_pc[17]~30_combout  & (\Add1~30_combout )) # (!\new_pc[17]~30_combout  & ((\nextpc[17]~30_combout )))))

	.dataa(\Add1~30_combout ),
	.datab(\pc[31]~1_combout ),
	.datac(\nextpc[17]~30_combout ),
	.datad(\new_pc[17]~30_combout ),
	.cin(gnd),
	.combout(\new_pc[17]~31_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[17]~31 .lut_mask = 16'hEE30;
defparam \new_pc[17]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N14
cycloneive_lcell_comb \new_pc[16]~32 (
// Equation(s):
// \new_pc[16]~32_combout  = (\pc[31]~2_combout  & (((\pc[31]~1_combout )))) # (!\pc[31]~2_combout  & ((\pc[31]~1_combout  & ((idex_ifrdat1_o_16))) # (!\pc[31]~1_combout  & (\nextpc[16]~28_combout ))))

	.dataa(\nextpc[16]~28_combout ),
	.datab(\IDEX|idex_if.rdat1_o [16]),
	.datac(\pc[31]~2_combout ),
	.datad(\pc[31]~1_combout ),
	.cin(gnd),
	.combout(\new_pc[16]~32_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[16]~32 .lut_mask = 16'hFC0A;
defparam \new_pc[16]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N8
cycloneive_lcell_comb \new_pc[16]~33 (
// Equation(s):
// \new_pc[16]~33_combout  = (\pc[31]~2_combout  & ((\new_pc[16]~32_combout  & ((idex_ifimm_26_o_14))) # (!\new_pc[16]~32_combout  & (\Add1~28_combout )))) # (!\pc[31]~2_combout  & (((\new_pc[16]~32_combout ))))

	.dataa(\Add1~28_combout ),
	.datab(\IDEX|idex_if.imm_26_o [14]),
	.datac(\pc[31]~2_combout ),
	.datad(\new_pc[16]~32_combout ),
	.cin(gnd),
	.combout(\new_pc[16]~33_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[16]~33 .lut_mask = 16'hCFA0;
defparam \new_pc[16]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N2
cycloneive_lcell_comb \Add1~32 (
// Equation(s):
// \Add1~32_combout  = ((idex_ifnext_pc_o_18 $ (idex_ifimm_o_15 $ (!\Add1~31 )))) # (GND)
// \Add1~33  = CARRY((idex_ifnext_pc_o_18 & ((idex_ifimm_o_15) # (!\Add1~31 ))) # (!idex_ifnext_pc_o_18 & (idex_ifimm_o_15 & !\Add1~31 )))

	.dataa(\IDEX|idex_if.next_pc_o [18]),
	.datab(\IDEX|idex_if.imm_o [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~31 ),
	.combout(\Add1~32_combout ),
	.cout(\Add1~33 ));
// synopsys translate_off
defparam \Add1~32 .lut_mask = 16'h698E;
defparam \Add1~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N4
cycloneive_lcell_comb \Add1~34 (
// Equation(s):
// \Add1~34_combout  = (idex_ifnext_pc_o_19 & ((idex_ifimm_o_15 & (\Add1~33  & VCC)) # (!idex_ifimm_o_15 & (!\Add1~33 )))) # (!idex_ifnext_pc_o_19 & ((idex_ifimm_o_15 & (!\Add1~33 )) # (!idex_ifimm_o_15 & ((\Add1~33 ) # (GND)))))
// \Add1~35  = CARRY((idex_ifnext_pc_o_19 & (!idex_ifimm_o_15 & !\Add1~33 )) # (!idex_ifnext_pc_o_19 & ((!\Add1~33 ) # (!idex_ifimm_o_15))))

	.dataa(\IDEX|idex_if.next_pc_o [19]),
	.datab(\IDEX|idex_if.imm_o [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~33 ),
	.combout(\Add1~34_combout ),
	.cout(\Add1~35 ));
// synopsys translate_off
defparam \Add1~34 .lut_mask = 16'h9617;
defparam \Add1~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N4
cycloneive_lcell_comb \nextpc[19]~34 (
// Equation(s):
// \nextpc[19]~34_combout  = (pc_19 & (!\nextpc[18]~33 )) # (!pc_19 & ((\nextpc[18]~33 ) # (GND)))
// \nextpc[19]~35  = CARRY((!\nextpc[18]~33 ) # (!pc_19))

	.dataa(pc_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[18]~33 ),
	.combout(\nextpc[19]~34_combout ),
	.cout(\nextpc[19]~35 ));
// synopsys translate_off
defparam \nextpc[19]~34 .lut_mask = 16'h5A5F;
defparam \nextpc[19]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N6
cycloneive_lcell_comb \new_pc[19]~34 (
// Equation(s):
// \new_pc[19]~34_combout  = (\pc[31]~1_combout  & ((\pc[31]~2_combout  & (idex_ifimm_26_o_17)) # (!\pc[31]~2_combout  & ((idex_ifrdat1_o_19))))) # (!\pc[31]~1_combout  & (((\pc[31]~2_combout ))))

	.dataa(\IDEX|idex_if.imm_26_o [17]),
	.datab(\pc[31]~1_combout ),
	.datac(\IDEX|idex_if.rdat1_o [19]),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[19]~34_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[19]~34 .lut_mask = 16'hBBC0;
defparam \new_pc[19]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N14
cycloneive_lcell_comb \new_pc[19]~35 (
// Equation(s):
// \new_pc[19]~35_combout  = (\pc[31]~1_combout  & (((\new_pc[19]~34_combout )))) # (!\pc[31]~1_combout  & ((\new_pc[19]~34_combout  & (\Add1~34_combout )) # (!\new_pc[19]~34_combout  & ((\nextpc[19]~34_combout )))))

	.dataa(\Add1~34_combout ),
	.datab(\pc[31]~1_combout ),
	.datac(\nextpc[19]~34_combout ),
	.datad(\new_pc[19]~34_combout ),
	.cin(gnd),
	.combout(\new_pc[19]~35_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[19]~35 .lut_mask = 16'hEE30;
defparam \new_pc[19]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N26
cycloneive_lcell_comb \new_pc[18]~36 (
// Equation(s):
// \new_pc[18]~36_combout  = (\pc[31]~1_combout  & (((idex_ifrdat1_o_18) # (\pc[31]~2_combout )))) # (!\pc[31]~1_combout  & (\nextpc[18]~32_combout  & ((!\pc[31]~2_combout ))))

	.dataa(\nextpc[18]~32_combout ),
	.datab(\pc[31]~1_combout ),
	.datac(\IDEX|idex_if.rdat1_o [18]),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[18]~36_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[18]~36 .lut_mask = 16'hCCE2;
defparam \new_pc[18]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N4
cycloneive_lcell_comb \new_pc[18]~37 (
// Equation(s):
// \new_pc[18]~37_combout  = (\new_pc[18]~36_combout  & ((idex_ifimm_26_o_16) # ((!\pc[31]~2_combout )))) # (!\new_pc[18]~36_combout  & (((\Add1~32_combout  & \pc[31]~2_combout ))))

	.dataa(\IDEX|idex_if.imm_26_o [16]),
	.datab(\Add1~32_combout ),
	.datac(\new_pc[18]~36_combout ),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[18]~37_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[18]~37 .lut_mask = 16'hACF0;
defparam \new_pc[18]~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N6
cycloneive_lcell_comb \Add1~36 (
// Equation(s):
// \Add1~36_combout  = ((idex_ifnext_pc_o_20 $ (idex_ifimm_o_15 $ (!\Add1~35 )))) # (GND)
// \Add1~37  = CARRY((idex_ifnext_pc_o_20 & ((idex_ifimm_o_15) # (!\Add1~35 ))) # (!idex_ifnext_pc_o_20 & (idex_ifimm_o_15 & !\Add1~35 )))

	.dataa(\IDEX|idex_if.next_pc_o [20]),
	.datab(\IDEX|idex_if.imm_o [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~35 ),
	.combout(\Add1~36_combout ),
	.cout(\Add1~37 ));
// synopsys translate_off
defparam \Add1~36 .lut_mask = 16'h698E;
defparam \Add1~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N8
cycloneive_lcell_comb \Add1~38 (
// Equation(s):
// \Add1~38_combout  = (idex_ifnext_pc_o_21 & ((idex_ifimm_o_15 & (\Add1~37  & VCC)) # (!idex_ifimm_o_15 & (!\Add1~37 )))) # (!idex_ifnext_pc_o_21 & ((idex_ifimm_o_15 & (!\Add1~37 )) # (!idex_ifimm_o_15 & ((\Add1~37 ) # (GND)))))
// \Add1~39  = CARRY((idex_ifnext_pc_o_21 & (!idex_ifimm_o_15 & !\Add1~37 )) # (!idex_ifnext_pc_o_21 & ((!\Add1~37 ) # (!idex_ifimm_o_15))))

	.dataa(\IDEX|idex_if.next_pc_o [21]),
	.datab(\IDEX|idex_if.imm_o [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~37 ),
	.combout(\Add1~38_combout ),
	.cout(\Add1~39 ));
// synopsys translate_off
defparam \Add1~38 .lut_mask = 16'h9617;
defparam \Add1~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N6
cycloneive_lcell_comb \nextpc[20]~36 (
// Equation(s):
// \nextpc[20]~36_combout  = (pc_20 & (\nextpc[19]~35  $ (GND))) # (!pc_20 & (!\nextpc[19]~35  & VCC))
// \nextpc[20]~37  = CARRY((pc_20 & !\nextpc[19]~35 ))

	.dataa(pc_20),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[19]~35 ),
	.combout(\nextpc[20]~36_combout ),
	.cout(\nextpc[20]~37 ));
// synopsys translate_off
defparam \nextpc[20]~36 .lut_mask = 16'hA50A;
defparam \nextpc[20]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N8
cycloneive_lcell_comb \nextpc[21]~38 (
// Equation(s):
// \nextpc[21]~38_combout  = (pc_21 & (!\nextpc[20]~37 )) # (!pc_21 & ((\nextpc[20]~37 ) # (GND)))
// \nextpc[21]~39  = CARRY((!\nextpc[20]~37 ) # (!pc_21))

	.dataa(pc_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[20]~37 ),
	.combout(\nextpc[21]~38_combout ),
	.cout(\nextpc[21]~39 ));
// synopsys translate_off
defparam \nextpc[21]~38 .lut_mask = 16'h5A5F;
defparam \nextpc[21]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N6
cycloneive_lcell_comb \new_pc[21]~38 (
// Equation(s):
// \new_pc[21]~38_combout  = (\pc[31]~1_combout  & ((\pc[31]~2_combout  & (idex_ifimm_26_o_19)) # (!\pc[31]~2_combout  & ((idex_ifrdat1_o_21))))) # (!\pc[31]~1_combout  & (((\pc[31]~2_combout ))))

	.dataa(\IDEX|idex_if.imm_26_o [19]),
	.datab(\IDEX|idex_if.rdat1_o [21]),
	.datac(\pc[31]~1_combout ),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[21]~38_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[21]~38 .lut_mask = 16'hAFC0;
defparam \new_pc[21]~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N4
cycloneive_lcell_comb \new_pc[21]~39 (
// Equation(s):
// \new_pc[21]~39_combout  = (\pc[31]~1_combout  & (((\new_pc[21]~38_combout )))) # (!\pc[31]~1_combout  & ((\new_pc[21]~38_combout  & (\Add1~38_combout )) # (!\new_pc[21]~38_combout  & ((\nextpc[21]~38_combout )))))

	.dataa(\Add1~38_combout ),
	.datab(\nextpc[21]~38_combout ),
	.datac(\pc[31]~1_combout ),
	.datad(\new_pc[21]~38_combout ),
	.cin(gnd),
	.combout(\new_pc[21]~39_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[21]~39 .lut_mask = 16'hFA0C;
defparam \new_pc[21]~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N14
cycloneive_lcell_comb \new_pc[20]~40 (
// Equation(s):
// \new_pc[20]~40_combout  = (\pc[31]~1_combout  & ((idex_ifrdat1_o_20) # ((\pc[31]~2_combout )))) # (!\pc[31]~1_combout  & (((\nextpc[20]~36_combout  & !\pc[31]~2_combout ))))

	.dataa(\IDEX|idex_if.rdat1_o [20]),
	.datab(\pc[31]~1_combout ),
	.datac(\nextpc[20]~36_combout ),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[20]~40_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[20]~40 .lut_mask = 16'hCCB8;
defparam \new_pc[20]~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N0
cycloneive_lcell_comb \new_pc[20]~41 (
// Equation(s):
// \new_pc[20]~41_combout  = (\new_pc[20]~40_combout  & (((idex_ifimm_26_o_18) # (!\pc[31]~2_combout )))) # (!\new_pc[20]~40_combout  & (\Add1~36_combout  & ((\pc[31]~2_combout ))))

	.dataa(\Add1~36_combout ),
	.datab(\IDEX|idex_if.imm_26_o [18]),
	.datac(\new_pc[20]~40_combout ),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[20]~41_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[20]~41 .lut_mask = 16'hCAF0;
defparam \new_pc[20]~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N10
cycloneive_lcell_comb \Add1~40 (
// Equation(s):
// \Add1~40_combout  = ((idex_ifnext_pc_o_22 $ (idex_ifimm_o_15 $ (!\Add1~39 )))) # (GND)
// \Add1~41  = CARRY((idex_ifnext_pc_o_22 & ((idex_ifimm_o_15) # (!\Add1~39 ))) # (!idex_ifnext_pc_o_22 & (idex_ifimm_o_15 & !\Add1~39 )))

	.dataa(\IDEX|idex_if.next_pc_o [22]),
	.datab(\IDEX|idex_if.imm_o [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~39 ),
	.combout(\Add1~40_combout ),
	.cout(\Add1~41 ));
// synopsys translate_off
defparam \Add1~40 .lut_mask = 16'h698E;
defparam \Add1~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N12
cycloneive_lcell_comb \Add1~42 (
// Equation(s):
// \Add1~42_combout  = (idex_ifimm_o_15 & ((idex_ifnext_pc_o_23 & (\Add1~41  & VCC)) # (!idex_ifnext_pc_o_23 & (!\Add1~41 )))) # (!idex_ifimm_o_15 & ((idex_ifnext_pc_o_23 & (!\Add1~41 )) # (!idex_ifnext_pc_o_23 & ((\Add1~41 ) # (GND)))))
// \Add1~43  = CARRY((idex_ifimm_o_15 & (!idex_ifnext_pc_o_23 & !\Add1~41 )) # (!idex_ifimm_o_15 & ((!\Add1~41 ) # (!idex_ifnext_pc_o_23))))

	.dataa(\IDEX|idex_if.imm_o [15]),
	.datab(\IDEX|idex_if.next_pc_o [23]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~41 ),
	.combout(\Add1~42_combout ),
	.cout(\Add1~43 ));
// synopsys translate_off
defparam \Add1~42 .lut_mask = 16'h9617;
defparam \Add1~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N10
cycloneive_lcell_comb \nextpc[22]~40 (
// Equation(s):
// \nextpc[22]~40_combout  = (pc_22 & (\nextpc[21]~39  $ (GND))) # (!pc_22 & (!\nextpc[21]~39  & VCC))
// \nextpc[22]~41  = CARRY((pc_22 & !\nextpc[21]~39 ))

	.dataa(pc_22),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[21]~39 ),
	.combout(\nextpc[22]~40_combout ),
	.cout(\nextpc[22]~41 ));
// synopsys translate_off
defparam \nextpc[22]~40 .lut_mask = 16'hA50A;
defparam \nextpc[22]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N12
cycloneive_lcell_comb \nextpc[23]~42 (
// Equation(s):
// \nextpc[23]~42_combout  = (pc_23 & (!\nextpc[22]~41 )) # (!pc_23 & ((\nextpc[22]~41 ) # (GND)))
// \nextpc[23]~43  = CARRY((!\nextpc[22]~41 ) # (!pc_23))

	.dataa(gnd),
	.datab(pc_23),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[22]~41 ),
	.combout(\nextpc[23]~42_combout ),
	.cout(\nextpc[23]~43 ));
// synopsys translate_off
defparam \nextpc[23]~42 .lut_mask = 16'h3C3F;
defparam \nextpc[23]~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N28
cycloneive_lcell_comb \new_pc[23]~42 (
// Equation(s):
// \new_pc[23]~42_combout  = (\pc[31]~1_combout  & ((\pc[31]~2_combout  & ((idex_ifimm_26_o_21))) # (!\pc[31]~2_combout  & (idex_ifrdat1_o_23)))) # (!\pc[31]~1_combout  & (((\pc[31]~2_combout ))))

	.dataa(\IDEX|idex_if.rdat1_o [23]),
	.datab(\pc[31]~1_combout ),
	.datac(\IDEX|idex_if.imm_26_o [21]),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[23]~42_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[23]~42 .lut_mask = 16'hF388;
defparam \new_pc[23]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N22
cycloneive_lcell_comb \new_pc[23]~43 (
// Equation(s):
// \new_pc[23]~43_combout  = (\pc[31]~1_combout  & (((\new_pc[23]~42_combout )))) # (!\pc[31]~1_combout  & ((\new_pc[23]~42_combout  & (\Add1~42_combout )) # (!\new_pc[23]~42_combout  & ((\nextpc[23]~42_combout )))))

	.dataa(\Add1~42_combout ),
	.datab(\pc[31]~1_combout ),
	.datac(\nextpc[23]~42_combout ),
	.datad(\new_pc[23]~42_combout ),
	.cin(gnd),
	.combout(\new_pc[23]~43_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[23]~43 .lut_mask = 16'hEE30;
defparam \new_pc[23]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N0
cycloneive_lcell_comb \new_pc[22]~44 (
// Equation(s):
// \new_pc[22]~44_combout  = (\pc[31]~1_combout  & ((idex_ifrdat1_o_22) # ((\pc[31]~2_combout )))) # (!\pc[31]~1_combout  & (((\nextpc[22]~40_combout  & !\pc[31]~2_combout ))))

	.dataa(\IDEX|idex_if.rdat1_o [22]),
	.datab(\pc[31]~1_combout ),
	.datac(\nextpc[22]~40_combout ),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[22]~44_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[22]~44 .lut_mask = 16'hCCB8;
defparam \new_pc[22]~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N28
cycloneive_lcell_comb \new_pc[22]~45 (
// Equation(s):
// \new_pc[22]~45_combout  = (\pc[31]~2_combout  & ((\new_pc[22]~44_combout  & ((idex_ifimm_26_o_20))) # (!\new_pc[22]~44_combout  & (\Add1~40_combout )))) # (!\pc[31]~2_combout  & (((\new_pc[22]~44_combout ))))

	.dataa(\Add1~40_combout ),
	.datab(\IDEX|idex_if.imm_26_o [20]),
	.datac(\pc[31]~2_combout ),
	.datad(\new_pc[22]~44_combout ),
	.cin(gnd),
	.combout(\new_pc[22]~45_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[22]~45 .lut_mask = 16'hCFA0;
defparam \new_pc[22]~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N16
cycloneive_lcell_comb \nextpc[25]~46 (
// Equation(s):
// \nextpc[25]~46_combout  = (pc_25 & (!\nextpc[24]~45 )) # (!pc_25 & ((\nextpc[24]~45 ) # (GND)))
// \nextpc[25]~47  = CARRY((!\nextpc[24]~45 ) # (!pc_25))

	.dataa(pc_25),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[24]~45 ),
	.combout(\nextpc[25]~46_combout ),
	.cout(\nextpc[25]~47 ));
// synopsys translate_off
defparam \nextpc[25]~46 .lut_mask = 16'h5A5F;
defparam \nextpc[25]~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N14
cycloneive_lcell_comb \Add1~44 (
// Equation(s):
// \Add1~44_combout  = ((idex_ifimm_o_15 $ (idex_ifnext_pc_o_24 $ (!\Add1~43 )))) # (GND)
// \Add1~45  = CARRY((idex_ifimm_o_15 & ((idex_ifnext_pc_o_24) # (!\Add1~43 ))) # (!idex_ifimm_o_15 & (idex_ifnext_pc_o_24 & !\Add1~43 )))

	.dataa(\IDEX|idex_if.imm_o [15]),
	.datab(\IDEX|idex_if.next_pc_o [24]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~43 ),
	.combout(\Add1~44_combout ),
	.cout(\Add1~45 ));
// synopsys translate_off
defparam \Add1~44 .lut_mask = 16'h698E;
defparam \Add1~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N16
cycloneive_lcell_comb \Add1~46 (
// Equation(s):
// \Add1~46_combout  = (idex_ifimm_o_15 & ((idex_ifnext_pc_o_25 & (\Add1~45  & VCC)) # (!idex_ifnext_pc_o_25 & (!\Add1~45 )))) # (!idex_ifimm_o_15 & ((idex_ifnext_pc_o_25 & (!\Add1~45 )) # (!idex_ifnext_pc_o_25 & ((\Add1~45 ) # (GND)))))
// \Add1~47  = CARRY((idex_ifimm_o_15 & (!idex_ifnext_pc_o_25 & !\Add1~45 )) # (!idex_ifimm_o_15 & ((!\Add1~45 ) # (!idex_ifnext_pc_o_25))))

	.dataa(\IDEX|idex_if.imm_o [15]),
	.datab(\IDEX|idex_if.next_pc_o [25]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~45 ),
	.combout(\Add1~46_combout ),
	.cout(\Add1~47 ));
// synopsys translate_off
defparam \Add1~46 .lut_mask = 16'h9617;
defparam \Add1~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N10
cycloneive_lcell_comb \new_pc[25]~46 (
// Equation(s):
// \new_pc[25]~46_combout  = (\pc[31]~1_combout  & ((\pc[31]~2_combout  & ((idex_ifimm_26_o_23))) # (!\pc[31]~2_combout  & (idex_ifrdat1_o_25)))) # (!\pc[31]~1_combout  & (((\pc[31]~2_combout ))))

	.dataa(\pc[31]~1_combout ),
	.datab(\IDEX|idex_if.rdat1_o [25]),
	.datac(\IDEX|idex_if.imm_26_o [23]),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[25]~46_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[25]~46 .lut_mask = 16'hF588;
defparam \new_pc[25]~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N24
cycloneive_lcell_comb \new_pc[25]~47 (
// Equation(s):
// \new_pc[25]~47_combout  = (\pc[31]~1_combout  & (((\new_pc[25]~46_combout )))) # (!\pc[31]~1_combout  & ((\new_pc[25]~46_combout  & ((\Add1~46_combout ))) # (!\new_pc[25]~46_combout  & (\nextpc[25]~46_combout ))))

	.dataa(\pc[31]~1_combout ),
	.datab(\nextpc[25]~46_combout ),
	.datac(\Add1~46_combout ),
	.datad(\new_pc[25]~46_combout ),
	.cin(gnd),
	.combout(\new_pc[25]~47_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[25]~47 .lut_mask = 16'hFA44;
defparam \new_pc[25]~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N22
cycloneive_lcell_comb \new_pc[24]~48 (
// Equation(s):
// \new_pc[24]~48_combout  = (\pc[31]~1_combout  & (((idex_ifrdat1_o_24) # (\pc[31]~2_combout )))) # (!\pc[31]~1_combout  & (\nextpc[24]~44_combout  & ((!\pc[31]~2_combout ))))

	.dataa(\nextpc[24]~44_combout ),
	.datab(\IDEX|idex_if.rdat1_o [24]),
	.datac(\pc[31]~1_combout ),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[24]~48_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[24]~48 .lut_mask = 16'hF0CA;
defparam \new_pc[24]~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N26
cycloneive_lcell_comb \new_pc[24]~49 (
// Equation(s):
// \new_pc[24]~49_combout  = (\new_pc[24]~48_combout  & (((idex_ifimm_26_o_22) # (!\pc[31]~2_combout )))) # (!\new_pc[24]~48_combout  & (\Add1~44_combout  & ((\pc[31]~2_combout ))))

	.dataa(\Add1~44_combout ),
	.datab(\IDEX|idex_if.imm_26_o [22]),
	.datac(\new_pc[24]~48_combout ),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[24]~49_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[24]~49 .lut_mask = 16'hCAF0;
defparam \new_pc[24]~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N20
cycloneive_lcell_comb \nextpc[27]~50 (
// Equation(s):
// \nextpc[27]~50_combout  = (pc_27 & (!\nextpc[26]~49 )) # (!pc_27 & ((\nextpc[26]~49 ) # (GND)))
// \nextpc[27]~51  = CARRY((!\nextpc[26]~49 ) # (!pc_27))

	.dataa(gnd),
	.datab(pc_27),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[26]~49 ),
	.combout(\nextpc[27]~50_combout ),
	.cout(\nextpc[27]~51 ));
// synopsys translate_off
defparam \nextpc[27]~50 .lut_mask = 16'h3C3F;
defparam \nextpc[27]~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N18
cycloneive_lcell_comb \Add1~48 (
// Equation(s):
// \Add1~48_combout  = ((idex_ifimm_o_15 $ (idex_ifnext_pc_o_26 $ (!\Add1~47 )))) # (GND)
// \Add1~49  = CARRY((idex_ifimm_o_15 & ((idex_ifnext_pc_o_26) # (!\Add1~47 ))) # (!idex_ifimm_o_15 & (idex_ifnext_pc_o_26 & !\Add1~47 )))

	.dataa(\IDEX|idex_if.imm_o [15]),
	.datab(\IDEX|idex_if.next_pc_o [26]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~47 ),
	.combout(\Add1~48_combout ),
	.cout(\Add1~49 ));
// synopsys translate_off
defparam \Add1~48 .lut_mask = 16'h698E;
defparam \Add1~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N20
cycloneive_lcell_comb \Add1~50 (
// Equation(s):
// \Add1~50_combout  = (idex_ifimm_o_15 & ((idex_ifnext_pc_o_27 & (\Add1~49  & VCC)) # (!idex_ifnext_pc_o_27 & (!\Add1~49 )))) # (!idex_ifimm_o_15 & ((idex_ifnext_pc_o_27 & (!\Add1~49 )) # (!idex_ifnext_pc_o_27 & ((\Add1~49 ) # (GND)))))
// \Add1~51  = CARRY((idex_ifimm_o_15 & (!idex_ifnext_pc_o_27 & !\Add1~49 )) # (!idex_ifimm_o_15 & ((!\Add1~49 ) # (!idex_ifnext_pc_o_27))))

	.dataa(\IDEX|idex_if.imm_o [15]),
	.datab(\IDEX|idex_if.next_pc_o [27]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~49 ),
	.combout(\Add1~50_combout ),
	.cout(\Add1~51 ));
// synopsys translate_off
defparam \Add1~50 .lut_mask = 16'h9617;
defparam \Add1~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N16
cycloneive_lcell_comb \new_pc[27]~50 (
// Equation(s):
// \new_pc[27]~50_combout  = (\pc[31]~1_combout  & ((\pc[31]~2_combout  & (idex_ifimm_26_o_25)) # (!\pc[31]~2_combout  & ((idex_ifrdat1_o_27))))) # (!\pc[31]~1_combout  & (((\pc[31]~2_combout ))))

	.dataa(\pc[31]~1_combout ),
	.datab(\IDEX|idex_if.imm_26_o [25]),
	.datac(\IDEX|idex_if.rdat1_o [27]),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[27]~50_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[27]~50 .lut_mask = 16'hDDA0;
defparam \new_pc[27]~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N12
cycloneive_lcell_comb \new_pc[27]~51 (
// Equation(s):
// \new_pc[27]~51_combout  = (\pc[31]~1_combout  & (((\new_pc[27]~50_combout )))) # (!\pc[31]~1_combout  & ((\new_pc[27]~50_combout  & ((\Add1~50_combout ))) # (!\new_pc[27]~50_combout  & (\nextpc[27]~50_combout ))))

	.dataa(\pc[31]~1_combout ),
	.datab(\nextpc[27]~50_combout ),
	.datac(\Add1~50_combout ),
	.datad(\new_pc[27]~50_combout ),
	.cin(gnd),
	.combout(\new_pc[27]~51_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[27]~51 .lut_mask = 16'hFA44;
defparam \new_pc[27]~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N14
cycloneive_lcell_comb \new_pc[26]~52 (
// Equation(s):
// \new_pc[26]~52_combout  = (\pc[31]~1_combout  & (((idex_ifrdat1_o_26) # (\pc[31]~2_combout )))) # (!\pc[31]~1_combout  & (\nextpc[26]~48_combout  & ((!\pc[31]~2_combout ))))

	.dataa(\nextpc[26]~48_combout ),
	.datab(\IDEX|idex_if.rdat1_o [26]),
	.datac(\pc[31]~1_combout ),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[26]~52_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[26]~52 .lut_mask = 16'hF0CA;
defparam \new_pc[26]~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N8
cycloneive_lcell_comb \new_pc[26]~53 (
// Equation(s):
// \new_pc[26]~53_combout  = (\new_pc[26]~52_combout  & ((idex_ifimm_26_o_24) # ((!\pc[31]~2_combout )))) # (!\new_pc[26]~52_combout  & (((\Add1~48_combout  & \pc[31]~2_combout ))))

	.dataa(\IDEX|idex_if.imm_26_o [24]),
	.datab(\Add1~48_combout ),
	.datac(\new_pc[26]~52_combout ),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[26]~53_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[26]~53 .lut_mask = 16'hACF0;
defparam \new_pc[26]~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N22
cycloneive_lcell_comb \Add1~52 (
// Equation(s):
// \Add1~52_combout  = ((idex_ifimm_o_15 $ (idex_ifnext_pc_o_28 $ (!\Add1~51 )))) # (GND)
// \Add1~53  = CARRY((idex_ifimm_o_15 & ((idex_ifnext_pc_o_28) # (!\Add1~51 ))) # (!idex_ifimm_o_15 & (idex_ifnext_pc_o_28 & !\Add1~51 )))

	.dataa(\IDEX|idex_if.imm_o [15]),
	.datab(\IDEX|idex_if.next_pc_o [28]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~51 ),
	.combout(\Add1~52_combout ),
	.cout(\Add1~53 ));
// synopsys translate_off
defparam \Add1~52 .lut_mask = 16'h698E;
defparam \Add1~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N24
cycloneive_lcell_comb \Add1~54 (
// Equation(s):
// \Add1~54_combout  = (idex_ifimm_o_15 & ((idex_ifnext_pc_o_29 & (\Add1~53  & VCC)) # (!idex_ifnext_pc_o_29 & (!\Add1~53 )))) # (!idex_ifimm_o_15 & ((idex_ifnext_pc_o_29 & (!\Add1~53 )) # (!idex_ifnext_pc_o_29 & ((\Add1~53 ) # (GND)))))
// \Add1~55  = CARRY((idex_ifimm_o_15 & (!idex_ifnext_pc_o_29 & !\Add1~53 )) # (!idex_ifimm_o_15 & ((!\Add1~53 ) # (!idex_ifnext_pc_o_29))))

	.dataa(\IDEX|idex_if.imm_o [15]),
	.datab(\IDEX|idex_if.next_pc_o [29]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~53 ),
	.combout(\Add1~54_combout ),
	.cout(\Add1~55 ));
// synopsys translate_off
defparam \Add1~54 .lut_mask = 16'h9617;
defparam \Add1~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N24
cycloneive_lcell_comb \nextpc[29]~54 (
// Equation(s):
// \nextpc[29]~54_combout  = (pc_29 & (!\nextpc[28]~53 )) # (!pc_29 & ((\nextpc[28]~53 ) # (GND)))
// \nextpc[29]~55  = CARRY((!\nextpc[28]~53 ) # (!pc_29))

	.dataa(gnd),
	.datab(pc_29),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[28]~53 ),
	.combout(\nextpc[29]~54_combout ),
	.cout(\nextpc[29]~55 ));
// synopsys translate_off
defparam \nextpc[29]~54 .lut_mask = 16'h3C3F;
defparam \nextpc[29]~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N16
cycloneive_lcell_comb \new_pc[29]~54 (
// Equation(s):
// \new_pc[29]~54_combout  = (\pc[31]~1_combout  & ((\pc[31]~2_combout  & (idex_ifnext_pc_o_29)) # (!\pc[31]~2_combout  & ((idex_ifrdat1_o_29))))) # (!\pc[31]~1_combout  & (((\pc[31]~2_combout ))))

	.dataa(\pc[31]~1_combout ),
	.datab(\IDEX|idex_if.next_pc_o [29]),
	.datac(\IDEX|idex_if.rdat1_o [29]),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[29]~54_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[29]~54 .lut_mask = 16'hDDA0;
defparam \new_pc[29]~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N4
cycloneive_lcell_comb \new_pc[29]~55 (
// Equation(s):
// \new_pc[29]~55_combout  = (\pc[31]~1_combout  & (((\new_pc[29]~54_combout )))) # (!\pc[31]~1_combout  & ((\new_pc[29]~54_combout  & (\Add1~54_combout )) # (!\new_pc[29]~54_combout  & ((\nextpc[29]~54_combout )))))

	.dataa(\pc[31]~1_combout ),
	.datab(\Add1~54_combout ),
	.datac(\nextpc[29]~54_combout ),
	.datad(\new_pc[29]~54_combout ),
	.cin(gnd),
	.combout(\new_pc[29]~55_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[29]~55 .lut_mask = 16'hEE50;
defparam \new_pc[29]~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N12
cycloneive_lcell_comb \new_pc[28]~56 (
// Equation(s):
// \new_pc[28]~56_combout  = (\pc[31]~1_combout  & (((idex_ifrdat1_o_28) # (\pc[31]~2_combout )))) # (!\pc[31]~1_combout  & (\nextpc[28]~52_combout  & ((!\pc[31]~2_combout ))))

	.dataa(\nextpc[28]~52_combout ),
	.datab(\IDEX|idex_if.rdat1_o [28]),
	.datac(\pc[31]~1_combout ),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[28]~56_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[28]~56 .lut_mask = 16'hF0CA;
defparam \new_pc[28]~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N28
cycloneive_lcell_comb \new_pc[28]~57 (
// Equation(s):
// \new_pc[28]~57_combout  = (\pc[31]~2_combout  & ((\new_pc[28]~56_combout  & (idex_ifnext_pc_o_28)) # (!\new_pc[28]~56_combout  & ((\Add1~52_combout ))))) # (!\pc[31]~2_combout  & (((\new_pc[28]~56_combout ))))

	.dataa(\pc[31]~2_combout ),
	.datab(\IDEX|idex_if.next_pc_o [28]),
	.datac(\Add1~52_combout ),
	.datad(\new_pc[28]~56_combout ),
	.cin(gnd),
	.combout(\new_pc[28]~57_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[28]~57 .lut_mask = 16'hDDA0;
defparam \new_pc[28]~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N26
cycloneive_lcell_comb \nextpc[30]~56 (
// Equation(s):
// \nextpc[30]~56_combout  = (pc_30 & (\nextpc[29]~55  $ (GND))) # (!pc_30 & (!\nextpc[29]~55  & VCC))
// \nextpc[30]~57  = CARRY((pc_30 & !\nextpc[29]~55 ))

	.dataa(pc_30),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nextpc[29]~55 ),
	.combout(\nextpc[30]~56_combout ),
	.cout(\nextpc[30]~57 ));
// synopsys translate_off
defparam \nextpc[30]~56 .lut_mask = 16'hA50A;
defparam \nextpc[30]~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N28
cycloneive_lcell_comb \nextpc[31]~58 (
// Equation(s):
// \nextpc[31]~58_combout  = \nextpc[30]~57  $ (pc_31)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(pc_31),
	.cin(\nextpc[30]~57 ),
	.combout(\nextpc[31]~58_combout ),
	.cout());
// synopsys translate_off
defparam \nextpc[31]~58 .lut_mask = 16'h0FF0;
defparam \nextpc[31]~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N26
cycloneive_lcell_comb \Add1~56 (
// Equation(s):
// \Add1~56_combout  = ((idex_ifnext_pc_o_30 $ (idex_ifimm_o_15 $ (!\Add1~55 )))) # (GND)
// \Add1~57  = CARRY((idex_ifnext_pc_o_30 & ((idex_ifimm_o_15) # (!\Add1~55 ))) # (!idex_ifnext_pc_o_30 & (idex_ifimm_o_15 & !\Add1~55 )))

	.dataa(\IDEX|idex_if.next_pc_o [30]),
	.datab(\IDEX|idex_if.imm_o [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~55 ),
	.combout(\Add1~56_combout ),
	.cout(\Add1~57 ));
// synopsys translate_off
defparam \Add1~56 .lut_mask = 16'h698E;
defparam \Add1~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N28
cycloneive_lcell_comb \Add1~58 (
// Equation(s):
// \Add1~58_combout  = idex_ifnext_pc_o_31 $ (\Add1~57  $ (idex_ifimm_o_15))

	.dataa(gnd),
	.datab(\IDEX|idex_if.next_pc_o [31]),
	.datac(gnd),
	.datad(\IDEX|idex_if.imm_o [15]),
	.cin(\Add1~57 ),
	.combout(\Add1~58_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~58 .lut_mask = 16'hC33C;
defparam \Add1~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N10
cycloneive_lcell_comb \new_pc[31]~58 (
// Equation(s):
// \new_pc[31]~58_combout  = (\pc[31]~1_combout  & ((\pc[31]~2_combout  & ((idex_ifnext_pc_o_31))) # (!\pc[31]~2_combout  & (idex_ifrdat1_o_31)))) # (!\pc[31]~1_combout  & (((\pc[31]~2_combout ))))

	.dataa(\pc[31]~1_combout ),
	.datab(\IDEX|idex_if.rdat1_o [31]),
	.datac(\pc[31]~2_combout ),
	.datad(\IDEX|idex_if.next_pc_o [31]),
	.cin(gnd),
	.combout(\new_pc[31]~58_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[31]~58 .lut_mask = 16'hF858;
defparam \new_pc[31]~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N18
cycloneive_lcell_comb \new_pc[31]~59 (
// Equation(s):
// \new_pc[31]~59_combout  = (\pc[31]~1_combout  & (((\new_pc[31]~58_combout )))) # (!\pc[31]~1_combout  & ((\new_pc[31]~58_combout  & ((\Add1~58_combout ))) # (!\new_pc[31]~58_combout  & (\nextpc[31]~58_combout ))))

	.dataa(\pc[31]~1_combout ),
	.datab(\nextpc[31]~58_combout ),
	.datac(\Add1~58_combout ),
	.datad(\new_pc[31]~58_combout ),
	.cin(gnd),
	.combout(\new_pc[31]~59_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[31]~59 .lut_mask = 16'hFA44;
defparam \new_pc[31]~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N18
cycloneive_lcell_comb \new_pc[30]~60 (
// Equation(s):
// \new_pc[30]~60_combout  = (\pc[31]~1_combout  & ((\pc[31]~2_combout  & (idex_ifnext_pc_o_30)) # (!\pc[31]~2_combout  & ((idex_ifrdat1_o_30))))) # (!\pc[31]~1_combout  & (((\pc[31]~2_combout ))))

	.dataa(\IDEX|idex_if.next_pc_o [30]),
	.datab(\IDEX|idex_if.rdat1_o [30]),
	.datac(\pc[31]~1_combout ),
	.datad(\pc[31]~2_combout ),
	.cin(gnd),
	.combout(\new_pc[30]~60_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[30]~60 .lut_mask = 16'hAFC0;
defparam \new_pc[30]~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N8
cycloneive_lcell_comb \new_pc[30]~61 (
// Equation(s):
// \new_pc[30]~61_combout  = (\pc[31]~1_combout  & (((\new_pc[30]~60_combout )))) # (!\pc[31]~1_combout  & ((\new_pc[30]~60_combout  & ((\Add1~56_combout ))) # (!\new_pc[30]~60_combout  & (\nextpc[30]~56_combout ))))

	.dataa(\nextpc[30]~56_combout ),
	.datab(\Add1~56_combout ),
	.datac(\pc[31]~1_combout ),
	.datad(\new_pc[30]~60_combout ),
	.cin(gnd),
	.combout(\new_pc[30]~61_combout ),
	.cout());
// synopsys translate_off
defparam \new_pc[30]~61 .lut_mask = 16'hFC0A;
defparam \new_pc[30]~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y29_N21
dffeas \dpif.halt~_Duplicate_1 (
	.clk(CLK),
	.d(\dpif.halt~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\dpif.halt~_Duplicate_1_q ),
	.prn(vcc));
// synopsys translate_off
defparam \dpif.halt~_Duplicate_1 .is_wysiwyg = "true";
defparam \dpif.halt~_Duplicate_1 .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y29_N20
cycloneive_lcell_comb \dpif.halt~0 (
// Equation(s):
// \dpif.halt~0_combout  = (\dpif.halt~_Duplicate_1_q ) # (exmem_ifhalt_o)

	.dataa(gnd),
	.datab(gnd),
	.datac(\dpif.halt~_Duplicate_1_q ),
	.datad(\EXMEM|exmem_if.halt_o~q ),
	.cin(gnd),
	.combout(\dpif.halt~0_combout ),
	.cout());
// synopsys translate_off
defparam \dpif.halt~0 .lut_mask = 16'hFFF0;
defparam \dpif.halt~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module alu_file (
	idex_ifaluop_o_1,
	port_b,
	fuifrtReplace_1,
	port_b1,
	always0,
	rdat1_1,
	port_b2,
	port_b3,
	fuifrtReplace_0,
	port_b4,
	rdat1_0,
	idex_ifaluop_o_2,
	rdat1_2,
	rdat1_4,
	mem_data,
	rdat1_41,
	rdat1_3,
	mem_data1,
	rdat1_31,
	port_b5,
	fuifrtReplace_2,
	port_b6,
	rdat1_8,
	rdat1_7,
	rdat1_6,
	rdat1_5,
	port_b7,
	rdat1_16,
	rdat1_15,
	rdat1_14,
	rdat1_13,
	rdat1_12,
	rdat1_11,
	rdat1_10,
	rdat1_9,
	port_b8,
	rdat1_311,
	rdat1_29,
	rdat1_30,
	rdat1_28,
	rdat1_26,
	rdat1_27,
	rdat1_25,
	rdat1_24,
	rdat1_22,
	rdat1_23,
	rdat1_21,
	rdat1_20,
	rdat1_18,
	rdat1_19,
	rdat1_17,
	port_b9,
	fuifrtReplace_31,
	port_b10,
	port_b11,
	fuifrtReplace_16,
	port_b12,
	port_b13,
	fuifrtReplace_17,
	port_b14,
	port_b15,
	fuifrtReplace_18,
	port_b16,
	port_b17,
	fuifrtReplace_19,
	port_b18,
	port_b19,
	fuifrtReplace_20,
	port_b20,
	port_b21,
	fuifrtReplace_21,
	port_b22,
	port_b23,
	fuifrtReplace_22,
	port_b24,
	port_b25,
	fuifrtReplace_23,
	port_b26,
	port_b27,
	fuifrtReplace_24,
	port_b28,
	port_b29,
	fuifrtReplace_25,
	port_b30,
	port_b31,
	fuifrtReplace_26,
	port_b32,
	port_b33,
	fuifrtReplace_5,
	port_b34,
	port_b35,
	fuifrtReplace_6,
	port_b36,
	port_b37,
	fuifrtReplace_7,
	port_b38,
	port_b39,
	fuifrtReplace_8,
	port_b40,
	port_b41,
	fuifrtReplace_27,
	port_b42,
	port_b43,
	fuifrtReplace_28,
	port_b44,
	port_b45,
	fuifrtReplace_29,
	port_b46,
	port_b47,
	fuifrtReplace_30,
	port_b48,
	port_b49,
	fuifrtReplace_9,
	port_b50,
	port_b51,
	fuifrtReplace_14,
	port_b52,
	fuifrtReplace_15,
	port_b53,
	port_b54,
	fuifrtReplace_10,
	port_b55,
	port_b56,
	fuifrtReplace_11,
	port_b57,
	port_b58,
	fuifrtReplace_12,
	port_b59,
	fuifrtReplace_13,
	port_b60,
	idex_ifaluop_o_0,
	idex_ifaluop_o_3,
	myifout_1,
	myifout_6,
	myifout_4,
	port_b61,
	port_b62,
	myifout_24,
	myifout_26,
	myifout_25,
	myifout_27,
	myifout_5,
	myifout_7,
	myifout_13,
	myifout_9,
	myifout_8,
	myifout_14,
	myifout_12,
	myifout_15,
	myifout_10,
	myifout_11,
	myifout_23,
	myifout_16,
	myifout_17,
	myifout_18,
	myifout_19,
	myifout_30,
	myifout_21,
	myifnegative,
	myifout_22,
	myifout_20,
	myifout_0,
	Equal10,
	myifout_28,
	myifout_29,
	myifout_2,
	myifout_3,
	myifout_31,
	myifout_210,
	Equal101,
	myifout_32,
	devpor,
	devclrn,
	devoe);
input 	idex_ifaluop_o_1;
input 	port_b;
input 	fuifrtReplace_1;
input 	port_b1;
input 	always0;
input 	rdat1_1;
input 	port_b2;
input 	port_b3;
input 	fuifrtReplace_0;
input 	port_b4;
input 	rdat1_0;
input 	idex_ifaluop_o_2;
input 	rdat1_2;
input 	rdat1_4;
input 	mem_data;
input 	rdat1_41;
input 	rdat1_3;
input 	mem_data1;
input 	rdat1_31;
input 	port_b5;
input 	fuifrtReplace_2;
input 	port_b6;
input 	rdat1_8;
input 	rdat1_7;
input 	rdat1_6;
input 	rdat1_5;
input 	port_b7;
input 	rdat1_16;
input 	rdat1_15;
input 	rdat1_14;
input 	rdat1_13;
input 	rdat1_12;
input 	rdat1_11;
input 	rdat1_10;
input 	rdat1_9;
input 	port_b8;
input 	rdat1_311;
input 	rdat1_29;
input 	rdat1_30;
input 	rdat1_28;
input 	rdat1_26;
input 	rdat1_27;
input 	rdat1_25;
input 	rdat1_24;
input 	rdat1_22;
input 	rdat1_23;
input 	rdat1_21;
input 	rdat1_20;
input 	rdat1_18;
input 	rdat1_19;
input 	rdat1_17;
input 	port_b9;
input 	fuifrtReplace_31;
input 	port_b10;
input 	port_b11;
input 	fuifrtReplace_16;
input 	port_b12;
input 	port_b13;
input 	fuifrtReplace_17;
input 	port_b14;
input 	port_b15;
input 	fuifrtReplace_18;
input 	port_b16;
input 	port_b17;
input 	fuifrtReplace_19;
input 	port_b18;
input 	port_b19;
input 	fuifrtReplace_20;
input 	port_b20;
input 	port_b21;
input 	fuifrtReplace_21;
input 	port_b22;
input 	port_b23;
input 	fuifrtReplace_22;
input 	port_b24;
input 	port_b25;
input 	fuifrtReplace_23;
input 	port_b26;
input 	port_b27;
input 	fuifrtReplace_24;
input 	port_b28;
input 	port_b29;
input 	fuifrtReplace_25;
input 	port_b30;
input 	port_b31;
input 	fuifrtReplace_26;
input 	port_b32;
input 	port_b33;
input 	fuifrtReplace_5;
input 	port_b34;
input 	port_b35;
input 	fuifrtReplace_6;
input 	port_b36;
input 	port_b37;
input 	fuifrtReplace_7;
input 	port_b38;
input 	port_b39;
input 	fuifrtReplace_8;
input 	port_b40;
input 	port_b41;
input 	fuifrtReplace_27;
input 	port_b42;
input 	port_b43;
input 	fuifrtReplace_28;
input 	port_b44;
input 	port_b45;
input 	fuifrtReplace_29;
input 	port_b46;
input 	port_b47;
input 	fuifrtReplace_30;
input 	port_b48;
input 	port_b49;
input 	fuifrtReplace_9;
input 	port_b50;
input 	port_b51;
input 	fuifrtReplace_14;
input 	port_b52;
input 	fuifrtReplace_15;
input 	port_b53;
input 	port_b54;
input 	fuifrtReplace_10;
input 	port_b55;
input 	port_b56;
input 	fuifrtReplace_11;
input 	port_b57;
input 	port_b58;
input 	fuifrtReplace_12;
input 	port_b59;
input 	fuifrtReplace_13;
input 	port_b60;
input 	idex_ifaluop_o_0;
input 	idex_ifaluop_o_3;
output 	myifout_1;
output 	myifout_6;
output 	myifout_4;
input 	port_b61;
input 	port_b62;
output 	myifout_24;
output 	myifout_26;
output 	myifout_25;
output 	myifout_27;
output 	myifout_5;
output 	myifout_7;
output 	myifout_13;
output 	myifout_9;
output 	myifout_8;
output 	myifout_14;
output 	myifout_12;
output 	myifout_15;
output 	myifout_10;
output 	myifout_11;
output 	myifout_23;
output 	myifout_16;
output 	myifout_17;
output 	myifout_18;
output 	myifout_19;
output 	myifout_30;
output 	myifout_21;
output 	myifnegative;
output 	myifout_22;
output 	myifout_20;
output 	myifout_0;
output 	Equal10;
output 	myifout_28;
output 	myifout_29;
output 	myifout_2;
output 	myifout_3;
output 	myifout_31;
output 	myifout_210;
output 	Equal101;
output 	myifout_32;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~32_combout ;
wire \Add0~16_combout ;
wire \Add0~18_combout ;
wire \Add0~26_combout ;
wire \Add0~28_combout ;
wire \Add0~46_combout ;
wire \LessThan0~1_cout ;
wire \LessThan0~3_cout ;
wire \LessThan0~5_cout ;
wire \LessThan0~7_cout ;
wire \LessThan0~9_cout ;
wire \LessThan0~11_cout ;
wire \LessThan0~13_cout ;
wire \LessThan0~15_cout ;
wire \LessThan0~17_cout ;
wire \LessThan0~19_cout ;
wire \LessThan0~21_cout ;
wire \LessThan0~23_cout ;
wire \LessThan0~25_cout ;
wire \LessThan0~27_cout ;
wire \LessThan0~29_cout ;
wire \LessThan0~31_cout ;
wire \LessThan0~33_cout ;
wire \LessThan0~35_cout ;
wire \LessThan0~37_cout ;
wire \LessThan0~39_cout ;
wire \LessThan0~41_cout ;
wire \LessThan0~43_cout ;
wire \LessThan0~45_cout ;
wire \LessThan0~47_cout ;
wire \LessThan0~49_cout ;
wire \LessThan0~51_cout ;
wire \LessThan0~53_cout ;
wire \LessThan0~55_cout ;
wire \LessThan0~57_cout ;
wire \LessThan0~59_cout ;
wire \LessThan0~61_cout ;
wire \LessThan0~62_combout ;
wire \ShiftLeft0~3_combout ;
wire \ShiftLeft0~6_combout ;
wire \ShiftLeft0~14_combout ;
wire \ShiftRight0~32_combout ;
wire \ShiftRight0~34_combout ;
wire \myif.out[6]~18_combout ;
wire \ShiftRight0~57_combout ;
wire \ShiftRight0~66_combout ;
wire \ShiftLeft0~31_combout ;
wire \out~13_combout ;
wire \ShiftLeft0~62_combout ;
wire \ShiftLeft0~63_combout ;
wire \ShiftLeft0~79_combout ;
wire \ShiftLeft0~80_combout ;
wire \ShiftLeft0~81_combout ;
wire \myif.out[7]~73_combout ;
wire \myif.out[7]~74_combout ;
wire \ShiftRight0~91_combout ;
wire \ShiftRight0~95_combout ;
wire \ShiftLeft0~95_combout ;
wire \out~44_combout ;
wire \out~49_combout ;
wire \myif.out[17]~166_combout ;
wire \out~57_combout ;
wire \myif.out[19]~188_combout ;
wire \myif.out[30]~197_combout ;
wire \out~61_combout ;
wire \myif.out[21]~212_combout ;
wire \myif.negative~3_combout ;
wire \myif.negative~4_combout ;
wire \out~65_combout ;
wire \out~71_combout ;
wire \ShiftRight0~106_combout ;
wire \ShiftRight0~108_combout ;
wire \ShiftRight0~109_combout ;
wire \ShiftRight0~110_combout ;
wire \myif.out[0]~233_combout ;
wire \myif.out[0]~234_combout ;
wire \out~79_combout ;
wire \myif.out[1]~10_combout ;
wire \myif.out[1]~11_combout ;
wire \ShiftLeft0~4_combout ;
wire \ShiftLeft0~7_combout ;
wire \ShiftLeft0~5_combout ;
wire \ShiftLeft0~8_combout ;
wire \ShiftLeft0~9_combout ;
wire \ShiftLeft0~10_combout ;
wire \ShiftLeft0~2_combout ;
wire \ShiftLeft0~11_combout ;
wire \myif.out[1]~13_combout ;
wire \Add0~1 ;
wire \Add0~2_combout ;
wire \myif.out[1]~12_combout ;
wire \myif.out[1]~14_combout ;
wire \myif.out[1]~8_combout ;
wire \myif.out[1]~6_combout ;
wire \Add1~1 ;
wire \Add1~2_combout ;
wire \myif.out[1]~7_combout ;
wire \ShiftRight0~19_combout ;
wire \ShiftRight0~20_combout ;
wire \ShiftRight0~21_combout ;
wire \ShiftRight0~22_combout ;
wire \ShiftRight0~27_combout ;
wire \ShiftRight0~26_combout ;
wire \ShiftRight0~28_combout ;
wire \ShiftRight0~24_combout ;
wire \ShiftRight0~23_combout ;
wire \ShiftRight0~25_combout ;
wire \ShiftRight0~29_combout ;
wire \ShiftRight0~30_combout ;
wire \ShiftRight0~12_combout ;
wire \ShiftRight0~13_combout ;
wire \ShiftRight0~14_combout ;
wire \ShiftRight0~9_combout ;
wire \ShiftRight0~10_combout ;
wire \ShiftRight0~11_combout ;
wire \ShiftRight0~15_combout ;
wire \ShiftRight0~2_combout ;
wire \ShiftRight0~3_combout ;
wire \ShiftRight0~4_combout ;
wire \ShiftRight0~5_combout ;
wire \ShiftRight0~6_combout ;
wire \ShiftRight0~7_combout ;
wire \ShiftRight0~8_combout ;
wire \ShiftRight0~16_combout ;
wire \ShiftRight0~31_combout ;
wire \myif.out[1]~9_combout ;
wire \out~9_combout ;
wire \Add0~3 ;
wire \Add0~5 ;
wire \Add0~7 ;
wire \Add0~9 ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \out~10_combout ;
wire \ShiftLeft0~18_combout ;
wire \ShiftLeft0~17_combout ;
wire \ShiftLeft0~19_combout ;
wire \ShiftLeft0~20_combout ;
wire \myif.out[13]~23_combout ;
wire \myif.out[6]~24_combout ;
wire \myif.out[6]~25_combout ;
wire \out~8_combout ;
wire \Add1~3 ;
wire \Add1~5 ;
wire \Add1~7 ;
wire \Add1~9 ;
wire \Add1~11 ;
wire \Add1~12_combout ;
wire \myif.out[5]~20_combout ;
wire \myif.out[5]~16_combout ;
wire \ShiftRight0~35_combout ;
wire \ShiftRight0~36_combout ;
wire \ShiftRight0~37_combout ;
wire \ShiftRight0~38_combout ;
wire \ShiftRight0~45_combout ;
wire \ShiftRight0~46_combout ;
wire \ShiftRight0~47_combout ;
wire \ShiftRight0~49_combout ;
wire \ShiftRight0~48_combout ;
wire \ShiftRight0~50_combout ;
wire \ShiftRight0~51_combout ;
wire \ShiftLeft0~13_combout ;
wire \ShiftRight0~53_combout ;
wire \myif.out[6]~19_combout ;
wire \myif.out[6]~21_combout ;
wire \myif.out[6]~22_combout ;
wire \Add1~8_combout ;
wire \out~77_combout ;
wire \myif.out[5]~17_combout ;
wire \ShiftRight0~43_combout ;
wire \ShiftRight0~60_combout ;
wire \ShiftRight0~55_combout ;
wire \ShiftRight0~56_combout ;
wire \ShiftRight0~58_combout ;
wire \myif.out[4]~27_combout ;
wire \ShiftRight0~61_combout ;
wire \ShiftRight0~62_combout ;
wire \ShiftRight0~63_combout ;
wire \ShiftRight0~64_combout ;
wire \ShiftRight0~65_combout ;
wire \ShiftRight0~68_combout ;
wire \myif.out[4]~28_combout ;
wire \myif.out[4]~29_combout ;
wire \myif.out[4]~30_combout ;
wire \out~78_combout ;
wire \Add0~8_combout ;
wire \ShiftLeft0~22_combout ;
wire \ShiftLeft0~23_combout ;
wire \ShiftLeft0~21_combout ;
wire \ShiftLeft0~24_combout ;
wire \myif.out[4]~31_combout ;
wire \myif.out[4]~32_combout ;
wire \Add0~13 ;
wire \Add0~15 ;
wire \Add0~17 ;
wire \Add0~19 ;
wire \Add0~21 ;
wire \Add0~23 ;
wire \Add0~25 ;
wire \Add0~27 ;
wire \Add0~29 ;
wire \Add0~31 ;
wire \Add0~33 ;
wire \Add0~35 ;
wire \Add0~37 ;
wire \Add0~39 ;
wire \Add0~41 ;
wire \Add0~43 ;
wire \Add0~45 ;
wire \Add0~47 ;
wire \Add0~48_combout ;
wire \out~12_combout ;
wire \ShiftLeft0~34_combout ;
wire \ShiftLeft0~35_combout ;
wire \ShiftLeft0~36_combout ;
wire \myif.out[24]~36_combout ;
wire \ShiftLeft0~25_combout ;
wire \ShiftLeft0~26_combout ;
wire \ShiftLeft0~27_combout ;
wire \ShiftLeft0~28_combout ;
wire \ShiftLeft0~30_combout ;
wire \ShiftLeft0~37_combout ;
wire \ShiftLeft0~38_combout ;
wire \ShiftLeft0~39_combout ;
wire \ShiftLeft0~40_combout ;
wire \myif.out[24]~37_combout ;
wire \myif.out[24]~38_combout ;
wire \myif.out[24]~39_combout ;
wire \out~11_combout ;
wire \Add1~13 ;
wire \Add1~15 ;
wire \Add1~17 ;
wire \Add1~19 ;
wire \Add1~21 ;
wire \Add1~23 ;
wire \Add1~25 ;
wire \Add1~27 ;
wire \Add1~29 ;
wire \Add1~31 ;
wire \Add1~33 ;
wire \Add1~35 ;
wire \Add1~37 ;
wire \Add1~39 ;
wire \Add1~41 ;
wire \Add1~43 ;
wire \Add1~45 ;
wire \Add1~47 ;
wire \Add1~48_combout ;
wire \ShiftRight0~52_combout ;
wire \ShiftRight0~67_combout ;
wire \ShiftRight0~69_combout ;
wire \myif.out[24]~34_combout ;
wire \myif.out[24]~35_combout ;
wire \out~14_combout ;
wire \ShiftRight0~70_combout ;
wire \ShiftRight0~71_combout ;
wire \myif.out[26]~41_combout ;
wire \Add1~49 ;
wire \Add1~51 ;
wire \Add1~52_combout ;
wire \myif.out[26]~42_combout ;
wire \out~15_combout ;
wire \out~16_combout ;
wire \ShiftLeft0~15_combout ;
wire \ShiftLeft0~16_combout ;
wire \ShiftLeft0~52_combout ;
wire \ShiftLeft0~53_combout ;
wire \ShiftLeft0~54_combout ;
wire \ShiftLeft0~44_combout ;
wire \ShiftLeft0~45_combout ;
wire \ShiftLeft0~46_combout ;
wire \ShiftLeft0~47_combout ;
wire \ShiftLeft0~48_combout ;
wire \myif.out[26]~43_combout ;
wire \myif.out[26]~44_combout ;
wire \myif.out[26]~45_combout ;
wire \Add0~49 ;
wire \Add0~51 ;
wire \Add0~52_combout ;
wire \myif.out[26]~46_combout ;
wire \out~17_combout ;
wire \ShiftRight0~17_combout ;
wire \ShiftRight0~18_combout ;
wire \ShiftRight0~72_combout ;
wire \myif.out[25]~48_combout ;
wire \Add1~50_combout ;
wire \myif.out[25]~49_combout ;
wire \Add0~50_combout ;
wire \out~18_combout ;
wire \out~19_combout ;
wire \ShiftLeft0~64_combout ;
wire \ShiftLeft0~65_combout ;
wire \myif.out[25]~50_combout ;
wire \ShiftLeft0~55_combout ;
wire \ShiftLeft0~56_combout ;
wire \ShiftLeft0~57_combout ;
wire \ShiftLeft0~58_combout ;
wire \ShiftLeft0~59_combout ;
wire \ShiftLeft0~60_combout ;
wire \ShiftLeft0~61_combout ;
wire \ShiftLeft0~67_combout ;
wire \ShiftLeft0~68_combout ;
wire \ShiftLeft0~70_combout ;
wire \ShiftLeft0~71_combout ;
wire \ShiftLeft0~72_combout ;
wire \ShiftLeft0~73_combout ;
wire \myif.out[25]~51_combout ;
wire \myif.out[25]~52_combout ;
wire \myif.out[25]~53_combout ;
wire \out~21_combout ;
wire \out~22_combout ;
wire \ShiftLeft0~12_combout ;
wire \ShiftLeft0~66_combout ;
wire \ShiftLeft0~85_combout ;
wire \ShiftLeft0~69_combout ;
wire \ShiftLeft0~82_combout ;
wire \ShiftLeft0~83_combout ;
wire \ShiftLeft0~84_combout ;
wire \ShiftLeft0~86_combout ;
wire \ShiftLeft0~75_combout ;
wire \ShiftLeft0~76_combout ;
wire \ShiftLeft0~32_combout ;
wire \ShiftLeft0~77_combout ;
wire \ShiftLeft0~78_combout ;
wire \myif.out[27]~57_combout ;
wire \myif.out[27]~58_combout ;
wire \myif.out[27]~59_combout ;
wire \Add0~53 ;
wire \Add0~54_combout ;
wire \myif.out[27]~60_combout ;
wire \out~20_combout ;
wire \Add1~53 ;
wire \Add1~54_combout ;
wire \ShiftRight0~74_combout ;
wire \ShiftRight0~75_combout ;
wire \ShiftRight0~76_combout ;
wire \myif.out[27]~55_combout ;
wire \myif.out[27]~56_combout ;
wire \out~24_combout ;
wire \ShiftLeft0~87_combout ;
wire \ShiftLeft0~88_combout ;
wire \out~25_combout ;
wire \myif.out[5]~66_combout ;
wire \Add0~10_combout ;
wire \myif.out[5]~67_combout ;
wire \Add1~10_combout ;
wire \out~23_combout ;
wire \myif.out[5]~62_combout ;
wire \ShiftRight0~77_combout ;
wire \ShiftRight0~78_combout ;
wire \ShiftRight0~79_combout ;
wire \myif.out[5]~63_combout ;
wire \myif.out[5]~64_combout ;
wire \myif.out[5]~65_combout ;
wire \ShiftLeft0~89_combout ;
wire \Add0~14_combout ;
wire \myif.out[7]~75_combout ;
wire \myif.out[7]~76_combout ;
wire \myif.out[7]~77_combout ;
wire \myif.out[7]~78_combout ;
wire \myif.out[7]~79_combout ;
wire \myif.out[7]~80_combout ;
wire \Add1~14_combout ;
wire \out~26_combout ;
wire \ShiftRight0~80_combout ;
wire \ShiftRight0~86_combout ;
wire \ShiftRight0~81_combout ;
wire \ShiftRight0~33_combout ;
wire \ShiftRight0~82_combout ;
wire \ShiftRight0~83_combout ;
wire \ShiftRight0~84_combout ;
wire \ShiftRight0~85_combout ;
wire \myif.out[7]~69_combout ;
wire \myif.out[7]~70_combout ;
wire \myif.out[7]~71_combout ;
wire \myif.out[7]~72_combout ;
wire \out~27_combout ;
wire \myif.out[13]~87_combout ;
wire \myif.out[13]~82_combout ;
wire \myif.out[13]~83_combout ;
wire \myif.out[13]~84_combout ;
wire \myif.out[13]~85_combout ;
wire \myif.out[13]~86_combout ;
wire \myif.out[13]~88_combout ;
wire \Add1~26_combout ;
wire \out~28_combout ;
wire \out~29_combout ;
wire \ShiftLeft0~90_combout ;
wire \ShiftLeft0~91_combout ;
wire \myif.out[13]~89_combout ;
wire \myif.out[13]~90_combout ;
wire \myif.out[13]~91_combout ;
wire \out~30_combout ;
wire \Add1~18_combout ;
wire \myif.out[9]~93_combout ;
wire \myif.out[9]~94_combout ;
wire \out~32_combout ;
wire \myif.out[9]~95_combout ;
wire \out~31_combout ;
wire \myif.out[9]~96_combout ;
wire \myif.out[9]~97_combout ;
wire \ShiftRight0~40_combout ;
wire \ShiftRight0~42_combout ;
wire \ShiftRight0~54_combout ;
wire \ShiftRight0~92_combout ;
wire \ShiftRight0~93_combout ;
wire \myif.out[8]~99_combout ;
wire \myif.out[8]~100_combout ;
wire \Add1~16_combout ;
wire \out~35_combout ;
wire \myif.out[8]~101_combout ;
wire \out~34_combout ;
wire \myif.out[8]~102_combout ;
wire \myif.out[8]~103_combout ;
wire \out~33_combout ;
wire \Add1~28_combout ;
wire \out~36_combout ;
wire \out~37_combout ;
wire \out~38_combout ;
wire \ShiftLeft0~92_combout ;
wire \ShiftLeft0~93_combout ;
wire \ShiftLeft0~94_combout ;
wire \myif.out[14]~107_combout ;
wire \myif.out[14]~108_combout ;
wire \ShiftRight0~94_combout ;
wire \myif.out[14]~105_combout ;
wire \myif.out[14]~106_combout ;
wire \myif.out[14]~109_combout ;
wire \out~39_combout ;
wire \Add1~24_combout ;
wire \Add0~24_combout ;
wire \out~40_combout ;
wire \ShiftLeft0~96_combout ;
wire \ShiftLeft0~97_combout ;
wire \out~41_combout ;
wire \myif.out[12]~113_combout ;
wire \myif.out[12]~114_combout ;
wire \myif.out[12]~115_combout ;
wire \myif.out[12]~111_combout ;
wire \myif.out[12]~112_combout ;
wire \out~42_combout ;
wire \Add1~30_combout ;
wire \ShiftRight0~87_combout ;
wire \ShiftRight0~88_combout ;
wire \ShiftRight0~89_combout ;
wire \ShiftRight0~73_combout ;
wire \ShiftRight0~96_combout ;
wire \myif.out[15]~117_combout ;
wire \myif.out[15]~118_combout ;
wire \out~43_combout ;
wire \Add0~30_combout ;
wire \ShiftLeft0~98_combout ;
wire \ShiftLeft0~99_combout ;
wire \ShiftLeft0~100_combout ;
wire \myif.out[15]~119_combout ;
wire \myif.out[15]~120_combout ;
wire \myif.out[15]~121_combout ;
wire \out~45_combout ;
wire \ShiftRight0~98_combout ;
wire \ShiftRight0~39_combout ;
wire \ShiftRight0~41_combout ;
wire \ShiftRight0~97_combout ;
wire \myif.out[10]~123_combout ;
wire \myif.out[10]~124_combout ;
wire \Add1~20_combout ;
wire \out~46_combout ;
wire \Add0~20_combout ;
wire \out~47_combout ;
wire \myif.out[10]~125_combout ;
wire \myif.out[10]~126_combout ;
wire \myif.out[10]~127_combout ;
wire \Add1~22_combout ;
wire \out~48_combout ;
wire \ShiftRight0~100_combout ;
wire \myif.out[11]~129_combout ;
wire \myif.out[11]~130_combout ;
wire \Add0~22_combout ;
wire \out~50_combout ;
wire \myif.out[11]~131_combout ;
wire \myif.out[11]~132_combout ;
wire \myif.out[11]~133_combout ;
wire \myif.out[23]~135_combout ;
wire \out~51_combout ;
wire \myif.out[23]~136_combout ;
wire \ShiftLeft0~42_combout ;
wire \ShiftLeft0~74_combout ;
wire \ShiftLeft0~101_combout ;
wire \myif.out[23]~137_combout ;
wire \myif.out[23]~150_combout ;
wire \myif.out[23]~138_combout ;
wire \Add1~46_combout ;
wire \myif.out[23]~140_combout ;
wire \myif.out[23]~141_combout ;
wire \myif.out[23]~151_combout ;
wire \myif.out[23]~139_combout ;
wire \myif.out[23]~147_combout ;
wire \myif.out[23]~142_combout ;
wire \myif.out[23]~143_combout ;
wire \ShiftRight0~90_combout ;
wire \myif.out[23]~144_combout ;
wire \myif.out[23]~145_combout ;
wire \myif.out[23]~146_combout ;
wire \myif.out[23]~148_combout ;
wire \myif.out[23]~149_combout ;
wire \Add0~32_combout ;
wire \out~54_combout ;
wire \out~53_combout ;
wire \myif.out[16]~155_combout ;
wire \myif.out[16]~156_combout ;
wire \out~52_combout ;
wire \ShiftRight0~101_combout ;
wire \ShiftRight0~102_combout ;
wire \myif.out[16]~153_combout ;
wire \myif.out[16]~154_combout ;
wire \myif.out[16]~157_combout ;
wire \out~55_combout ;
wire \myif.out[17]~159_combout ;
wire \myif.out[17]~160_combout ;
wire \Add0~34_combout ;
wire \Add1~34_combout ;
wire \myif.out[17]~163_combout ;
wire \myif.out[17]~164_combout ;
wire \myif.out[17]~161_combout ;
wire \myif.out[17]~162_combout ;
wire \myif.out[17]~165_combout ;
wire \myif.out[17]~170_combout ;
wire \myif.out[17]~167_combout ;
wire \myif.out[17]~168_combout ;
wire \myif.out[17]~169_combout ;
wire \myif.out[17]~171_combout ;
wire \myif.out[17]~172_combout ;
wire \myif.out[17]~173_combout ;
wire \out~58_combout ;
wire \Add0~36_combout ;
wire \out~56_combout ;
wire \ShiftRight0~103_combout ;
wire \myif.out[18]~175_combout ;
wire \Add1~36_combout ;
wire \myif.out[18]~176_combout ;
wire \ShiftLeft0~103_combout ;
wire \myif.out[18]~177_combout ;
wire \myif.out[18]~178_combout ;
wire \myif.out[18]~179_combout ;
wire \myif.out[19]~183_combout ;
wire \Add0~38_combout ;
wire \Add1~38_combout ;
wire \myif.out[19]~185_combout ;
wire \myif.out[19]~186_combout ;
wire \myif.out[19]~195_combout ;
wire \out~59_combout ;
wire \myif.out[19]~181_combout ;
wire \myif.out[19]~182_combout ;
wire \myif.out[19]~184_combout ;
wire \myif.out[19]~187_combout ;
wire \myif.out[19]~192_combout ;
wire \ShiftRight0~104_combout ;
wire \ShiftRight0~105_combout ;
wire \myif.out[19]~189_combout ;
wire \myif.out[19]~190_combout ;
wire \myif.out[19]~191_combout ;
wire \myif.out[19]~193_combout ;
wire \myif.out[19]~194_combout ;
wire \out~62_combout ;
wire \Add0~55 ;
wire \Add0~57 ;
wire \Add0~59 ;
wire \Add0~60_combout ;
wire \ShiftLeft0~41_combout ;
wire \ShiftLeft0~43_combout ;
wire \ShiftLeft0~105_combout ;
wire \myif.negative~0_combout ;
wire \ShiftLeft0~50_combout ;
wire \ShiftLeft0~49_combout ;
wire \ShiftLeft0~51_combout ;
wire \ShiftLeft0~104_combout ;
wire \myif.out[30]~199_combout ;
wire \myif.out[30]~200_combout ;
wire \myif.out[30]~201_combout ;
wire \myif.out[30]~202_combout ;
wire \Add1~55 ;
wire \Add1~57 ;
wire \Add1~59 ;
wire \Add1~60_combout ;
wire \out~60_combout ;
wire \myif.out[30]~198_combout ;
wire \myif.out[30]~203_combout ;
wire \Add1~42_combout ;
wire \myif.out[21]~207_combout ;
wire \myif.out[21]~209_combout ;
wire \Add0~42_combout ;
wire \myif.out[21]~210_combout ;
wire \myif.out[21]~219_combout ;
wire \ShiftLeft0~106_combout ;
wire \out~63_combout ;
wire \myif.out[21]~205_combout ;
wire \myif.out[21]~206_combout ;
wire \myif.out[21]~208_combout ;
wire \myif.out[21]~211_combout ;
wire \myif.out[21]~216_combout ;
wire \myif.out[21]~213_combout ;
wire \myif.out[21]~214_combout ;
wire \myif.out[21]~215_combout ;
wire \myif.out[21]~217_combout ;
wire \myif.out[21]~218_combout ;
wire \out~66_combout ;
wire \out~64_combout ;
wire \myif.negative~1_combout ;
wire \Add1~61 ;
wire \Add1~62_combout ;
wire \myif.negative~2_combout ;
wire \myif.negative~5_combout ;
wire \myif.negative~6_combout ;
wire \Add0~61 ;
wire \Add0~62_combout ;
wire \myif.negative~7_combout ;
wire \out~69_combout ;
wire \out~68_combout ;
wire \myif.out[22]~223_combout ;
wire \myif.out[22]~224_combout ;
wire \out~67_combout ;
wire \myif.out[22]~221_combout ;
wire \Add1~44_combout ;
wire \myif.out[22]~222_combout ;
wire \myif.out[22]~225_combout ;
wire \Add0~44_combout ;
wire \out~72_combout ;
wire \Add0~40_combout ;
wire \ShiftLeft0~29_combout ;
wire \ShiftLeft0~33_combout ;
wire \ShiftLeft0~108_combout ;
wire \myif.out[20]~229_combout ;
wire \myif.out[20]~230_combout ;
wire \out~70_combout ;
wire \myif.out[20]~227_combout ;
wire \Add1~40_combout ;
wire \myif.out[20]~228_combout ;
wire \myif.out[20]~231_combout ;
wire \Add1~0_combout ;
wire \Add0~0_combout ;
wire \myif.out[0]~237_combout ;
wire \out~73_combout ;
wire \myif.out[0]~238_combout ;
wire \ShiftLeft0~102_combout ;
wire \myif.out[0]~235_combout ;
wire \ShiftRight0~111_combout ;
wire \myif.out[0]~236_combout ;
wire \LessThan1~1_cout ;
wire \LessThan1~3_cout ;
wire \LessThan1~5_cout ;
wire \LessThan1~7_cout ;
wire \LessThan1~9_cout ;
wire \LessThan1~11_cout ;
wire \LessThan1~13_cout ;
wire \LessThan1~15_cout ;
wire \LessThan1~17_cout ;
wire \LessThan1~19_cout ;
wire \LessThan1~21_cout ;
wire \LessThan1~23_cout ;
wire \LessThan1~25_cout ;
wire \LessThan1~27_cout ;
wire \LessThan1~29_cout ;
wire \LessThan1~31_cout ;
wire \LessThan1~33_cout ;
wire \LessThan1~35_cout ;
wire \LessThan1~37_cout ;
wire \LessThan1~39_cout ;
wire \LessThan1~41_cout ;
wire \LessThan1~43_cout ;
wire \LessThan1~45_cout ;
wire \LessThan1~47_cout ;
wire \LessThan1~49_cout ;
wire \LessThan1~51_cout ;
wire \LessThan1~53_cout ;
wire \LessThan1~55_cout ;
wire \LessThan1~57_cout ;
wire \LessThan1~59_cout ;
wire \LessThan1~61_cout ;
wire \LessThan1~62_combout ;
wire \myif.out[0]~294_combout ;
wire \myif.out[0]~295_combout ;
wire \Equal10~8_combout ;
wire \Equal10~9_combout ;
wire \Equal10~4_combout ;
wire \Equal10~3_combout ;
wire \Equal10~6_combout ;
wire \Equal10~5_combout ;
wire \Equal10~7_combout ;
wire \Equal10~1_combout ;
wire \Equal10~0_combout ;
wire \Equal10~2_combout ;
wire \myif.out[3]~246_combout ;
wire \myif.out[28]~247_combout ;
wire \Add1~56_combout ;
wire \out~75_combout ;
wire \myif.out[28]~249_combout ;
wire \myif.out[28]~292_combout ;
wire \myif.out[28]~293_combout ;
wire \out~74_combout ;
wire \myif.out[3]~240_combout ;
wire \myif.out[3]~241_combout ;
wire \myif.out[28]~242_combout ;
wire \myif.out[28]~243_combout ;
wire \myif.out[28]~244_combout ;
wire \myif.out[28]~248_combout ;
wire \Add0~56_combout ;
wire \myif.out[28]~251_combout ;
wire \myif.out[5]~245_combout ;
wire \myif.out[28]~250_combout ;
wire \myif.out[28]~290_combout ;
wire \myif.out[29]~260_combout ;
wire \myif.out[29]~261_combout ;
wire \Add1~58_combout ;
wire \myif.out[29]~253_combout ;
wire \myif.out[29]~262_combout ;
wire \myif.out[29]~263_combout ;
wire \myif.out[29]~259_combout ;
wire \Add0~58_combout ;
wire \myif.out[29]~254_combout ;
wire \ShiftLeft0~107_combout ;
wire \myif.out[29]~255_combout ;
wire \myif.out[29]~256_combout ;
wire \myif.out[29]~257_combout ;
wire \myif.out[29]~258_combout ;
wire \myif.out[3]~273_combout ;
wire \out~76_combout ;
wire \myif.out[2]~265_combout ;
wire \myif.out[2]~266_combout ;
wire \Add0~4_combout ;
wire \myif.out[2]~267_combout ;
wire \myif.out[2]~268_combout ;
wire \myif.out[2]~269_combout ;
wire \myif.out[2]~270_combout ;
wire \myif.out[2]~271_combout ;
wire \myif.out[2]~272_combout ;
wire \Add1~6_combout ;
wire \out~80_combout ;
wire \ShiftRight0~99_combout ;
wire \ShiftRight0~112_combout ;
wire \myif.out[3]~280_combout ;
wire \myif.out[3]~281_combout ;
wire \myif.out[3]~282_combout ;
wire \myif.out[5]~284_combout ;
wire \Add1~4_combout ;
wire \ShiftRight0~59_combout ;
wire \ShiftRight0~107_combout ;
wire \ShiftRight0~44_combout ;
wire \myif.out[2]~286_combout ;
wire \myif.out[2]~287_combout ;
wire \myif.out[2]~288_combout ;
wire \Equal10~11_combout ;
wire \Add0~6_combout ;
wire \ShiftLeft0~109_combout ;
wire \myif.out[3]~276_combout ;
wire \myif.out[3]~277_combout ;
wire \myif.out[3]~278_combout ;
wire \myif.out[3]~279_combout ;
wire \myif.out[3]~275_combout ;


// Location: LCCOMB_X58_Y33_N0
cycloneive_lcell_comb \Add1~32 (
// Equation(s):
// \Add1~32_combout  = ((\port_b~22_combout  $ (\rdat1[16]~19_combout  $ (\Add1~31 )))) # (GND)
// \Add1~33  = CARRY((\port_b~22_combout  & (\rdat1[16]~19_combout  & !\Add1~31 )) # (!\port_b~22_combout  & ((\rdat1[16]~19_combout ) # (!\Add1~31 ))))

	.dataa(port_b12),
	.datab(rdat1_16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~31 ),
	.combout(\Add1~32_combout ),
	.cout(\Add1~33 ));
// synopsys translate_off
defparam \Add1~32 .lut_mask = 16'h964D;
defparam \Add1~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N16
cycloneive_lcell_comb \Add0~16 (
// Equation(s):
// \Add0~16_combout  = ((\rdat1[8]~11_combout  $ (\port_b~50_combout  $ (!\Add0~15 )))) # (GND)
// \Add0~17  = CARRY((\rdat1[8]~11_combout  & ((\port_b~50_combout ) # (!\Add0~15 ))) # (!\rdat1[8]~11_combout  & (\port_b~50_combout  & !\Add0~15 )))

	.dataa(rdat1_8),
	.datab(port_b40),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
// synopsys translate_off
defparam \Add0~16 .lut_mask = 16'h698E;
defparam \Add0~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N18
cycloneive_lcell_comb \Add0~18 (
// Equation(s):
// \Add0~18_combout  = (\port_b~60_combout  & ((\rdat1[9]~33_combout  & (\Add0~17  & VCC)) # (!\rdat1[9]~33_combout  & (!\Add0~17 )))) # (!\port_b~60_combout  & ((\rdat1[9]~33_combout  & (!\Add0~17 )) # (!\rdat1[9]~33_combout  & ((\Add0~17 ) # (GND)))))
// \Add0~19  = CARRY((\port_b~60_combout  & (!\rdat1[9]~33_combout  & !\Add0~17 )) # (!\port_b~60_combout  & ((!\Add0~17 ) # (!\rdat1[9]~33_combout ))))

	.dataa(port_b50),
	.datab(rdat1_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
// synopsys translate_off
defparam \Add0~18 .lut_mask = 16'h9617;
defparam \Add0~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N26
cycloneive_lcell_comb \Add0~26 (
// Equation(s):
// \Add0~26_combout  = (\port_b~70_combout  & ((\rdat1[13]~25_combout  & (\Add0~25  & VCC)) # (!\rdat1[13]~25_combout  & (!\Add0~25 )))) # (!\port_b~70_combout  & ((\rdat1[13]~25_combout  & (!\Add0~25 )) # (!\rdat1[13]~25_combout  & ((\Add0~25 ) # (GND)))))
// \Add0~27  = CARRY((\port_b~70_combout  & (!\rdat1[13]~25_combout  & !\Add0~25 )) # (!\port_b~70_combout  & ((!\Add0~25 ) # (!\rdat1[13]~25_combout ))))

	.dataa(port_b60),
	.datab(rdat1_13),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout(\Add0~27 ));
// synopsys translate_off
defparam \Add0~26 .lut_mask = 16'h9617;
defparam \Add0~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N28
cycloneive_lcell_comb \Add0~28 (
// Equation(s):
// \Add0~28_combout  = ((\rdat1[14]~23_combout  $ (\port_b~71_combout  $ (!\Add0~27 )))) # (GND)
// \Add0~29  = CARRY((\rdat1[14]~23_combout  & ((\port_b~71_combout ) # (!\Add0~27 ))) # (!\rdat1[14]~23_combout  & (\port_b~71_combout  & !\Add0~27 )))

	.dataa(rdat1_14),
	.datab(port_b61),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~27 ),
	.combout(\Add0~28_combout ),
	.cout(\Add0~29 ));
// synopsys translate_off
defparam \Add0~28 .lut_mask = 16'h698E;
defparam \Add0~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N14
cycloneive_lcell_comb \Add0~46 (
// Equation(s):
// \Add0~46_combout  = (\port_b~36_combout  & ((\rdat1[23]~53_combout  & (\Add0~45  & VCC)) # (!\rdat1[23]~53_combout  & (!\Add0~45 )))) # (!\port_b~36_combout  & ((\rdat1[23]~53_combout  & (!\Add0~45 )) # (!\rdat1[23]~53_combout  & ((\Add0~45 ) # (GND)))))
// \Add0~47  = CARRY((\port_b~36_combout  & (!\rdat1[23]~53_combout  & !\Add0~45 )) # (!\port_b~36_combout  & ((!\Add0~45 ) # (!\rdat1[23]~53_combout ))))

	.dataa(port_b26),
	.datab(rdat1_23),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~45 ),
	.combout(\Add0~46_combout ),
	.cout(\Add0~47 ));
// synopsys translate_off
defparam \Add0~46 .lut_mask = 16'h9617;
defparam \Add0~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N0
cycloneive_lcell_comb \LessThan0~1 (
// Equation(s):
// \LessThan0~1_cout  = CARRY((!\rdat1[0]~3_combout  & \port_b~7_combout ))

	.dataa(rdat1_0),
	.datab(port_b4),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan0~1_cout ));
// synopsys translate_off
defparam \LessThan0~1 .lut_mask = 16'h0044;
defparam \LessThan0~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N2
cycloneive_lcell_comb \LessThan0~3 (
// Equation(s):
// \LessThan0~3_cout  = CARRY((\port_b~4_combout  & (\rdat1[1]~1_combout  & !\LessThan0~1_cout )) # (!\port_b~4_combout  & ((\rdat1[1]~1_combout ) # (!\LessThan0~1_cout ))))

	.dataa(port_b2),
	.datab(rdat1_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~1_cout ),
	.combout(),
	.cout(\LessThan0~3_cout ));
// synopsys translate_off
defparam \LessThan0~3 .lut_mask = 16'h004D;
defparam \LessThan0~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N4
cycloneive_lcell_comb \LessThan0~5 (
// Equation(s):
// \LessThan0~5_cout  = CARRY((\rdat1[2]~5_combout  & (\port_b~10_combout  & !\LessThan0~3_cout )) # (!\rdat1[2]~5_combout  & ((\port_b~10_combout ) # (!\LessThan0~3_cout ))))

	.dataa(rdat1_2),
	.datab(port_b6),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~3_cout ),
	.combout(),
	.cout(\LessThan0~5_cout ));
// synopsys translate_off
defparam \LessThan0~5 .lut_mask = 16'h004D;
defparam \LessThan0~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N6
cycloneive_lcell_comb \LessThan0~7 (
// Equation(s):
// \LessThan0~7_cout  = CARRY((\port_b~14_combout  & (\rdat1[3]~9_combout  & !\LessThan0~5_cout )) # (!\port_b~14_combout  & ((\rdat1[3]~9_combout ) # (!\LessThan0~5_cout ))))

	.dataa(port_b7),
	.datab(rdat1_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~5_cout ),
	.combout(),
	.cout(\LessThan0~7_cout ));
// synopsys translate_off
defparam \LessThan0~7 .lut_mask = 16'h004D;
defparam \LessThan0~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N8
cycloneive_lcell_comb \LessThan0~9 (
// Equation(s):
// \LessThan0~9_cout  = CARRY((\port_b~17_combout  & ((!\LessThan0~7_cout ) # (!\rdat1[4]~7_combout ))) # (!\port_b~17_combout  & (!\rdat1[4]~7_combout  & !\LessThan0~7_cout )))

	.dataa(port_b8),
	.datab(rdat1_41),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~7_cout ),
	.combout(),
	.cout(\LessThan0~9_cout ));
// synopsys translate_off
defparam \LessThan0~9 .lut_mask = 16'h002B;
defparam \LessThan0~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N10
cycloneive_lcell_comb \LessThan0~11 (
// Equation(s):
// \LessThan0~11_cout  = CARRY((\port_b~44_combout  & (\rdat1[5]~17_combout  & !\LessThan0~9_cout )) # (!\port_b~44_combout  & ((\rdat1[5]~17_combout ) # (!\LessThan0~9_cout ))))

	.dataa(port_b34),
	.datab(rdat1_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~9_cout ),
	.combout(),
	.cout(\LessThan0~11_cout ));
// synopsys translate_off
defparam \LessThan0~11 .lut_mask = 16'h004D;
defparam \LessThan0~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N12
cycloneive_lcell_comb \LessThan0~13 (
// Equation(s):
// \LessThan0~13_cout  = CARRY((\rdat1[6]~15_combout  & (\port_b~46_combout  & !\LessThan0~11_cout )) # (!\rdat1[6]~15_combout  & ((\port_b~46_combout ) # (!\LessThan0~11_cout ))))

	.dataa(rdat1_6),
	.datab(port_b36),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~11_cout ),
	.combout(),
	.cout(\LessThan0~13_cout ));
// synopsys translate_off
defparam \LessThan0~13 .lut_mask = 16'h004D;
defparam \LessThan0~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N14
cycloneive_lcell_comb \LessThan0~15 (
// Equation(s):
// \LessThan0~15_cout  = CARRY((\port_b~48_combout  & (\rdat1[7]~13_combout  & !\LessThan0~13_cout )) # (!\port_b~48_combout  & ((\rdat1[7]~13_combout ) # (!\LessThan0~13_cout ))))

	.dataa(port_b38),
	.datab(rdat1_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~13_cout ),
	.combout(),
	.cout(\LessThan0~15_cout ));
// synopsys translate_off
defparam \LessThan0~15 .lut_mask = 16'h004D;
defparam \LessThan0~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N16
cycloneive_lcell_comb \LessThan0~17 (
// Equation(s):
// \LessThan0~17_cout  = CARRY((\port_b~50_combout  & ((!\LessThan0~15_cout ) # (!\rdat1[8]~11_combout ))) # (!\port_b~50_combout  & (!\rdat1[8]~11_combout  & !\LessThan0~15_cout )))

	.dataa(port_b40),
	.datab(rdat1_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~15_cout ),
	.combout(),
	.cout(\LessThan0~17_cout ));
// synopsys translate_off
defparam \LessThan0~17 .lut_mask = 16'h002B;
defparam \LessThan0~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N18
cycloneive_lcell_comb \LessThan0~19 (
// Equation(s):
// \LessThan0~19_cout  = CARRY((\port_b~60_combout  & (\rdat1[9]~33_combout  & !\LessThan0~17_cout )) # (!\port_b~60_combout  & ((\rdat1[9]~33_combout ) # (!\LessThan0~17_cout ))))

	.dataa(port_b50),
	.datab(rdat1_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~17_cout ),
	.combout(),
	.cout(\LessThan0~19_cout ));
// synopsys translate_off
defparam \LessThan0~19 .lut_mask = 16'h004D;
defparam \LessThan0~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N20
cycloneive_lcell_comb \LessThan0~21 (
// Equation(s):
// \LessThan0~21_cout  = CARRY((\rdat1[10]~31_combout  & (\port_b~65_combout  & !\LessThan0~19_cout )) # (!\rdat1[10]~31_combout  & ((\port_b~65_combout ) # (!\LessThan0~19_cout ))))

	.dataa(rdat1_10),
	.datab(port_b55),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~19_cout ),
	.combout(),
	.cout(\LessThan0~21_cout ));
// synopsys translate_off
defparam \LessThan0~21 .lut_mask = 16'h004D;
defparam \LessThan0~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N22
cycloneive_lcell_comb \LessThan0~23 (
// Equation(s):
// \LessThan0~23_cout  = CARRY((\rdat1[11]~29_combout  & ((!\LessThan0~21_cout ) # (!\port_b~67_combout ))) # (!\rdat1[11]~29_combout  & (!\port_b~67_combout  & !\LessThan0~21_cout )))

	.dataa(rdat1_11),
	.datab(port_b57),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~21_cout ),
	.combout(),
	.cout(\LessThan0~23_cout ));
// synopsys translate_off
defparam \LessThan0~23 .lut_mask = 16'h002B;
defparam \LessThan0~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N24
cycloneive_lcell_comb \LessThan0~25 (
// Equation(s):
// \LessThan0~25_cout  = CARRY((\port_b~72_combout  & ((!\LessThan0~23_cout ) # (!\rdat1[12]~27_combout ))) # (!\port_b~72_combout  & (!\rdat1[12]~27_combout  & !\LessThan0~23_cout )))

	.dataa(port_b62),
	.datab(rdat1_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~23_cout ),
	.combout(),
	.cout(\LessThan0~25_cout ));
// synopsys translate_off
defparam \LessThan0~25 .lut_mask = 16'h002B;
defparam \LessThan0~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N26
cycloneive_lcell_comb \LessThan0~27 (
// Equation(s):
// \LessThan0~27_cout  = CARRY((\rdat1[13]~25_combout  & ((!\LessThan0~25_cout ) # (!\port_b~70_combout ))) # (!\rdat1[13]~25_combout  & (!\port_b~70_combout  & !\LessThan0~25_cout )))

	.dataa(rdat1_13),
	.datab(port_b60),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~25_cout ),
	.combout(),
	.cout(\LessThan0~27_cout ));
// synopsys translate_off
defparam \LessThan0~27 .lut_mask = 16'h002B;
defparam \LessThan0~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N28
cycloneive_lcell_comb \LessThan0~29 (
// Equation(s):
// \LessThan0~29_cout  = CARRY((\rdat1[14]~23_combout  & (\port_b~71_combout  & !\LessThan0~27_cout )) # (!\rdat1[14]~23_combout  & ((\port_b~71_combout ) # (!\LessThan0~27_cout ))))

	.dataa(rdat1_14),
	.datab(port_b61),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~27_cout ),
	.combout(),
	.cout(\LessThan0~29_cout ));
// synopsys translate_off
defparam \LessThan0~29 .lut_mask = 16'h004D;
defparam \LessThan0~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N30
cycloneive_lcell_comb \LessThan0~31 (
// Equation(s):
// \LessThan0~31_cout  = CARRY((\rdat1[15]~21_combout  & ((!\LessThan0~29_cout ) # (!\port_b~63_combout ))) # (!\rdat1[15]~21_combout  & (!\port_b~63_combout  & !\LessThan0~29_cout )))

	.dataa(rdat1_15),
	.datab(port_b53),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~29_cout ),
	.combout(),
	.cout(\LessThan0~31_cout ));
// synopsys translate_off
defparam \LessThan0~31 .lut_mask = 16'h002B;
defparam \LessThan0~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N0
cycloneive_lcell_comb \LessThan0~33 (
// Equation(s):
// \LessThan0~33_cout  = CARRY((\rdat1[16]~19_combout  & (\port_b~22_combout  & !\LessThan0~31_cout )) # (!\rdat1[16]~19_combout  & ((\port_b~22_combout ) # (!\LessThan0~31_cout ))))

	.dataa(rdat1_16),
	.datab(port_b12),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~31_cout ),
	.combout(),
	.cout(\LessThan0~33_cout ));
// synopsys translate_off
defparam \LessThan0~33 .lut_mask = 16'h004D;
defparam \LessThan0~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N2
cycloneive_lcell_comb \LessThan0~35 (
// Equation(s):
// \LessThan0~35_cout  = CARRY((\rdat1[17]~63_combout  & ((!\LessThan0~33_cout ) # (!\port_b~24_combout ))) # (!\rdat1[17]~63_combout  & (!\port_b~24_combout  & !\LessThan0~33_cout )))

	.dataa(rdat1_17),
	.datab(port_b14),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~33_cout ),
	.combout(),
	.cout(\LessThan0~35_cout ));
// synopsys translate_off
defparam \LessThan0~35 .lut_mask = 16'h002B;
defparam \LessThan0~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N4
cycloneive_lcell_comb \LessThan0~37 (
// Equation(s):
// \LessThan0~37_cout  = CARRY((\rdat1[18]~59_combout  & (\port_b~26_combout  & !\LessThan0~35_cout )) # (!\rdat1[18]~59_combout  & ((\port_b~26_combout ) # (!\LessThan0~35_cout ))))

	.dataa(rdat1_18),
	.datab(port_b16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~35_cout ),
	.combout(),
	.cout(\LessThan0~37_cout ));
// synopsys translate_off
defparam \LessThan0~37 .lut_mask = 16'h004D;
defparam \LessThan0~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N6
cycloneive_lcell_comb \LessThan0~39 (
// Equation(s):
// \LessThan0~39_cout  = CARRY((\rdat1[19]~61_combout  & ((!\LessThan0~37_cout ) # (!\port_b~28_combout ))) # (!\rdat1[19]~61_combout  & (!\port_b~28_combout  & !\LessThan0~37_cout )))

	.dataa(rdat1_19),
	.datab(port_b18),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~37_cout ),
	.combout(),
	.cout(\LessThan0~39_cout ));
// synopsys translate_off
defparam \LessThan0~39 .lut_mask = 16'h002B;
defparam \LessThan0~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N8
cycloneive_lcell_comb \LessThan0~41 (
// Equation(s):
// \LessThan0~41_cout  = CARRY((\rdat1[20]~57_combout  & (\port_b~30_combout  & !\LessThan0~39_cout )) # (!\rdat1[20]~57_combout  & ((\port_b~30_combout ) # (!\LessThan0~39_cout ))))

	.dataa(rdat1_20),
	.datab(port_b20),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~39_cout ),
	.combout(),
	.cout(\LessThan0~41_cout ));
// synopsys translate_off
defparam \LessThan0~41 .lut_mask = 16'h004D;
defparam \LessThan0~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N10
cycloneive_lcell_comb \LessThan0~43 (
// Equation(s):
// \LessThan0~43_cout  = CARRY((\port_b~32_combout  & (\rdat1[21]~55_combout  & !\LessThan0~41_cout )) # (!\port_b~32_combout  & ((\rdat1[21]~55_combout ) # (!\LessThan0~41_cout ))))

	.dataa(port_b22),
	.datab(rdat1_21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~41_cout ),
	.combout(),
	.cout(\LessThan0~43_cout ));
// synopsys translate_off
defparam \LessThan0~43 .lut_mask = 16'h004D;
defparam \LessThan0~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N12
cycloneive_lcell_comb \LessThan0~45 (
// Equation(s):
// \LessThan0~45_cout  = CARRY((\rdat1[22]~51_combout  & (\port_b~34_combout  & !\LessThan0~43_cout )) # (!\rdat1[22]~51_combout  & ((\port_b~34_combout ) # (!\LessThan0~43_cout ))))

	.dataa(rdat1_22),
	.datab(port_b24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~43_cout ),
	.combout(),
	.cout(\LessThan0~45_cout ));
// synopsys translate_off
defparam \LessThan0~45 .lut_mask = 16'h004D;
defparam \LessThan0~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N14
cycloneive_lcell_comb \LessThan0~47 (
// Equation(s):
// \LessThan0~47_cout  = CARRY((\rdat1[23]~53_combout  & ((!\LessThan0~45_cout ) # (!\port_b~36_combout ))) # (!\rdat1[23]~53_combout  & (!\port_b~36_combout  & !\LessThan0~45_cout )))

	.dataa(rdat1_23),
	.datab(port_b26),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~45_cout ),
	.combout(),
	.cout(\LessThan0~47_cout ));
// synopsys translate_off
defparam \LessThan0~47 .lut_mask = 16'h002B;
defparam \LessThan0~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N16
cycloneive_lcell_comb \LessThan0~49 (
// Equation(s):
// \LessThan0~49_cout  = CARRY((\port_b~38_combout  & ((!\LessThan0~47_cout ) # (!\rdat1[24]~49_combout ))) # (!\port_b~38_combout  & (!\rdat1[24]~49_combout  & !\LessThan0~47_cout )))

	.dataa(port_b28),
	.datab(rdat1_24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~47_cout ),
	.combout(),
	.cout(\LessThan0~49_cout ));
// synopsys translate_off
defparam \LessThan0~49 .lut_mask = 16'h002B;
defparam \LessThan0~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N18
cycloneive_lcell_comb \LessThan0~51 (
// Equation(s):
// \LessThan0~51_cout  = CARRY((\port_b~40_combout  & (\rdat1[25]~47_combout  & !\LessThan0~49_cout )) # (!\port_b~40_combout  & ((\rdat1[25]~47_combout ) # (!\LessThan0~49_cout ))))

	.dataa(port_b30),
	.datab(rdat1_25),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~49_cout ),
	.combout(),
	.cout(\LessThan0~51_cout ));
// synopsys translate_off
defparam \LessThan0~51 .lut_mask = 16'h004D;
defparam \LessThan0~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N20
cycloneive_lcell_comb \LessThan0~53 (
// Equation(s):
// \LessThan0~53_cout  = CARRY((\rdat1[26]~43_combout  & (\port_b~42_combout  & !\LessThan0~51_cout )) # (!\rdat1[26]~43_combout  & ((\port_b~42_combout ) # (!\LessThan0~51_cout ))))

	.dataa(rdat1_26),
	.datab(port_b32),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~51_cout ),
	.combout(),
	.cout(\LessThan0~53_cout ));
// synopsys translate_off
defparam \LessThan0~53 .lut_mask = 16'h004D;
defparam \LessThan0~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N22
cycloneive_lcell_comb \LessThan0~55 (
// Equation(s):
// \LessThan0~55_cout  = CARRY((\port_b~52_combout  & (\rdat1[27]~45_combout  & !\LessThan0~53_cout )) # (!\port_b~52_combout  & ((\rdat1[27]~45_combout ) # (!\LessThan0~53_cout ))))

	.dataa(port_b42),
	.datab(rdat1_27),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~53_cout ),
	.combout(),
	.cout(\LessThan0~55_cout ));
// synopsys translate_off
defparam \LessThan0~55 .lut_mask = 16'h004D;
defparam \LessThan0~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N24
cycloneive_lcell_comb \LessThan0~57 (
// Equation(s):
// \LessThan0~57_cout  = CARRY((\port_b~54_combout  & ((!\LessThan0~55_cout ) # (!\rdat1[28]~41_combout ))) # (!\port_b~54_combout  & (!\rdat1[28]~41_combout  & !\LessThan0~55_cout )))

	.dataa(port_b44),
	.datab(rdat1_28),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~55_cout ),
	.combout(),
	.cout(\LessThan0~57_cout ));
// synopsys translate_off
defparam \LessThan0~57 .lut_mask = 16'h002B;
defparam \LessThan0~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N26
cycloneive_lcell_comb \LessThan0~59 (
// Equation(s):
// \LessThan0~59_cout  = CARRY((\rdat1[29]~37_combout  & ((!\LessThan0~57_cout ) # (!\port_b~56_combout ))) # (!\rdat1[29]~37_combout  & (!\port_b~56_combout  & !\LessThan0~57_cout )))

	.dataa(rdat1_29),
	.datab(port_b46),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~57_cout ),
	.combout(),
	.cout(\LessThan0~59_cout ));
// synopsys translate_off
defparam \LessThan0~59 .lut_mask = 16'h002B;
defparam \LessThan0~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N28
cycloneive_lcell_comb \LessThan0~61 (
// Equation(s):
// \LessThan0~61_cout  = CARRY((\port_b~58_combout  & ((!\LessThan0~59_cout ) # (!\rdat1[30]~39_combout ))) # (!\port_b~58_combout  & (!\rdat1[30]~39_combout  & !\LessThan0~59_cout )))

	.dataa(port_b48),
	.datab(rdat1_30),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~59_cout ),
	.combout(),
	.cout(\LessThan0~61_cout ));
// synopsys translate_off
defparam \LessThan0~61 .lut_mask = 16'h002B;
defparam \LessThan0~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N30
cycloneive_lcell_comb \LessThan0~62 (
// Equation(s):
// \LessThan0~62_combout  = (\rdat1[31]~35_combout  & ((\LessThan0~61_cout ) # (!\port_b~20_combout ))) # (!\rdat1[31]~35_combout  & (\LessThan0~61_cout  & !\port_b~20_combout ))

	.dataa(rdat1_311),
	.datab(gnd),
	.datac(gnd),
	.datad(port_b10),
	.cin(\LessThan0~61_cout ),
	.combout(\LessThan0~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan0~62 .lut_mask = 16'hA0FA;
defparam \LessThan0~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N16
cycloneive_lcell_comb \ShiftLeft0~3 (
// Equation(s):
// \ShiftLeft0~3_combout  = (\port_b~28_combout ) # ((\port_b~30_combout ) # ((\port_b~34_combout ) # (\port_b~32_combout )))

	.dataa(port_b18),
	.datab(port_b20),
	.datac(port_b24),
	.datad(port_b22),
	.cin(gnd),
	.combout(\ShiftLeft0~3_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~3 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N20
cycloneive_lcell_comb \ShiftLeft0~6 (
// Equation(s):
// \ShiftLeft0~6_combout  = (\port_b~54_combout ) # ((\port_b~52_combout ) # ((\port_b~56_combout ) # (\port_b~58_combout )))

	.dataa(port_b44),
	.datab(port_b42),
	.datac(port_b46),
	.datad(port_b48),
	.cin(gnd),
	.combout(\ShiftLeft0~6_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~6 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N24
cycloneive_lcell_comb \ShiftLeft0~14 (
// Equation(s):
// \ShiftLeft0~14_combout  = (\ShiftLeft0~12_combout  & (!\ShiftLeft0~13_combout  & !\port_b~14_combout ))

	.dataa(\ShiftLeft0~12_combout ),
	.datab(gnd),
	.datac(\ShiftLeft0~13_combout ),
	.datad(port_b7),
	.cin(gnd),
	.combout(\ShiftLeft0~14_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~14 .lut_mask = 16'h000A;
defparam \ShiftLeft0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N30
cycloneive_lcell_comb \ShiftRight0~32 (
// Equation(s):
// \ShiftRight0~32_combout  = (!\port_b~7_combout  & ((\port_b~4_combout  & (\rdat1[20]~57_combout )) # (!\port_b~4_combout  & ((\rdat1[18]~59_combout )))))

	.dataa(port_b2),
	.datab(rdat1_20),
	.datac(rdat1_18),
	.datad(port_b4),
	.cin(gnd),
	.combout(\ShiftRight0~32_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~32 .lut_mask = 16'h00D8;
defparam \ShiftRight0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N12
cycloneive_lcell_comb \ShiftRight0~34 (
// Equation(s):
// \ShiftRight0~34_combout  = (\ShiftRight0~32_combout ) # ((\port_b~7_combout  & \ShiftRight0~33_combout ))

	.dataa(port_b4),
	.datab(gnd),
	.datac(\ShiftRight0~33_combout ),
	.datad(\ShiftRight0~32_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~34_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~34 .lut_mask = 16'hFFA0;
defparam \ShiftRight0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N22
cycloneive_lcell_comb \myif.out[6]~18 (
// Equation(s):
// \myif.out[6]~18_combout  = (\myif.out[5]~16_combout  & (\myif.out[5]~17_combout )) # (!\myif.out[5]~16_combout  & ((\myif.out[5]~17_combout  & (\ShiftRight0~41_combout )) # (!\myif.out[5]~17_combout  & ((\ShiftRight0~44_combout )))))

	.dataa(\myif.out[5]~16_combout ),
	.datab(\myif.out[5]~17_combout ),
	.datac(\ShiftRight0~41_combout ),
	.datad(\ShiftRight0~44_combout ),
	.cin(gnd),
	.combout(\myif.out[6]~18_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[6]~18 .lut_mask = 16'hD9C8;
defparam \myif.out[6]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N10
cycloneive_lcell_comb \ShiftRight0~57 (
// Equation(s):
// \ShiftRight0~57_combout  = (\port_b~4_combout  & (\ShiftRight0~36_combout )) # (!\port_b~4_combout  & ((\ShiftRight0~39_combout )))

	.dataa(gnd),
	.datab(port_b2),
	.datac(\ShiftRight0~36_combout ),
	.datad(\ShiftRight0~39_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~57_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~57 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N26
cycloneive_lcell_comb \ShiftRight0~66 (
// Equation(s):
// \ShiftRight0~66_combout  = (!\port_b~4_combout  & ((\port_b~7_combout  & ((\rdat1[29]~37_combout ))) # (!\port_b~7_combout  & (\rdat1[28]~41_combout ))))

	.dataa(port_b4),
	.datab(port_b2),
	.datac(rdat1_28),
	.datad(rdat1_29),
	.cin(gnd),
	.combout(\ShiftRight0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~66 .lut_mask = 16'h3210;
defparam \ShiftRight0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N10
cycloneive_lcell_comb \ShiftLeft0~31 (
// Equation(s):
// \ShiftLeft0~31_combout  = (!\port_b~7_combout  & ((\port_b~4_combout  & (\rdat1[18]~59_combout )) # (!\port_b~4_combout  & ((\rdat1[20]~57_combout )))))

	.dataa(rdat1_18),
	.datab(port_b4),
	.datac(port_b2),
	.datad(rdat1_20),
	.cin(gnd),
	.combout(\ShiftLeft0~31_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~31 .lut_mask = 16'h2320;
defparam \ShiftLeft0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N6
cycloneive_lcell_comb \out~13 (
// Equation(s):
// \out~13_combout  = (\rdat1[24]~49_combout  & ((\port_b~37_combout ) # ((\port_b~0_combout  & fuifrtReplace_24))))

	.dataa(port_b),
	.datab(port_b27),
	.datac(fuifrtReplace_24),
	.datad(rdat1_24),
	.cin(gnd),
	.combout(\out~13_combout ),
	.cout());
// synopsys translate_off
defparam \out~13 .lut_mask = 16'hEC00;
defparam \out~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N2
cycloneive_lcell_comb \ShiftLeft0~62 (
// Equation(s):
// \ShiftLeft0~62_combout  = (\port_b~7_combout  & ((\port_b~4_combout  & ((\rdat1[18]~59_combout ))) # (!\port_b~4_combout  & (\rdat1[20]~57_combout ))))

	.dataa(port_b2),
	.datab(rdat1_20),
	.datac(port_b4),
	.datad(rdat1_18),
	.cin(gnd),
	.combout(\ShiftLeft0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~62 .lut_mask = 16'hE040;
defparam \ShiftLeft0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N12
cycloneive_lcell_comb \ShiftLeft0~63 (
// Equation(s):
// \ShiftLeft0~63_combout  = (\ShiftLeft0~62_combout ) # ((!\port_b~7_combout  & \ShiftLeft0~41_combout ))

	.dataa(gnd),
	.datab(port_b4),
	.datac(\ShiftLeft0~41_combout ),
	.datad(\ShiftLeft0~62_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~63 .lut_mask = 16'hFF30;
defparam \ShiftLeft0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N22
cycloneive_lcell_comb \ShiftLeft0~79 (
// Equation(s):
// \ShiftLeft0~79_combout  = (\port_b~4_combout  & ((\port_b~7_combout  & (\rdat1[24]~49_combout )) # (!\port_b~7_combout  & ((\rdat1[25]~47_combout )))))

	.dataa(rdat1_24),
	.datab(port_b4),
	.datac(rdat1_25),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftLeft0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~79 .lut_mask = 16'hB800;
defparam \ShiftLeft0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N10
cycloneive_lcell_comb \ShiftLeft0~80 (
// Equation(s):
// \ShiftLeft0~80_combout  = (\port_b~7_combout  & (\rdat1[26]~43_combout )) # (!\port_b~7_combout  & ((\rdat1[27]~45_combout )))

	.dataa(rdat1_26),
	.datab(port_b4),
	.datac(rdat1_27),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~80 .lut_mask = 16'hB8B8;
defparam \ShiftLeft0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N30
cycloneive_lcell_comb \ShiftLeft0~81 (
// Equation(s):
// \ShiftLeft0~81_combout  = (\ShiftLeft0~79_combout ) # ((!\port_b~4_combout  & \ShiftLeft0~80_combout ))

	.dataa(port_b2),
	.datab(\ShiftLeft0~79_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~80_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~81 .lut_mask = 16'hDDCC;
defparam \ShiftLeft0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N24
cycloneive_lcell_comb \myif.out[7]~73 (
// Equation(s):
// \myif.out[7]~73_combout  = (!\port_b~0_combout ) # (!fuifrtReplace_7)

	.dataa(gnd),
	.datab(gnd),
	.datac(fuifrtReplace_7),
	.datad(port_b),
	.cin(gnd),
	.combout(\myif.out[7]~73_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[7]~73 .lut_mask = 16'h0FFF;
defparam \myif.out[7]~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N18
cycloneive_lcell_comb \myif.out[7]~74 (
// Equation(s):
// \myif.out[7]~74_combout  = (\rdat1[7]~13_combout  $ (((\port_b~47_combout ) # (!\myif.out[7]~73_combout )))) # (!idex_ifaluop_o_1)

	.dataa(port_b37),
	.datab(idex_ifaluop_o_1),
	.datac(rdat1_7),
	.datad(\myif.out[7]~73_combout ),
	.cin(gnd),
	.combout(\myif.out[7]~74_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[7]~74 .lut_mask = 16'h7B3F;
defparam \myif.out[7]~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N28
cycloneive_lcell_comb \ShiftRight0~91 (
// Equation(s):
// \ShiftRight0~91_combout  = (\ShiftRight0~18_combout  & \ShiftRight0~112_combout )

	.dataa(\ShiftRight0~18_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\ShiftRight0~112_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~91_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~91 .lut_mask = 16'hAA00;
defparam \ShiftRight0~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N8
cycloneive_lcell_comb \ShiftRight0~95 (
// Equation(s):
// \ShiftRight0~95_combout  = (\ShiftRight0~112_combout  & ((\ShiftRight0~66_combout ) # ((\port_b~4_combout  & \ShiftRight0~52_combout ))))

	.dataa(\ShiftRight0~66_combout ),
	.datab(port_b2),
	.datac(\ShiftRight0~52_combout ),
	.datad(\ShiftRight0~112_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~95_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~95 .lut_mask = 16'hEA00;
defparam \ShiftRight0~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N10
cycloneive_lcell_comb \ShiftLeft0~95 (
// Equation(s):
// \ShiftLeft0~95_combout  = (\port_b~10_combout  & (\ShiftLeft0~21_combout )) # (!\port_b~10_combout  & ((\ShiftLeft0~23_combout )))

	.dataa(port_b6),
	.datab(\ShiftLeft0~21_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~23_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~95_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~95 .lut_mask = 16'hDD88;
defparam \ShiftLeft0~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N6
cycloneive_lcell_comb \out~44 (
// Equation(s):
// \out~44_combout  = (\rdat1[15]~21_combout  & ((\port_b~62_combout ) # ((\port_b~0_combout  & fuifrtReplace_15))))

	.dataa(port_b),
	.datab(port_b52),
	.datac(rdat1_15),
	.datad(fuifrtReplace_15),
	.cin(gnd),
	.combout(\out~44_combout ),
	.cout());
// synopsys translate_off
defparam \out~44 .lut_mask = 16'hE0C0;
defparam \out~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N20
cycloneive_lcell_comb \out~49 (
// Equation(s):
// \out~49_combout  = \rdat1[11]~29_combout  $ (((\port_b~66_combout ) # ((\port_b~0_combout  & fuifrtReplace_11))))

	.dataa(rdat1_11),
	.datab(port_b56),
	.datac(port_b),
	.datad(fuifrtReplace_11),
	.cin(gnd),
	.combout(\out~49_combout ),
	.cout());
// synopsys translate_off
defparam \out~49 .lut_mask = 16'h5666;
defparam \out~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N22
cycloneive_lcell_comb \myif.out[17]~166 (
// Equation(s):
// \myif.out[17]~166_combout  = (\rdat1[17]~63_combout  & (idex_ifaluop_o_1 $ (((!idex_ifaluop_o_2))))) # (!\rdat1[17]~63_combout  & ((idex_ifaluop_o_1 $ (!idex_ifaluop_o_2)) # (!\myif.out[17]~165_combout )))

	.dataa(rdat1_17),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[17]~165_combout ),
	.datad(idex_ifaluop_o_2),
	.cin(gnd),
	.combout(\myif.out[17]~166_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[17]~166 .lut_mask = 16'hCD37;
defparam \myif.out[17]~166 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N6
cycloneive_lcell_comb \out~57 (
// Equation(s):
// \out~57_combout  = (\rdat1[18]~59_combout  & ((\port_b~25_combout ) # ((fuifrtReplace_18 & \port_b~0_combout ))))

	.dataa(port_b15),
	.datab(fuifrtReplace_18),
	.datac(rdat1_18),
	.datad(port_b),
	.cin(gnd),
	.combout(\out~57_combout ),
	.cout());
// synopsys translate_off
defparam \out~57 .lut_mask = 16'hE0A0;
defparam \out~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N30
cycloneive_lcell_comb \myif.out[19]~188 (
// Equation(s):
// \myif.out[19]~188_combout  = (\myif.out[19]~187_combout  & (idex_ifaluop_o_2 $ ((!idex_ifaluop_o_1)))) # (!\myif.out[19]~187_combout  & ((idex_ifaluop_o_2 $ (!idex_ifaluop_o_1)) # (!\rdat1[19]~61_combout )))

	.dataa(idex_ifaluop_o_2),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[19]~187_combout ),
	.datad(rdat1_19),
	.cin(gnd),
	.combout(\myif.out[19]~188_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[19]~188 .lut_mask = 16'h999F;
defparam \myif.out[19]~188 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N12
cycloneive_lcell_comb \myif.out[30]~197 (
// Equation(s):
// \myif.out[30]~197_combout  = (\myif.out[13]~23_combout  & ((idex_ifaluop_o_2 & ((\out~60_combout ))) # (!idex_ifaluop_o_2 & (\ShiftRight0~94_combout )))) # (!\myif.out[13]~23_combout  & (idex_ifaluop_o_2))

	.dataa(\myif.out[13]~23_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\ShiftRight0~94_combout ),
	.datad(\out~60_combout ),
	.cin(gnd),
	.combout(\myif.out[30]~197_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[30]~197 .lut_mask = 16'hEC64;
defparam \myif.out[30]~197 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N10
cycloneive_lcell_comb \out~61 (
// Equation(s):
// \out~61_combout  = (\rdat1[30]~39_combout  & ((\port_b~57_combout ) # ((\port_b~0_combout  & fuifrtReplace_30))))

	.dataa(port_b),
	.datab(rdat1_30),
	.datac(port_b47),
	.datad(fuifrtReplace_30),
	.cin(gnd),
	.combout(\out~61_combout ),
	.cout());
// synopsys translate_off
defparam \out~61 .lut_mask = 16'hC8C0;
defparam \out~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N6
cycloneive_lcell_comb \myif.out[21]~212 (
// Equation(s):
// \myif.out[21]~212_combout  = (\rdat1[21]~55_combout  & (idex_ifaluop_o_1 $ ((!idex_ifaluop_o_2)))) # (!\rdat1[21]~55_combout  & ((idex_ifaluop_o_1 $ (!idex_ifaluop_o_2)) # (!\myif.out[21]~211_combout )))

	.dataa(idex_ifaluop_o_1),
	.datab(idex_ifaluop_o_2),
	.datac(rdat1_21),
	.datad(\myif.out[21]~211_combout ),
	.cin(gnd),
	.combout(\myif.out[21]~212_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[21]~212 .lut_mask = 16'h999F;
defparam \myif.out[21]~212 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N22
cycloneive_lcell_comb \myif.negative~3 (
// Equation(s):
// \myif.negative~3_combout  = (\ShiftLeft0~13_combout  & (((\ShiftLeft0~107_combout ) # (\myif.negative~0_combout )))) # (!\ShiftLeft0~13_combout  & (\rdat1[31]~35_combout  & ((!\myif.negative~0_combout ))))

	.dataa(\ShiftLeft0~13_combout ),
	.datab(rdat1_311),
	.datac(\ShiftLeft0~107_combout ),
	.datad(\myif.negative~0_combout ),
	.cin(gnd),
	.combout(\myif.negative~3_combout ),
	.cout());
// synopsys translate_off
defparam \myif.negative~3 .lut_mask = 16'hAAE4;
defparam \myif.negative~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N12
cycloneive_lcell_comb \myif.negative~4 (
// Equation(s):
// \myif.negative~4_combout  = (\myif.negative~0_combout  & ((\myif.negative~3_combout  & (\ShiftLeft0~81_combout )) # (!\myif.negative~3_combout  & ((\rdat1[30]~39_combout ))))) # (!\myif.negative~0_combout  & (((\myif.negative~3_combout ))))

	.dataa(\ShiftLeft0~81_combout ),
	.datab(\myif.negative~0_combout ),
	.datac(\myif.negative~3_combout ),
	.datad(rdat1_30),
	.cin(gnd),
	.combout(\myif.negative~4_combout ),
	.cout());
// synopsys translate_off
defparam \myif.negative~4 .lut_mask = 16'hBCB0;
defparam \myif.negative~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N28
cycloneive_lcell_comb \out~65 (
// Equation(s):
// \out~65_combout  = (\rdat1[31]~35_combout  & ((\port_b~19_combout ) # ((\port_b~0_combout  & fuifrtReplace_31))))

	.dataa(port_b),
	.datab(port_b9),
	.datac(rdat1_311),
	.datad(fuifrtReplace_31),
	.cin(gnd),
	.combout(\out~65_combout ),
	.cout());
// synopsys translate_off
defparam \out~65 .lut_mask = 16'hE0C0;
defparam \out~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N16
cycloneive_lcell_comb \out~71 (
// Equation(s):
// \out~71_combout  = (\rdat1[20]~57_combout  & ((\port_b~29_combout ) # ((\port_b~0_combout  & fuifrtReplace_20))))

	.dataa(port_b19),
	.datab(port_b),
	.datac(rdat1_20),
	.datad(fuifrtReplace_20),
	.cin(gnd),
	.combout(\out~71_combout ),
	.cout());
// synopsys translate_off
defparam \out~71 .lut_mask = 16'hE0A0;
defparam \out~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N30
cycloneive_lcell_comb \ShiftRight0~106 (
// Equation(s):
// \ShiftRight0~106_combout  = (!\port_b~4_combout  & ((\port_b~7_combout  & ((\rdat1[1]~1_combout ))) # (!\port_b~7_combout  & (\rdat1[0]~3_combout ))))

	.dataa(port_b2),
	.datab(port_b4),
	.datac(rdat1_0),
	.datad(rdat1_1),
	.cin(gnd),
	.combout(\ShiftRight0~106_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~106 .lut_mask = 16'h5410;
defparam \ShiftRight0~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N10
cycloneive_lcell_comb \ShiftRight0~108 (
// Equation(s):
// \ShiftRight0~108_combout  = (!\port_b~10_combout  & ((\ShiftRight0~106_combout ) # ((\port_b~4_combout  & \ShiftRight0~107_combout ))))

	.dataa(port_b2),
	.datab(port_b6),
	.datac(\ShiftRight0~106_combout ),
	.datad(\ShiftRight0~107_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~108_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~108 .lut_mask = 16'h3230;
defparam \ShiftRight0~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N4
cycloneive_lcell_comb \ShiftRight0~109 (
// Equation(s):
// \ShiftRight0~109_combout  = (!\port_b~14_combout  & ((\ShiftRight0~108_combout ) # ((\ShiftRight0~60_combout  & \port_b~10_combout ))))

	.dataa(\ShiftRight0~60_combout ),
	.datab(port_b7),
	.datac(port_b6),
	.datad(\ShiftRight0~108_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~109_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~109 .lut_mask = 16'h3320;
defparam \ShiftRight0~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N22
cycloneive_lcell_comb \ShiftRight0~110 (
// Equation(s):
// \ShiftRight0~110_combout  = (\ShiftRight0~109_combout ) # ((\port_b~14_combout  & \ShiftRight0~92_combout ))

	.dataa(gnd),
	.datab(port_b7),
	.datac(\ShiftRight0~109_combout ),
	.datad(\ShiftRight0~92_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~110_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~110 .lut_mask = 16'hFCF0;
defparam \ShiftRight0~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N4
cycloneive_lcell_comb \myif.out[0]~233 (
// Equation(s):
// \myif.out[0]~233_combout  = (\rdat1[0]~3_combout  & ((\port_b~6_combout ) # ((fuifrtReplace_0 & \port_b~0_combout ))))

	.dataa(fuifrtReplace_0),
	.datab(port_b),
	.datac(port_b3),
	.datad(rdat1_0),
	.cin(gnd),
	.combout(\myif.out[0]~233_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[0]~233 .lut_mask = 16'hF800;
defparam \myif.out[0]~233 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N8
cycloneive_lcell_comb \myif.out[0]~234 (
// Equation(s):
// \myif.out[0]~234_combout  = (idex_ifaluop_o_2 & ((idex_ifaluop_o_0) # ((\myif.out[0]~233_combout )))) # (!idex_ifaluop_o_2 & (!idex_ifaluop_o_0 & ((!\port_b~17_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(idex_ifaluop_o_0),
	.datac(\myif.out[0]~233_combout ),
	.datad(port_b8),
	.cin(gnd),
	.combout(\myif.out[0]~234_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[0]~234 .lut_mask = 16'hA8B9;
defparam \myif.out[0]~234 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N6
cycloneive_lcell_comb \out~79 (
// Equation(s):
// \out~79_combout  = (\port_b~17_combout  & ((\rdat1[4]~6_combout ) # ((always03 & \mem_data~10_combout ))))

	.dataa(always0),
	.datab(rdat1_4),
	.datac(mem_data),
	.datad(port_b8),
	.cin(gnd),
	.combout(\out~79_combout ),
	.cout());
// synopsys translate_off
defparam \out~79 .lut_mask = 16'hEC00;
defparam \out~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N6
cycloneive_lcell_comb \myif.out[1]~15 (
// Equation(s):
// myifout_1 = (!idex_ifaluop_o_3 & ((idex_ifaluop_o_0 & ((\myif.out[1]~9_combout ))) # (!idex_ifaluop_o_0 & (\myif.out[1]~14_combout ))))

	.dataa(idex_ifaluop_o_3),
	.datab(idex_ifaluop_o_0),
	.datac(\myif.out[1]~14_combout ),
	.datad(\myif.out[1]~9_combout ),
	.cin(gnd),
	.combout(myifout_1),
	.cout());
// synopsys translate_off
defparam \myif.out[1]~15 .lut_mask = 16'h5410;
defparam \myif.out[1]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N4
cycloneive_lcell_comb \myif.out[6]~26 (
// Equation(s):
// myifout_6 = (!idex_ifaluop_o_3 & ((idex_ifaluop_o_0 & ((\myif.out[6]~22_combout ))) # (!idex_ifaluop_o_0 & (\myif.out[6]~25_combout ))))

	.dataa(idex_ifaluop_o_3),
	.datab(idex_ifaluop_o_0),
	.datac(\myif.out[6]~25_combout ),
	.datad(\myif.out[6]~22_combout ),
	.cin(gnd),
	.combout(myifout_6),
	.cout());
// synopsys translate_off
defparam \myif.out[6]~26 .lut_mask = 16'h5410;
defparam \myif.out[6]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N14
cycloneive_lcell_comb \myif.out[4]~33 (
// Equation(s):
// myifout_4 = (!idex_ifaluop_o_3 & ((idex_ifaluop_o_0 & (\myif.out[4]~30_combout )) # (!idex_ifaluop_o_0 & ((\myif.out[4]~32_combout )))))

	.dataa(idex_ifaluop_o_3),
	.datab(idex_ifaluop_o_0),
	.datac(\myif.out[4]~30_combout ),
	.datad(\myif.out[4]~32_combout ),
	.cin(gnd),
	.combout(myifout_4),
	.cout());
// synopsys translate_off
defparam \myif.out[4]~33 .lut_mask = 16'h5140;
defparam \myif.out[4]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N12
cycloneive_lcell_comb \myif.out[24]~40 (
// Equation(s):
// myifout_24 = (!idex_ifaluop_o_3 & ((idex_ifaluop_o_0 & ((\myif.out[24]~35_combout ))) # (!idex_ifaluop_o_0 & (\myif.out[24]~39_combout ))))

	.dataa(idex_ifaluop_o_0),
	.datab(idex_ifaluop_o_3),
	.datac(\myif.out[24]~39_combout ),
	.datad(\myif.out[24]~35_combout ),
	.cin(gnd),
	.combout(myifout_24),
	.cout());
// synopsys translate_off
defparam \myif.out[24]~40 .lut_mask = 16'h3210;
defparam \myif.out[24]~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N30
cycloneive_lcell_comb \myif.out[26]~47 (
// Equation(s):
// myifout_26 = (!idex_ifaluop_o_3 & ((idex_ifaluop_o_0 & (\myif.out[26]~42_combout )) # (!idex_ifaluop_o_0 & ((\myif.out[26]~46_combout )))))

	.dataa(idex_ifaluop_o_0),
	.datab(idex_ifaluop_o_3),
	.datac(\myif.out[26]~42_combout ),
	.datad(\myif.out[26]~46_combout ),
	.cin(gnd),
	.combout(myifout_26),
	.cout());
// synopsys translate_off
defparam \myif.out[26]~47 .lut_mask = 16'h3120;
defparam \myif.out[26]~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N2
cycloneive_lcell_comb \myif.out[25]~54 (
// Equation(s):
// myifout_25 = (!idex_ifaluop_o_3 & ((idex_ifaluop_o_0 & (\myif.out[25]~49_combout )) # (!idex_ifaluop_o_0 & ((\myif.out[25]~53_combout )))))

	.dataa(idex_ifaluop_o_0),
	.datab(idex_ifaluop_o_3),
	.datac(\myif.out[25]~49_combout ),
	.datad(\myif.out[25]~53_combout ),
	.cin(gnd),
	.combout(myifout_25),
	.cout());
// synopsys translate_off
defparam \myif.out[25]~54 .lut_mask = 16'h3120;
defparam \myif.out[25]~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N28
cycloneive_lcell_comb \myif.out[27]~61 (
// Equation(s):
// myifout_27 = (!idex_ifaluop_o_3 & ((idex_ifaluop_o_0 & ((\myif.out[27]~56_combout ))) # (!idex_ifaluop_o_0 & (\myif.out[27]~60_combout ))))

	.dataa(idex_ifaluop_o_0),
	.datab(idex_ifaluop_o_3),
	.datac(\myif.out[27]~60_combout ),
	.datad(\myif.out[27]~56_combout ),
	.cin(gnd),
	.combout(myifout_27),
	.cout());
// synopsys translate_off
defparam \myif.out[27]~61 .lut_mask = 16'h3210;
defparam \myif.out[27]~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N14
cycloneive_lcell_comb \myif.out[5]~68 (
// Equation(s):
// myifout_5 = (!idex_ifaluop_o_3 & ((idex_ifaluop_o_0 & ((\myif.out[5]~65_combout ))) # (!idex_ifaluop_o_0 & (\myif.out[5]~67_combout ))))

	.dataa(idex_ifaluop_o_0),
	.datab(\myif.out[5]~67_combout ),
	.datac(\myif.out[5]~65_combout ),
	.datad(idex_ifaluop_o_3),
	.cin(gnd),
	.combout(myifout_5),
	.cout());
// synopsys translate_off
defparam \myif.out[5]~68 .lut_mask = 16'h00E4;
defparam \myif.out[5]~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N24
cycloneive_lcell_comb \myif.out[7]~81 (
// Equation(s):
// myifout_7 = (!idex_ifaluop_o_3 & ((idex_ifaluop_o_0 & ((\myif.out[7]~72_combout ))) # (!idex_ifaluop_o_0 & (\myif.out[7]~80_combout ))))

	.dataa(\myif.out[7]~80_combout ),
	.datab(idex_ifaluop_o_0),
	.datac(idex_ifaluop_o_3),
	.datad(\myif.out[7]~72_combout ),
	.cin(gnd),
	.combout(myifout_7),
	.cout());
// synopsys translate_off
defparam \myif.out[7]~81 .lut_mask = 16'h0E02;
defparam \myif.out[7]~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N4
cycloneive_lcell_comb \myif.out[13]~92 (
// Equation(s):
// myifout_13 = (\myif.out[13]~87_combout  & ((\myif.out[13]~91_combout  & (!\out~27_combout )) # (!\myif.out[13]~91_combout  & ((\myif.out[13]~86_combout ))))) # (!\myif.out[13]~87_combout  & (((\myif.out[13]~91_combout ))))

	.dataa(\out~27_combout ),
	.datab(\myif.out[13]~87_combout ),
	.datac(\myif.out[13]~86_combout ),
	.datad(\myif.out[13]~91_combout ),
	.cin(gnd),
	.combout(myifout_13),
	.cout());
// synopsys translate_off
defparam \myif.out[13]~92 .lut_mask = 16'h77C0;
defparam \myif.out[13]~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N24
cycloneive_lcell_comb \myif.out[9]~98 (
// Equation(s):
// myifout_9 = (\myif.out[13]~88_combout  & ((\myif.out[9]~97_combout  & (!\out~30_combout )) # (!\myif.out[9]~97_combout  & ((\Add1~18_combout ))))) # (!\myif.out[13]~88_combout  & (((\myif.out[9]~97_combout ))))

	.dataa(\myif.out[13]~88_combout ),
	.datab(\out~30_combout ),
	.datac(\Add1~18_combout ),
	.datad(\myif.out[9]~97_combout ),
	.cin(gnd),
	.combout(myifout_9),
	.cout());
// synopsys translate_off
defparam \myif.out[9]~98 .lut_mask = 16'h77A0;
defparam \myif.out[9]~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N12
cycloneive_lcell_comb \myif.out[8]~104 (
// Equation(s):
// myifout_8 = (\myif.out[13]~87_combout  & ((\myif.out[8]~103_combout  & ((!\out~33_combout ))) # (!\myif.out[8]~103_combout  & (\myif.out[8]~100_combout )))) # (!\myif.out[13]~87_combout  & (((\myif.out[8]~103_combout ))))

	.dataa(\myif.out[8]~100_combout ),
	.datab(\myif.out[13]~87_combout ),
	.datac(\myif.out[8]~103_combout ),
	.datad(\out~33_combout ),
	.cin(gnd),
	.combout(myifout_8),
	.cout());
// synopsys translate_off
defparam \myif.out[8]~104 .lut_mask = 16'h38F8;
defparam \myif.out[8]~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N2
cycloneive_lcell_comb \myif.out[14]~110 (
// Equation(s):
// myifout_14 = (\myif.out[13]~88_combout  & ((\myif.out[14]~109_combout  & ((!\out~36_combout ))) # (!\myif.out[14]~109_combout  & (\Add1~28_combout )))) # (!\myif.out[13]~88_combout  & (((\myif.out[14]~109_combout ))))

	.dataa(\myif.out[13]~88_combout ),
	.datab(\Add1~28_combout ),
	.datac(\out~36_combout ),
	.datad(\myif.out[14]~109_combout ),
	.cin(gnd),
	.combout(myifout_14),
	.cout());
// synopsys translate_off
defparam \myif.out[14]~110 .lut_mask = 16'h5F88;
defparam \myif.out[14]~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N26
cycloneive_lcell_comb \myif.out[12]~116 (
// Equation(s):
// myifout_12 = (\myif.out[13]~87_combout  & ((\myif.out[12]~115_combout  & (!\out~39_combout )) # (!\myif.out[12]~115_combout  & ((\myif.out[12]~112_combout ))))) # (!\myif.out[13]~87_combout  & (((\myif.out[12]~115_combout ))))

	.dataa(\myif.out[13]~87_combout ),
	.datab(\out~39_combout ),
	.datac(\myif.out[12]~115_combout ),
	.datad(\myif.out[12]~112_combout ),
	.cin(gnd),
	.combout(myifout_12),
	.cout());
// synopsys translate_off
defparam \myif.out[12]~116 .lut_mask = 16'h7A70;
defparam \myif.out[12]~116 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N4
cycloneive_lcell_comb \myif.out[15]~122 (
// Equation(s):
// myifout_15 = (\myif.out[13]~88_combout  & ((\myif.out[15]~121_combout  & (!\out~42_combout )) # (!\myif.out[15]~121_combout  & ((\Add1~30_combout ))))) # (!\myif.out[13]~88_combout  & (((\myif.out[15]~121_combout ))))

	.dataa(\out~42_combout ),
	.datab(\myif.out[13]~88_combout ),
	.datac(\Add1~30_combout ),
	.datad(\myif.out[15]~121_combout ),
	.cin(gnd),
	.combout(myifout_15),
	.cout());
// synopsys translate_off
defparam \myif.out[15]~122 .lut_mask = 16'h77C0;
defparam \myif.out[15]~122 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N30
cycloneive_lcell_comb \myif.out[10]~128 (
// Equation(s):
// myifout_10 = (\myif.out[13]~87_combout  & ((\myif.out[10]~127_combout  & (!\out~45_combout )) # (!\myif.out[10]~127_combout  & ((\myif.out[10]~124_combout ))))) # (!\myif.out[13]~87_combout  & (((\myif.out[10]~127_combout ))))

	.dataa(\myif.out[13]~87_combout ),
	.datab(\out~45_combout ),
	.datac(\myif.out[10]~124_combout ),
	.datad(\myif.out[10]~127_combout ),
	.cin(gnd),
	.combout(myifout_10),
	.cout());
// synopsys translate_off
defparam \myif.out[10]~128 .lut_mask = 16'h77A0;
defparam \myif.out[10]~128 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N4
cycloneive_lcell_comb \myif.out[11]~134 (
// Equation(s):
// myifout_11 = (\myif.out[13]~88_combout  & ((\myif.out[11]~133_combout  & ((!\out~48_combout ))) # (!\myif.out[11]~133_combout  & (\Add1~22_combout )))) # (!\myif.out[13]~88_combout  & (((\myif.out[11]~133_combout ))))

	.dataa(\Add1~22_combout ),
	.datab(\out~48_combout ),
	.datac(\myif.out[13]~88_combout ),
	.datad(\myif.out[11]~133_combout ),
	.cin(gnd),
	.combout(myifout_11),
	.cout());
// synopsys translate_off
defparam \myif.out[11]~134 .lut_mask = 16'h3FA0;
defparam \myif.out[11]~134 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N28
cycloneive_lcell_comb \myif.out[23]~152 (
// Equation(s):
// myifout_23 = (\myif.out[23]~135_combout  & (((\myif.out[23]~151_combout )))) # (!\myif.out[23]~135_combout  & ((\myif.out[23]~151_combout  & ((\myif.out[23]~149_combout ))) # (!\myif.out[23]~151_combout  & (\myif.out[23]~137_combout ))))

	.dataa(\myif.out[23]~135_combout ),
	.datab(\myif.out[23]~137_combout ),
	.datac(\myif.out[23]~151_combout ),
	.datad(\myif.out[23]~149_combout ),
	.cin(gnd),
	.combout(myifout_23),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~152 .lut_mask = 16'hF4A4;
defparam \myif.out[23]~152 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N2
cycloneive_lcell_comb \myif.out[16]~158 (
// Equation(s):
// myifout_16 = (\myif.out[23]~135_combout  & ((\myif.out[16]~157_combout  & ((\out~54_combout ))) # (!\myif.out[16]~157_combout  & (\Add0~32_combout )))) # (!\myif.out[23]~135_combout  & (((\myif.out[16]~157_combout ))))

	.dataa(\Add0~32_combout ),
	.datab(\out~54_combout ),
	.datac(\myif.out[23]~135_combout ),
	.datad(\myif.out[16]~157_combout ),
	.cin(gnd),
	.combout(myifout_16),
	.cout());
// synopsys translate_off
defparam \myif.out[16]~158 .lut_mask = 16'hCFA0;
defparam \myif.out[16]~158 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N10
cycloneive_lcell_comb \myif.out[17]~174 (
// Equation(s):
// myifout_17 = (\myif.out[23]~135_combout  & (((\myif.out[17]~173_combout )))) # (!\myif.out[23]~135_combout  & ((\myif.out[17]~173_combout  & ((\myif.out[17]~172_combout ))) # (!\myif.out[17]~173_combout  & (\myif.out[17]~160_combout ))))

	.dataa(\myif.out[17]~160_combout ),
	.datab(\myif.out[23]~135_combout ),
	.datac(\myif.out[17]~172_combout ),
	.datad(\myif.out[17]~173_combout ),
	.cin(gnd),
	.combout(myifout_17),
	.cout());
// synopsys translate_off
defparam \myif.out[17]~174 .lut_mask = 16'hFC22;
defparam \myif.out[17]~174 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N4
cycloneive_lcell_comb \myif.out[18]~180 (
// Equation(s):
// myifout_18 = (\myif.out[23]~135_combout  & ((\myif.out[18]~179_combout  & (\out~58_combout )) # (!\myif.out[18]~179_combout  & ((\Add0~36_combout ))))) # (!\myif.out[23]~135_combout  & (((\myif.out[18]~179_combout ))))

	.dataa(\myif.out[23]~135_combout ),
	.datab(\out~58_combout ),
	.datac(\Add0~36_combout ),
	.datad(\myif.out[18]~179_combout ),
	.cin(gnd),
	.combout(myifout_18),
	.cout());
// synopsys translate_off
defparam \myif.out[18]~180 .lut_mask = 16'hDDA0;
defparam \myif.out[18]~180 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N2
cycloneive_lcell_comb \myif.out[19]~196 (
// Equation(s):
// myifout_19 = (\myif.out[23]~135_combout  & (\myif.out[19]~195_combout )) # (!\myif.out[23]~135_combout  & ((\myif.out[19]~195_combout  & (\myif.out[19]~182_combout )) # (!\myif.out[19]~195_combout  & ((\myif.out[19]~194_combout )))))

	.dataa(\myif.out[23]~135_combout ),
	.datab(\myif.out[19]~195_combout ),
	.datac(\myif.out[19]~182_combout ),
	.datad(\myif.out[19]~194_combout ),
	.cin(gnd),
	.combout(myifout_19),
	.cout());
// synopsys translate_off
defparam \myif.out[19]~196 .lut_mask = 16'hD9C8;
defparam \myif.out[19]~196 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N30
cycloneive_lcell_comb \myif.out[30]~204 (
// Equation(s):
// myifout_30 = (\myif.out[23]~135_combout  & ((\myif.out[30]~203_combout  & (\out~62_combout )) # (!\myif.out[30]~203_combout  & ((\Add0~60_combout ))))) # (!\myif.out[23]~135_combout  & (((\myif.out[30]~203_combout ))))

	.dataa(\out~62_combout ),
	.datab(\myif.out[23]~135_combout ),
	.datac(\Add0~60_combout ),
	.datad(\myif.out[30]~203_combout ),
	.cin(gnd),
	.combout(myifout_30),
	.cout());
// synopsys translate_off
defparam \myif.out[30]~204 .lut_mask = 16'hBBC0;
defparam \myif.out[30]~204 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N10
cycloneive_lcell_comb \myif.out[21]~220 (
// Equation(s):
// myifout_21 = (\myif.out[23]~135_combout  & (\myif.out[21]~219_combout )) # (!\myif.out[23]~135_combout  & ((\myif.out[21]~219_combout  & ((\myif.out[21]~218_combout ))) # (!\myif.out[21]~219_combout  & (\myif.out[21]~206_combout ))))

	.dataa(\myif.out[23]~135_combout ),
	.datab(\myif.out[21]~219_combout ),
	.datac(\myif.out[21]~206_combout ),
	.datad(\myif.out[21]~218_combout ),
	.cin(gnd),
	.combout(myifout_21),
	.cout());
// synopsys translate_off
defparam \myif.out[21]~220 .lut_mask = 16'hDC98;
defparam \myif.out[21]~220 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N24
cycloneive_lcell_comb \myif.negative~8 (
// Equation(s):
// myifnegative = (\myif.out[23]~150_combout  & ((\myif.negative~7_combout  & (\out~66_combout )) # (!\myif.negative~7_combout  & ((\myif.negative~2_combout ))))) # (!\myif.out[23]~150_combout  & (((\myif.negative~7_combout ))))

	.dataa(\myif.out[23]~150_combout ),
	.datab(\out~66_combout ),
	.datac(\myif.negative~2_combout ),
	.datad(\myif.negative~7_combout ),
	.cin(gnd),
	.combout(myifnegative),
	.cout());
// synopsys translate_off
defparam \myif.negative~8 .lut_mask = 16'hDDA0;
defparam \myif.negative~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N12
cycloneive_lcell_comb \myif.out[22]~226 (
// Equation(s):
// myifout_22 = (\myif.out[23]~135_combout  & ((\myif.out[22]~225_combout  & (\out~69_combout )) # (!\myif.out[22]~225_combout  & ((\Add0~44_combout ))))) # (!\myif.out[23]~135_combout  & (((\myif.out[22]~225_combout ))))

	.dataa(\out~69_combout ),
	.datab(\myif.out[23]~135_combout ),
	.datac(\myif.out[22]~225_combout ),
	.datad(\Add0~44_combout ),
	.cin(gnd),
	.combout(myifout_22),
	.cout());
// synopsys translate_off
defparam \myif.out[22]~226 .lut_mask = 16'hBCB0;
defparam \myif.out[22]~226 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N30
cycloneive_lcell_comb \myif.out[20]~232 (
// Equation(s):
// myifout_20 = (\myif.out[23]~135_combout  & ((\myif.out[20]~231_combout  & (\out~72_combout )) # (!\myif.out[20]~231_combout  & ((\Add0~40_combout ))))) # (!\myif.out[23]~135_combout  & (((\myif.out[20]~231_combout ))))

	.dataa(\myif.out[23]~135_combout ),
	.datab(\out~72_combout ),
	.datac(\Add0~40_combout ),
	.datad(\myif.out[20]~231_combout ),
	.cin(gnd),
	.combout(myifout_20),
	.cout());
// synopsys translate_off
defparam \myif.out[20]~232 .lut_mask = 16'hDDA0;
defparam \myif.out[20]~232 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N10
cycloneive_lcell_comb \myif.out[0]~239 (
// Equation(s):
// myifout_0 = (\myif.out[0]~295_combout ) # ((!idex_ifaluop_o_3 & (idex_ifaluop_o_1 & \myif.out[0]~238_combout )))

	.dataa(idex_ifaluop_o_3),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[0]~238_combout ),
	.datad(\myif.out[0]~295_combout ),
	.cin(gnd),
	.combout(myifout_0),
	.cout());
// synopsys translate_off
defparam \myif.out[0]~239 .lut_mask = 16'hFF40;
defparam \myif.out[0]~239 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N16
cycloneive_lcell_comb \Equal10~10 (
// Equation(s):
// Equal10 = (\Equal10~9_combout  & (!myifout_0 & (\Equal10~7_combout  & \Equal10~2_combout )))

	.dataa(\Equal10~9_combout ),
	.datab(myifout_0),
	.datac(\Equal10~7_combout ),
	.datad(\Equal10~2_combout ),
	.cin(gnd),
	.combout(Equal10),
	.cout());
// synopsys translate_off
defparam \Equal10~10 .lut_mask = 16'h2000;
defparam \Equal10~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N20
cycloneive_lcell_comb \myif.out[28]~252 (
// Equation(s):
// myifout_28 = (\myif.out[28]~293_combout ) # ((\myif.out[28]~290_combout  & ((\myif.out[28]~244_combout ) # (\myif.out[28]~248_combout ))))

	.dataa(\myif.out[28]~293_combout ),
	.datab(\myif.out[28]~244_combout ),
	.datac(\myif.out[28]~248_combout ),
	.datad(\myif.out[28]~290_combout ),
	.cin(gnd),
	.combout(myifout_28),
	.cout());
// synopsys translate_off
defparam \myif.out[28]~252 .lut_mask = 16'hFEAA;
defparam \myif.out[28]~252 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N16
cycloneive_lcell_comb \myif.out[29]~264 (
// Equation(s):
// myifout_29 = (\myif.out[29]~263_combout  & ((\myif.out[29]~259_combout ) # ((\myif.out[28]~250_combout  & \myif.out[29]~258_combout )))) # (!\myif.out[29]~263_combout  & (\myif.out[28]~250_combout  & ((\myif.out[29]~258_combout ))))

	.dataa(\myif.out[29]~263_combout ),
	.datab(\myif.out[28]~250_combout ),
	.datac(\myif.out[29]~259_combout ),
	.datad(\myif.out[29]~258_combout ),
	.cin(gnd),
	.combout(myifout_29),
	.cout());
// synopsys translate_off
defparam \myif.out[29]~264 .lut_mask = 16'hECA0;
defparam \myif.out[29]~264 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N28
cycloneive_lcell_comb \myif.out[2]~274 (
// Equation(s):
// myifout_2 = (\myif.out[5]~245_combout  & ((\myif.out[2]~272_combout ) # ((\myif.out[3]~273_combout  & !\out~76_combout )))) # (!\myif.out[5]~245_combout  & (\myif.out[3]~273_combout  & (!\out~76_combout )))

	.dataa(\myif.out[5]~245_combout ),
	.datab(\myif.out[3]~273_combout ),
	.datac(\out~76_combout ),
	.datad(\myif.out[2]~272_combout ),
	.cin(gnd),
	.combout(myifout_2),
	.cout());
// synopsys translate_off
defparam \myif.out[2]~274 .lut_mask = 16'hAE0C;
defparam \myif.out[2]~274 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N22
cycloneive_lcell_comb \myif.out[3]~283 (
// Equation(s):
// myifout_3 = (\myif.out[3]~240_combout  & ((\myif.out[3]~282_combout  & (\Add1~6_combout )) # (!\myif.out[3]~282_combout  & ((\ShiftRight0~105_combout ))))) # (!\myif.out[3]~240_combout  & (((\myif.out[3]~282_combout ))))

	.dataa(\Add1~6_combout ),
	.datab(\myif.out[3]~240_combout ),
	.datac(\myif.out[3]~282_combout ),
	.datad(\ShiftRight0~105_combout ),
	.cin(gnd),
	.combout(myifout_3),
	.cout());
// synopsys translate_off
defparam \myif.out[3]~283 .lut_mask = 16'hBCB0;
defparam \myif.out[3]~283 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N22
cycloneive_lcell_comb \myif.out[3]~285 (
// Equation(s):
// myifout_31 = (!\myif.out[3]~246_combout  & (\myif.out[5]~284_combout  & ((!\ShiftLeft0~11_combout ) # (!\myif.out[1]~8_combout ))))

	.dataa(\myif.out[1]~8_combout ),
	.datab(\myif.out[3]~246_combout ),
	.datac(\myif.out[5]~284_combout ),
	.datad(\ShiftLeft0~11_combout ),
	.cin(gnd),
	.combout(myifout_31),
	.cout());
// synopsys translate_off
defparam \myif.out[3]~285 .lut_mask = 16'h1030;
defparam \myif.out[3]~285 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N30
cycloneive_lcell_comb \myif.out[2]~289 (
// Equation(s):
// myifout_210 = (\myif.out[1]~8_combout  & (((\myif.out[2]~288_combout )))) # (!\myif.out[1]~8_combout  & ((\myif.out[2]~288_combout  & (\Add1~4_combout )) # (!\myif.out[2]~288_combout  & ((\out~76_combout )))))

	.dataa(\myif.out[1]~8_combout ),
	.datab(\Add1~4_combout ),
	.datac(\out~76_combout ),
	.datad(\myif.out[2]~288_combout ),
	.cin(gnd),
	.combout(myifout_210),
	.cout());
// synopsys translate_off
defparam \myif.out[2]~289 .lut_mask = 16'hEE50;
defparam \myif.out[2]~289 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N4
cycloneive_lcell_comb \Equal10~12 (
// Equation(s):
// Equal101 = (!myifout_29 & (!myifout_2 & (\Equal10~11_combout  & !myifout_28)))

	.dataa(myifout_29),
	.datab(myifout_2),
	.datac(\Equal10~11_combout ),
	.datad(myifout_28),
	.cin(gnd),
	.combout(Equal101),
	.cout());
// synopsys translate_off
defparam \Equal10~12 .lut_mask = 16'h0010;
defparam \Equal10~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N24
cycloneive_lcell_comb \myif.out[3]~291 (
// Equation(s):
// myifout_32 = (\myif.out[3]~275_combout ) # ((!idex_ifaluop_o_0 & (!idex_ifaluop_o_3 & \myif.out[3]~279_combout )))

	.dataa(idex_ifaluop_o_0),
	.datab(idex_ifaluop_o_3),
	.datac(\myif.out[3]~279_combout ),
	.datad(\myif.out[3]~275_combout ),
	.cin(gnd),
	.combout(myifout_32),
	.cout());
// synopsys translate_off
defparam \myif.out[3]~291 .lut_mask = 16'hFF10;
defparam \myif.out[3]~291 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N12
cycloneive_lcell_comb \myif.out[1]~10 (
// Equation(s):
// \myif.out[1]~10_combout  = (\port_b~3_combout ) # ((\port_b~0_combout  & fuifrtReplace_1))

	.dataa(port_b1),
	.datab(port_b),
	.datac(gnd),
	.datad(fuifrtReplace_1),
	.cin(gnd),
	.combout(\myif.out[1]~10_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[1]~10 .lut_mask = 16'hEEAA;
defparam \myif.out[1]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N24
cycloneive_lcell_comb \myif.out[1]~11 (
// Equation(s):
// \myif.out[1]~11_combout  = (idex_ifaluop_o_2 & (\rdat1[1]~1_combout  & ((\myif.out[1]~10_combout )))) # (!idex_ifaluop_o_2 & (((!\port_b~17_combout ))))

	.dataa(rdat1_1),
	.datab(idex_ifaluop_o_2),
	.datac(port_b8),
	.datad(\myif.out[1]~10_combout ),
	.cin(gnd),
	.combout(\myif.out[1]~11_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[1]~11 .lut_mask = 16'h8B03;
defparam \myif.out[1]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N30
cycloneive_lcell_comb \ShiftLeft0~4 (
// Equation(s):
// \ShiftLeft0~4_combout  = (\port_b~38_combout ) # ((\port_b~36_combout ) # ((\port_b~40_combout ) # (\port_b~42_combout )))

	.dataa(port_b28),
	.datab(port_b26),
	.datac(port_b30),
	.datad(port_b32),
	.cin(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~4 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N10
cycloneive_lcell_comb \ShiftLeft0~7 (
// Equation(s):
// \ShiftLeft0~7_combout  = (\port_b~61_combout ) # ((\port_b~60_combout ) # ((\port_b~0_combout  & fuifrtReplace_14)))

	.dataa(port_b),
	.datab(fuifrtReplace_14),
	.datac(port_b51),
	.datad(port_b50),
	.cin(gnd),
	.combout(\ShiftLeft0~7_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~7 .lut_mask = 16'hFFF8;
defparam \ShiftLeft0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N24
cycloneive_lcell_comb \ShiftLeft0~5 (
// Equation(s):
// \ShiftLeft0~5_combout  = (\port_b~48_combout ) # ((\port_b~50_combout ) # ((\port_b~46_combout ) # (\port_b~44_combout )))

	.dataa(port_b38),
	.datab(port_b40),
	.datac(port_b36),
	.datad(port_b34),
	.cin(gnd),
	.combout(\ShiftLeft0~5_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~5 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N20
cycloneive_lcell_comb \ShiftLeft0~8 (
// Equation(s):
// \ShiftLeft0~8_combout  = (\port_b~68_combout ) # ((\port_b~67_combout ) # ((\port_b~0_combout  & fuifrtReplace_12)))

	.dataa(port_b58),
	.datab(port_b),
	.datac(port_b57),
	.datad(fuifrtReplace_12),
	.cin(gnd),
	.combout(\ShiftLeft0~8_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~8 .lut_mask = 16'hFEFA;
defparam \ShiftLeft0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N20
cycloneive_lcell_comb \ShiftLeft0~9 (
// Equation(s):
// \ShiftLeft0~9_combout  = (\port_b~63_combout ) # ((\port_b~70_combout ) # ((\port_b~65_combout ) # (\ShiftLeft0~8_combout )))

	.dataa(port_b53),
	.datab(port_b60),
	.datac(port_b55),
	.datad(\ShiftLeft0~8_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~9_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~9 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N14
cycloneive_lcell_comb \ShiftLeft0~10 (
// Equation(s):
// \ShiftLeft0~10_combout  = (\ShiftLeft0~6_combout ) # ((\ShiftLeft0~7_combout ) # ((\ShiftLeft0~5_combout ) # (\ShiftLeft0~9_combout )))

	.dataa(\ShiftLeft0~6_combout ),
	.datab(\ShiftLeft0~7_combout ),
	.datac(\ShiftLeft0~5_combout ),
	.datad(\ShiftLeft0~9_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~10_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~10 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N24
cycloneive_lcell_comb \ShiftLeft0~2 (
// Equation(s):
// \ShiftLeft0~2_combout  = (\port_b~20_combout ) # ((\port_b~26_combout ) # ((\port_b~24_combout ) # (\port_b~22_combout )))

	.dataa(port_b10),
	.datab(port_b16),
	.datac(port_b14),
	.datad(port_b12),
	.cin(gnd),
	.combout(\ShiftLeft0~2_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~2 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N24
cycloneive_lcell_comb \ShiftLeft0~11 (
// Equation(s):
// \ShiftLeft0~11_combout  = (\ShiftLeft0~3_combout ) # ((\ShiftLeft0~4_combout ) # ((\ShiftLeft0~10_combout ) # (\ShiftLeft0~2_combout )))

	.dataa(\ShiftLeft0~3_combout ),
	.datab(\ShiftLeft0~4_combout ),
	.datac(\ShiftLeft0~10_combout ),
	.datad(\ShiftLeft0~2_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~11_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~11 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N26
cycloneive_lcell_comb \myif.out[1]~13 (
// Equation(s):
// \myif.out[1]~13_combout  = (idex_ifaluop_o_2) # ((\ShiftLeft0~14_combout  & !\ShiftLeft0~11_combout ))

	.dataa(\ShiftLeft0~14_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(gnd),
	.datad(\ShiftLeft0~11_combout ),
	.cin(gnd),
	.combout(\myif.out[1]~13_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[1]~13 .lut_mask = 16'hCCEE;
defparam \myif.out[1]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N0
cycloneive_lcell_comb \Add0~0 (
// Equation(s):
// \Add0~0_combout  = (\rdat1[0]~3_combout  & (\port_b~7_combout  $ (VCC))) # (!\rdat1[0]~3_combout  & (\port_b~7_combout  & VCC))
// \Add0~1  = CARRY((\rdat1[0]~3_combout  & \port_b~7_combout ))

	.dataa(rdat1_0),
	.datab(port_b4),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
// synopsys translate_off
defparam \Add0~0 .lut_mask = 16'h6688;
defparam \Add0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N2
cycloneive_lcell_comb \Add0~2 (
// Equation(s):
// \Add0~2_combout  = (\port_b~4_combout  & ((\rdat1[1]~1_combout  & (\Add0~1  & VCC)) # (!\rdat1[1]~1_combout  & (!\Add0~1 )))) # (!\port_b~4_combout  & ((\rdat1[1]~1_combout  & (!\Add0~1 )) # (!\rdat1[1]~1_combout  & ((\Add0~1 ) # (GND)))))
// \Add0~3  = CARRY((\port_b~4_combout  & (!\rdat1[1]~1_combout  & !\Add0~1 )) # (!\port_b~4_combout  & ((!\Add0~1 ) # (!\rdat1[1]~1_combout ))))

	.dataa(port_b2),
	.datab(rdat1_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
// synopsys translate_off
defparam \Add0~2 .lut_mask = 16'h9617;
defparam \Add0~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N28
cycloneive_lcell_comb \myif.out[1]~12 (
// Equation(s):
// \myif.out[1]~12_combout  = (idex_ifaluop_o_2 & (\myif.out[1]~10_combout  $ (((\rdat1[1]~1_combout ))))) # (!idex_ifaluop_o_2 & (((\Add0~2_combout ))))

	.dataa(\myif.out[1]~10_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\Add0~2_combout ),
	.datad(rdat1_1),
	.cin(gnd),
	.combout(\myif.out[1]~12_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[1]~12 .lut_mask = 16'h74B8;
defparam \myif.out[1]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N8
cycloneive_lcell_comb \myif.out[1]~14 (
// Equation(s):
// \myif.out[1]~14_combout  = (idex_ifaluop_o_1 & (((\myif.out[1]~12_combout )))) # (!idex_ifaluop_o_1 & (\myif.out[1]~11_combout  & (\myif.out[1]~13_combout )))

	.dataa(idex_ifaluop_o_1),
	.datab(\myif.out[1]~11_combout ),
	.datac(\myif.out[1]~13_combout ),
	.datad(\myif.out[1]~12_combout ),
	.cin(gnd),
	.combout(\myif.out[1]~14_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[1]~14 .lut_mask = 16'hEA40;
defparam \myif.out[1]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N16
cycloneive_lcell_comb \myif.out[1]~8 (
// Equation(s):
// \myif.out[1]~8_combout  = (!idex_ifaluop_o_2 & !idex_ifaluop_o_1)

	.dataa(idex_ifaluop_o_2),
	.datab(gnd),
	.datac(gnd),
	.datad(idex_ifaluop_o_1),
	.cin(gnd),
	.combout(\myif.out[1]~8_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[1]~8 .lut_mask = 16'h0055;
defparam \myif.out[1]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N14
cycloneive_lcell_comb \myif.out[1]~6 (
// Equation(s):
// \myif.out[1]~6_combout  = (!\port_b~3_combout  & (!\rdat1[1]~1_combout  & ((!\port_b~0_combout ) # (!fuifrtReplace_1))))

	.dataa(port_b1),
	.datab(fuifrtReplace_1),
	.datac(port_b),
	.datad(rdat1_1),
	.cin(gnd),
	.combout(\myif.out[1]~6_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[1]~6 .lut_mask = 16'h0015;
defparam \myif.out[1]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N0
cycloneive_lcell_comb \Add1~0 (
// Equation(s):
// \Add1~0_combout  = (\rdat1[0]~3_combout  & ((GND) # (!\port_b~7_combout ))) # (!\rdat1[0]~3_combout  & (\port_b~7_combout  $ (GND)))
// \Add1~1  = CARRY((\rdat1[0]~3_combout ) # (!\port_b~7_combout ))

	.dataa(rdat1_0),
	.datab(port_b4),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h66BB;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N2
cycloneive_lcell_comb \Add1~2 (
// Equation(s):
// \Add1~2_combout  = (\port_b~4_combout  & ((\rdat1[1]~1_combout  & (!\Add1~1 )) # (!\rdat1[1]~1_combout  & ((\Add1~1 ) # (GND))))) # (!\port_b~4_combout  & ((\rdat1[1]~1_combout  & (\Add1~1  & VCC)) # (!\rdat1[1]~1_combout  & (!\Add1~1 ))))
// \Add1~3  = CARRY((\port_b~4_combout  & ((!\Add1~1 ) # (!\rdat1[1]~1_combout ))) # (!\port_b~4_combout  & (!\rdat1[1]~1_combout  & !\Add1~1 )))

	.dataa(port_b2),
	.datab(rdat1_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h692B;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N4
cycloneive_lcell_comb \myif.out[1]~7 (
// Equation(s):
// \myif.out[1]~7_combout  = (idex_ifaluop_o_2 & (idex_ifaluop_o_1 $ ((!\myif.out[1]~6_combout )))) # (!idex_ifaluop_o_2 & (idex_ifaluop_o_1 & ((\Add1~2_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(idex_ifaluop_o_2),
	.datac(\myif.out[1]~6_combout ),
	.datad(\Add1~2_combout ),
	.cin(gnd),
	.combout(\myif.out[1]~7_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[1]~7 .lut_mask = 16'hA684;
defparam \myif.out[1]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N30
cycloneive_lcell_comb \ShiftRight0~19 (
// Equation(s):
// \ShiftRight0~19_combout  = (\port_b~7_combout  & ((\port_b~4_combout  & (\rdat1[28]~41_combout )) # (!\port_b~4_combout  & ((\rdat1[26]~43_combout )))))

	.dataa(port_b2),
	.datab(port_b4),
	.datac(rdat1_28),
	.datad(rdat1_26),
	.cin(gnd),
	.combout(\ShiftRight0~19_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~19 .lut_mask = 16'hC480;
defparam \ShiftRight0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N20
cycloneive_lcell_comb \ShiftRight0~20 (
// Equation(s):
// \ShiftRight0~20_combout  = (\port_b~4_combout  & (\rdat1[27]~45_combout )) # (!\port_b~4_combout  & ((\rdat1[25]~47_combout )))

	.dataa(gnd),
	.datab(rdat1_27),
	.datac(rdat1_25),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftRight0~20_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~20 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N22
cycloneive_lcell_comb \ShiftRight0~21 (
// Equation(s):
// \ShiftRight0~21_combout  = (\ShiftRight0~19_combout ) # ((!\port_b~7_combout  & \ShiftRight0~20_combout ))

	.dataa(gnd),
	.datab(port_b4),
	.datac(\ShiftRight0~19_combout ),
	.datad(\ShiftRight0~20_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~21_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~21 .lut_mask = 16'hF3F0;
defparam \ShiftRight0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N4
cycloneive_lcell_comb \ShiftRight0~22 (
// Equation(s):
// \ShiftRight0~22_combout  = (\port_b~14_combout  & ((\port_b~10_combout  & (\ShiftRight0~18_combout )) # (!\port_b~10_combout  & ((\ShiftRight0~21_combout )))))

	.dataa(\ShiftRight0~18_combout ),
	.datab(port_b7),
	.datac(\ShiftRight0~21_combout ),
	.datad(port_b6),
	.cin(gnd),
	.combout(\ShiftRight0~22_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~22 .lut_mask = 16'h88C0;
defparam \ShiftRight0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N24
cycloneive_lcell_comb \ShiftRight0~27 (
// Equation(s):
// \ShiftRight0~27_combout  = (\port_b~4_combout  & ((\rdat1[19]~61_combout ))) # (!\port_b~4_combout  & (\rdat1[17]~63_combout ))

	.dataa(port_b2),
	.datab(rdat1_17),
	.datac(rdat1_19),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~27_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~27 .lut_mask = 16'hE4E4;
defparam \ShiftRight0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N2
cycloneive_lcell_comb \ShiftRight0~26 (
// Equation(s):
// \ShiftRight0~26_combout  = (\port_b~7_combout  & ((\port_b~4_combout  & (\rdat1[20]~57_combout )) # (!\port_b~4_combout  & ((\rdat1[18]~59_combout )))))

	.dataa(port_b4),
	.datab(rdat1_20),
	.datac(rdat1_18),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftRight0~26_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~26 .lut_mask = 16'h88A0;
defparam \ShiftRight0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N8
cycloneive_lcell_comb \ShiftRight0~28 (
// Equation(s):
// \ShiftRight0~28_combout  = (\ShiftRight0~26_combout ) # ((!\port_b~7_combout  & \ShiftRight0~27_combout ))

	.dataa(gnd),
	.datab(port_b4),
	.datac(\ShiftRight0~27_combout ),
	.datad(\ShiftRight0~26_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~28_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~28 .lut_mask = 16'hFF30;
defparam \ShiftRight0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N4
cycloneive_lcell_comb \ShiftRight0~24 (
// Equation(s):
// \ShiftRight0~24_combout  = (\port_b~4_combout  & ((\rdat1[23]~53_combout ))) # (!\port_b~4_combout  & (\rdat1[21]~55_combout ))

	.dataa(gnd),
	.datab(rdat1_21),
	.datac(port_b2),
	.datad(rdat1_23),
	.cin(gnd),
	.combout(\ShiftRight0~24_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~24 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N2
cycloneive_lcell_comb \ShiftRight0~23 (
// Equation(s):
// \ShiftRight0~23_combout  = (\port_b~7_combout  & ((\port_b~4_combout  & (\rdat1[24]~49_combout )) # (!\port_b~4_combout  & ((\rdat1[22]~51_combout )))))

	.dataa(rdat1_24),
	.datab(port_b4),
	.datac(port_b2),
	.datad(rdat1_22),
	.cin(gnd),
	.combout(\ShiftRight0~23_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~23 .lut_mask = 16'h8C80;
defparam \ShiftRight0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N30
cycloneive_lcell_comb \ShiftRight0~25 (
// Equation(s):
// \ShiftRight0~25_combout  = (\ShiftRight0~23_combout ) # ((!\port_b~7_combout  & \ShiftRight0~24_combout ))

	.dataa(gnd),
	.datab(port_b4),
	.datac(\ShiftRight0~24_combout ),
	.datad(\ShiftRight0~23_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~25_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~25 .lut_mask = 16'hFF30;
defparam \ShiftRight0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N10
cycloneive_lcell_comb \ShiftRight0~29 (
// Equation(s):
// \ShiftRight0~29_combout  = (\port_b~10_combout  & ((\ShiftRight0~25_combout ))) # (!\port_b~10_combout  & (\ShiftRight0~28_combout ))

	.dataa(gnd),
	.datab(port_b6),
	.datac(\ShiftRight0~28_combout ),
	.datad(\ShiftRight0~25_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~29_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~29 .lut_mask = 16'hFC30;
defparam \ShiftRight0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N28
cycloneive_lcell_comb \ShiftRight0~30 (
// Equation(s):
// \ShiftRight0~30_combout  = (\ShiftRight0~22_combout ) # ((!\port_b~14_combout  & \ShiftRight0~29_combout ))

	.dataa(gnd),
	.datab(port_b7),
	.datac(\ShiftRight0~22_combout ),
	.datad(\ShiftRight0~29_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~30_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~30 .lut_mask = 16'hF3F0;
defparam \ShiftRight0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N0
cycloneive_lcell_comb \ShiftRight0~12 (
// Equation(s):
// \ShiftRight0~12_combout  = (\port_b~7_combout  & (\rdat1[12]~27_combout )) # (!\port_b~7_combout  & ((\rdat1[11]~29_combout )))

	.dataa(rdat1_12),
	.datab(port_b4),
	.datac(gnd),
	.datad(rdat1_11),
	.cin(gnd),
	.combout(\ShiftRight0~12_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~12 .lut_mask = 16'hBB88;
defparam \ShiftRight0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N24
cycloneive_lcell_comb \ShiftRight0~13 (
// Equation(s):
// \ShiftRight0~13_combout  = (\port_b~7_combout  & (\rdat1[10]~31_combout )) # (!\port_b~7_combout  & ((\rdat1[9]~33_combout )))

	.dataa(port_b4),
	.datab(gnd),
	.datac(rdat1_10),
	.datad(rdat1_9),
	.cin(gnd),
	.combout(\ShiftRight0~13_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~13 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N20
cycloneive_lcell_comb \ShiftRight0~14 (
// Equation(s):
// \ShiftRight0~14_combout  = (\port_b~4_combout  & (\ShiftRight0~12_combout )) # (!\port_b~4_combout  & ((\ShiftRight0~13_combout )))

	.dataa(port_b2),
	.datab(gnd),
	.datac(\ShiftRight0~12_combout ),
	.datad(\ShiftRight0~13_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~14_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~14 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N14
cycloneive_lcell_comb \ShiftRight0~9 (
// Equation(s):
// \ShiftRight0~9_combout  = (\port_b~4_combout  & ((\port_b~7_combout  & ((\rdat1[16]~19_combout ))) # (!\port_b~7_combout  & (\rdat1[15]~21_combout ))))

	.dataa(port_b2),
	.datab(rdat1_15),
	.datac(rdat1_16),
	.datad(port_b4),
	.cin(gnd),
	.combout(\ShiftRight0~9_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~9 .lut_mask = 16'hA088;
defparam \ShiftRight0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N24
cycloneive_lcell_comb \ShiftRight0~10 (
// Equation(s):
// \ShiftRight0~10_combout  = (\port_b~7_combout  & ((\rdat1[14]~23_combout ))) # (!\port_b~7_combout  & (\rdat1[13]~25_combout ))

	.dataa(rdat1_13),
	.datab(gnd),
	.datac(rdat1_14),
	.datad(port_b4),
	.cin(gnd),
	.combout(\ShiftRight0~10_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~10 .lut_mask = 16'hF0AA;
defparam \ShiftRight0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N10
cycloneive_lcell_comb \ShiftRight0~11 (
// Equation(s):
// \ShiftRight0~11_combout  = (\ShiftRight0~9_combout ) # ((!\port_b~4_combout  & \ShiftRight0~10_combout ))

	.dataa(port_b2),
	.datab(gnd),
	.datac(\ShiftRight0~9_combout ),
	.datad(\ShiftRight0~10_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~11_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~11 .lut_mask = 16'hF5F0;
defparam \ShiftRight0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N30
cycloneive_lcell_comb \ShiftRight0~15 (
// Equation(s):
// \ShiftRight0~15_combout  = (\port_b~10_combout  & ((\ShiftRight0~11_combout ))) # (!\port_b~10_combout  & (\ShiftRight0~14_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~14_combout ),
	.datac(port_b6),
	.datad(\ShiftRight0~11_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~15_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~15 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N4
cycloneive_lcell_comb \ShiftRight0~2 (
// Equation(s):
// \ShiftRight0~2_combout  = (!\port_b~4_combout  & ((\port_b~7_combout  & (\rdat1[2]~5_combout )) # (!\port_b~7_combout  & ((\rdat1[1]~1_combout )))))

	.dataa(rdat1_2),
	.datab(port_b2),
	.datac(rdat1_1),
	.datad(port_b4),
	.cin(gnd),
	.combout(\ShiftRight0~2_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~2 .lut_mask = 16'h2230;
defparam \ShiftRight0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N18
cycloneive_lcell_comb \ShiftRight0~3 (
// Equation(s):
// \ShiftRight0~3_combout  = (\port_b~7_combout  & (\rdat1[4]~7_combout )) # (!\port_b~7_combout  & ((\rdat1[3]~9_combout )))

	.dataa(port_b4),
	.datab(gnd),
	.datac(rdat1_41),
	.datad(rdat1_31),
	.cin(gnd),
	.combout(\ShiftRight0~3_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~3 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N12
cycloneive_lcell_comb \ShiftRight0~4 (
// Equation(s):
// \ShiftRight0~4_combout  = (!\port_b~10_combout  & ((\ShiftRight0~2_combout ) # ((\port_b~4_combout  & \ShiftRight0~3_combout ))))

	.dataa(port_b6),
	.datab(\ShiftRight0~2_combout ),
	.datac(port_b2),
	.datad(\ShiftRight0~3_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~4_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~4 .lut_mask = 16'h5444;
defparam \ShiftRight0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N2
cycloneive_lcell_comb \ShiftRight0~5 (
// Equation(s):
// \ShiftRight0~5_combout  = (\port_b~7_combout  & ((\rdat1[8]~11_combout ))) # (!\port_b~7_combout  & (\rdat1[7]~13_combout ))

	.dataa(rdat1_7),
	.datab(gnd),
	.datac(rdat1_8),
	.datad(port_b4),
	.cin(gnd),
	.combout(\ShiftRight0~5_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~5 .lut_mask = 16'hF0AA;
defparam \ShiftRight0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N12
cycloneive_lcell_comb \ShiftRight0~6 (
// Equation(s):
// \ShiftRight0~6_combout  = (\port_b~7_combout  & ((\rdat1[6]~15_combout ))) # (!\port_b~7_combout  & (\rdat1[5]~17_combout ))

	.dataa(rdat1_5),
	.datab(port_b4),
	.datac(gnd),
	.datad(rdat1_6),
	.cin(gnd),
	.combout(\ShiftRight0~6_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~6 .lut_mask = 16'hEE22;
defparam \ShiftRight0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N26
cycloneive_lcell_comb \ShiftRight0~7 (
// Equation(s):
// \ShiftRight0~7_combout  = (\port_b~4_combout  & (\ShiftRight0~5_combout )) # (!\port_b~4_combout  & ((\ShiftRight0~6_combout )))

	.dataa(port_b2),
	.datab(\ShiftRight0~5_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~6_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~7_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~7 .lut_mask = 16'hDD88;
defparam \ShiftRight0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N28
cycloneive_lcell_comb \ShiftRight0~8 (
// Equation(s):
// \ShiftRight0~8_combout  = (!\port_b~14_combout  & ((\ShiftRight0~4_combout ) # ((\port_b~10_combout  & \ShiftRight0~7_combout ))))

	.dataa(port_b6),
	.datab(\ShiftRight0~4_combout ),
	.datac(\ShiftRight0~7_combout ),
	.datad(port_b7),
	.cin(gnd),
	.combout(\ShiftRight0~8_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~8 .lut_mask = 16'h00EC;
defparam \ShiftRight0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N16
cycloneive_lcell_comb \ShiftRight0~16 (
// Equation(s):
// \ShiftRight0~16_combout  = (!\port_b~17_combout  & ((\ShiftRight0~8_combout ) # ((\port_b~14_combout  & \ShiftRight0~15_combout ))))

	.dataa(port_b7),
	.datab(port_b8),
	.datac(\ShiftRight0~15_combout ),
	.datad(\ShiftRight0~8_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~16_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~16 .lut_mask = 16'h3320;
defparam \ShiftRight0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N10
cycloneive_lcell_comb \ShiftRight0~31 (
// Equation(s):
// \ShiftRight0~31_combout  = (\ShiftRight0~16_combout ) # ((\port_b~17_combout  & \ShiftRight0~30_combout ))

	.dataa(gnd),
	.datab(port_b8),
	.datac(\ShiftRight0~30_combout ),
	.datad(\ShiftRight0~16_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~31_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~31 .lut_mask = 16'hFFC0;
defparam \ShiftRight0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N18
cycloneive_lcell_comb \myif.out[1]~9 (
// Equation(s):
// \myif.out[1]~9_combout  = (\myif.out[1]~7_combout ) # ((\myif.out[1]~8_combout  & (!\ShiftLeft0~11_combout  & \ShiftRight0~31_combout )))

	.dataa(\myif.out[1]~8_combout ),
	.datab(\ShiftLeft0~11_combout ),
	.datac(\myif.out[1]~7_combout ),
	.datad(\ShiftRight0~31_combout ),
	.cin(gnd),
	.combout(\myif.out[1]~9_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[1]~9 .lut_mask = 16'hF2F0;
defparam \myif.out[1]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N22
cycloneive_lcell_comb \out~9 (
// Equation(s):
// \out~9_combout  = \rdat1[6]~15_combout  $ (((\port_b~45_combout ) # ((\port_b~0_combout  & fuifrtReplace_6))))

	.dataa(port_b),
	.datab(port_b35),
	.datac(rdat1_6),
	.datad(fuifrtReplace_6),
	.cin(gnd),
	.combout(\out~9_combout ),
	.cout());
// synopsys translate_off
defparam \out~9 .lut_mask = 16'h1E3C;
defparam \out~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N4
cycloneive_lcell_comb \Add0~4 (
// Equation(s):
// \Add0~4_combout  = ((\rdat1[2]~5_combout  $ (\port_b~10_combout  $ (!\Add0~3 )))) # (GND)
// \Add0~5  = CARRY((\rdat1[2]~5_combout  & ((\port_b~10_combout ) # (!\Add0~3 ))) # (!\rdat1[2]~5_combout  & (\port_b~10_combout  & !\Add0~3 )))

	.dataa(rdat1_2),
	.datab(port_b6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
// synopsys translate_off
defparam \Add0~4 .lut_mask = 16'h698E;
defparam \Add0~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N6
cycloneive_lcell_comb \Add0~6 (
// Equation(s):
// \Add0~6_combout  = (\rdat1[3]~9_combout  & ((\port_b~14_combout  & (\Add0~5  & VCC)) # (!\port_b~14_combout  & (!\Add0~5 )))) # (!\rdat1[3]~9_combout  & ((\port_b~14_combout  & (!\Add0~5 )) # (!\port_b~14_combout  & ((\Add0~5 ) # (GND)))))
// \Add0~7  = CARRY((\rdat1[3]~9_combout  & (!\port_b~14_combout  & !\Add0~5 )) # (!\rdat1[3]~9_combout  & ((!\Add0~5 ) # (!\port_b~14_combout ))))

	.dataa(rdat1_31),
	.datab(port_b7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
// synopsys translate_off
defparam \Add0~6 .lut_mask = 16'h9617;
defparam \Add0~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N8
cycloneive_lcell_comb \Add0~8 (
// Equation(s):
// \Add0~8_combout  = ((\rdat1[4]~7_combout  $ (\port_b~17_combout  $ (!\Add0~7 )))) # (GND)
// \Add0~9  = CARRY((\rdat1[4]~7_combout  & ((\port_b~17_combout ) # (!\Add0~7 ))) # (!\rdat1[4]~7_combout  & (\port_b~17_combout  & !\Add0~7 )))

	.dataa(rdat1_41),
	.datab(port_b8),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
// synopsys translate_off
defparam \Add0~8 .lut_mask = 16'h698E;
defparam \Add0~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N10
cycloneive_lcell_comb \Add0~10 (
// Equation(s):
// \Add0~10_combout  = (\port_b~44_combout  & ((\rdat1[5]~17_combout  & (\Add0~9  & VCC)) # (!\rdat1[5]~17_combout  & (!\Add0~9 )))) # (!\port_b~44_combout  & ((\rdat1[5]~17_combout  & (!\Add0~9 )) # (!\rdat1[5]~17_combout  & ((\Add0~9 ) # (GND)))))
// \Add0~11  = CARRY((\port_b~44_combout  & (!\rdat1[5]~17_combout  & !\Add0~9 )) # (!\port_b~44_combout  & ((!\Add0~9 ) # (!\rdat1[5]~17_combout ))))

	.dataa(port_b34),
	.datab(rdat1_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
// synopsys translate_off
defparam \Add0~10 .lut_mask = 16'h9617;
defparam \Add0~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N12
cycloneive_lcell_comb \Add0~12 (
// Equation(s):
// \Add0~12_combout  = ((\port_b~46_combout  $ (\rdat1[6]~15_combout  $ (!\Add0~11 )))) # (GND)
// \Add0~13  = CARRY((\port_b~46_combout  & ((\rdat1[6]~15_combout ) # (!\Add0~11 ))) # (!\port_b~46_combout  & (\rdat1[6]~15_combout  & !\Add0~11 )))

	.dataa(port_b36),
	.datab(rdat1_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
// synopsys translate_off
defparam \Add0~12 .lut_mask = 16'h698E;
defparam \Add0~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N28
cycloneive_lcell_comb \out~10 (
// Equation(s):
// \out~10_combout  = (\rdat1[6]~15_combout  & ((\port_b~45_combout ) # ((\port_b~0_combout  & fuifrtReplace_6))))

	.dataa(port_b),
	.datab(port_b35),
	.datac(rdat1_6),
	.datad(fuifrtReplace_6),
	.cin(gnd),
	.combout(\out~10_combout ),
	.cout());
// synopsys translate_off
defparam \out~10 .lut_mask = 16'hE0C0;
defparam \out~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N26
cycloneive_lcell_comb \ShiftLeft0~18 (
// Equation(s):
// \ShiftLeft0~18_combout  = (\port_b~7_combout  & ((\rdat1[5]~17_combout ))) # (!\port_b~7_combout  & (\rdat1[6]~15_combout ))

	.dataa(gnd),
	.datab(port_b4),
	.datac(rdat1_6),
	.datad(rdat1_5),
	.cin(gnd),
	.combout(\ShiftLeft0~18_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~18 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N24
cycloneive_lcell_comb \ShiftLeft0~17 (
// Equation(s):
// \ShiftLeft0~17_combout  = (\port_b~7_combout  & (\rdat1[3]~9_combout )) # (!\port_b~7_combout  & ((\rdat1[4]~7_combout )))

	.dataa(gnd),
	.datab(port_b4),
	.datac(rdat1_31),
	.datad(rdat1_41),
	.cin(gnd),
	.combout(\ShiftLeft0~17_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~17 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N20
cycloneive_lcell_comb \ShiftLeft0~19 (
// Equation(s):
// \ShiftLeft0~19_combout  = (\port_b~4_combout  & ((\ShiftLeft0~17_combout ))) # (!\port_b~4_combout  & (\ShiftLeft0~18_combout ))

	.dataa(port_b2),
	.datab(gnd),
	.datac(\ShiftLeft0~18_combout ),
	.datad(\ShiftLeft0~17_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~19_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~19 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N18
cycloneive_lcell_comb \ShiftLeft0~20 (
// Equation(s):
// \ShiftLeft0~20_combout  = (!\port_b~14_combout  & ((\port_b~10_combout  & (\ShiftLeft0~16_combout )) # (!\port_b~10_combout  & ((\ShiftLeft0~19_combout )))))

	.dataa(\ShiftLeft0~16_combout ),
	.datab(port_b6),
	.datac(port_b7),
	.datad(\ShiftLeft0~19_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~20_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~20 .lut_mask = 16'h0B08;
defparam \ShiftLeft0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N2
cycloneive_lcell_comb \myif.out[13]~23 (
// Equation(s):
// \myif.out[13]~23_combout  = (!idex_ifaluop_o_1 & ((idex_ifaluop_o_2) # ((!\port_b~17_combout  & !\ShiftLeft0~11_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(idex_ifaluop_o_2),
	.datac(port_b8),
	.datad(\ShiftLeft0~11_combout ),
	.cin(gnd),
	.combout(\myif.out[13]~23_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[13]~23 .lut_mask = 16'h4445;
defparam \myif.out[13]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N10
cycloneive_lcell_comb \myif.out[6]~24 (
// Equation(s):
// \myif.out[6]~24_combout  = (idex_ifaluop_o_2 & ((\out~10_combout ) # ((!\myif.out[13]~23_combout )))) # (!idex_ifaluop_o_2 & (((\ShiftLeft0~20_combout  & \myif.out[13]~23_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\out~10_combout ),
	.datac(\ShiftLeft0~20_combout ),
	.datad(\myif.out[13]~23_combout ),
	.cin(gnd),
	.combout(\myif.out[6]~24_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[6]~24 .lut_mask = 16'hD8AA;
defparam \myif.out[6]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N8
cycloneive_lcell_comb \myif.out[6]~25 (
// Equation(s):
// \myif.out[6]~25_combout  = (idex_ifaluop_o_1 & ((\myif.out[6]~24_combout  & (\out~9_combout )) # (!\myif.out[6]~24_combout  & ((\Add0~12_combout ))))) # (!idex_ifaluop_o_1 & (((\myif.out[6]~24_combout ))))

	.dataa(\out~9_combout ),
	.datab(idex_ifaluop_o_1),
	.datac(\Add0~12_combout ),
	.datad(\myif.out[6]~24_combout ),
	.cin(gnd),
	.combout(\myif.out[6]~25_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[6]~25 .lut_mask = 16'hBBC0;
defparam \myif.out[6]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N22
cycloneive_lcell_comb \out~8 (
// Equation(s):
// \out~8_combout  = (\rdat1[6]~15_combout ) # ((\port_b~45_combout ) # ((\port_b~0_combout  & fuifrtReplace_6)))

	.dataa(port_b),
	.datab(rdat1_6),
	.datac(port_b35),
	.datad(fuifrtReplace_6),
	.cin(gnd),
	.combout(\out~8_combout ),
	.cout());
// synopsys translate_off
defparam \out~8 .lut_mask = 16'hFEFC;
defparam \out~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N4
cycloneive_lcell_comb \Add1~4 (
// Equation(s):
// \Add1~4_combout  = ((\rdat1[2]~5_combout  $ (\port_b~10_combout  $ (\Add1~3 )))) # (GND)
// \Add1~5  = CARRY((\rdat1[2]~5_combout  & ((!\Add1~3 ) # (!\port_b~10_combout ))) # (!\rdat1[2]~5_combout  & (!\port_b~10_combout  & !\Add1~3 )))

	.dataa(rdat1_2),
	.datab(port_b6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'h962B;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N6
cycloneive_lcell_comb \Add1~6 (
// Equation(s):
// \Add1~6_combout  = (\port_b~14_combout  & ((\rdat1[3]~9_combout  & (!\Add1~5 )) # (!\rdat1[3]~9_combout  & ((\Add1~5 ) # (GND))))) # (!\port_b~14_combout  & ((\rdat1[3]~9_combout  & (\Add1~5  & VCC)) # (!\rdat1[3]~9_combout  & (!\Add1~5 ))))
// \Add1~7  = CARRY((\port_b~14_combout  & ((!\Add1~5 ) # (!\rdat1[3]~9_combout ))) # (!\port_b~14_combout  & (!\rdat1[3]~9_combout  & !\Add1~5 )))

	.dataa(port_b7),
	.datab(rdat1_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h692B;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N8
cycloneive_lcell_comb \Add1~8 (
// Equation(s):
// \Add1~8_combout  = ((\rdat1[4]~7_combout  $ (\port_b~17_combout  $ (\Add1~7 )))) # (GND)
// \Add1~9  = CARRY((\rdat1[4]~7_combout  & ((!\Add1~7 ) # (!\port_b~17_combout ))) # (!\rdat1[4]~7_combout  & (!\port_b~17_combout  & !\Add1~7 )))

	.dataa(rdat1_41),
	.datab(port_b8),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'h962B;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N10
cycloneive_lcell_comb \Add1~10 (
// Equation(s):
// \Add1~10_combout  = (\port_b~44_combout  & ((\rdat1[5]~17_combout  & (!\Add1~9 )) # (!\rdat1[5]~17_combout  & ((\Add1~9 ) # (GND))))) # (!\port_b~44_combout  & ((\rdat1[5]~17_combout  & (\Add1~9  & VCC)) # (!\rdat1[5]~17_combout  & (!\Add1~9 ))))
// \Add1~11  = CARRY((\port_b~44_combout  & ((!\Add1~9 ) # (!\rdat1[5]~17_combout ))) # (!\port_b~44_combout  & (!\rdat1[5]~17_combout  & !\Add1~9 )))

	.dataa(port_b34),
	.datab(rdat1_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h692B;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N12
cycloneive_lcell_comb \Add1~12 (
// Equation(s):
// \Add1~12_combout  = ((\rdat1[6]~15_combout  $ (\port_b~46_combout  $ (\Add1~11 )))) # (GND)
// \Add1~13  = CARRY((\rdat1[6]~15_combout  & ((!\Add1~11 ) # (!\port_b~46_combout ))) # (!\rdat1[6]~15_combout  & (!\port_b~46_combout  & !\Add1~11 )))

	.dataa(rdat1_6),
	.datab(port_b36),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout(\Add1~13 ));
// synopsys translate_off
defparam \Add1~12 .lut_mask = 16'h962B;
defparam \Add1~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N0
cycloneive_lcell_comb \myif.out[5]~20 (
// Equation(s):
// \myif.out[5]~20_combout  = (!idex_ifaluop_o_1 & ((idex_ifaluop_o_2) # (!\ShiftLeft0~11_combout )))

	.dataa(idex_ifaluop_o_1),
	.datab(idex_ifaluop_o_2),
	.datac(gnd),
	.datad(\ShiftLeft0~11_combout ),
	.cin(gnd),
	.combout(\myif.out[5]~20_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[5]~20 .lut_mask = 16'h4455;
defparam \myif.out[5]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N28
cycloneive_lcell_comb \myif.out[5]~16 (
// Equation(s):
// \myif.out[5]~16_combout  = (\port_b~14_combout ) # (\port_b~17_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(port_b7),
	.datad(port_b8),
	.cin(gnd),
	.combout(\myif.out[5]~16_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[5]~16 .lut_mask = 16'hFFF0;
defparam \myif.out[5]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N4
cycloneive_lcell_comb \ShiftRight0~35 (
// Equation(s):
// \ShiftRight0~35_combout  = (\port_b~4_combout  & ((\port_b~7_combout  & (\rdat1[17]~63_combout )) # (!\port_b~7_combout  & ((\rdat1[16]~19_combout )))))

	.dataa(port_b2),
	.datab(rdat1_17),
	.datac(port_b4),
	.datad(rdat1_16),
	.cin(gnd),
	.combout(\ShiftRight0~35_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~35 .lut_mask = 16'h8A80;
defparam \ShiftRight0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N26
cycloneive_lcell_comb \ShiftRight0~36 (
// Equation(s):
// \ShiftRight0~36_combout  = (\port_b~7_combout  & (\rdat1[15]~21_combout )) # (!\port_b~7_combout  & ((\rdat1[14]~23_combout )))

	.dataa(rdat1_15),
	.datab(gnd),
	.datac(rdat1_14),
	.datad(port_b4),
	.cin(gnd),
	.combout(\ShiftRight0~36_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~36 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N26
cycloneive_lcell_comb \ShiftRight0~37 (
// Equation(s):
// \ShiftRight0~37_combout  = (\ShiftRight0~35_combout ) # ((!\port_b~4_combout  & \ShiftRight0~36_combout ))

	.dataa(port_b2),
	.datab(gnd),
	.datac(\ShiftRight0~35_combout ),
	.datad(\ShiftRight0~36_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~37_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~37 .lut_mask = 16'hF5F0;
defparam \ShiftRight0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N14
cycloneive_lcell_comb \ShiftRight0~38 (
// Equation(s):
// \ShiftRight0~38_combout  = (\port_b~10_combout  & (\ShiftRight0~34_combout )) # (!\port_b~10_combout  & ((\ShiftRight0~37_combout )))

	.dataa(\ShiftRight0~34_combout ),
	.datab(port_b6),
	.datac(gnd),
	.datad(\ShiftRight0~37_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~38_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~38 .lut_mask = 16'hBB88;
defparam \ShiftRight0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N8
cycloneive_lcell_comb \ShiftRight0~45 (
// Equation(s):
// \ShiftRight0~45_combout  = (!\port_b~7_combout  & ((\port_b~4_combout  & (\rdat1[28]~41_combout )) # (!\port_b~4_combout  & ((\rdat1[26]~43_combout )))))

	.dataa(port_b4),
	.datab(rdat1_28),
	.datac(rdat1_26),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftRight0~45_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~45 .lut_mask = 16'h4450;
defparam \ShiftRight0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N2
cycloneive_lcell_comb \ShiftRight0~46 (
// Equation(s):
// \ShiftRight0~46_combout  = (\port_b~4_combout  & (\rdat1[29]~37_combout )) # (!\port_b~4_combout  & ((\rdat1[27]~45_combout )))

	.dataa(gnd),
	.datab(rdat1_29),
	.datac(rdat1_27),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftRight0~46_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~46 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N14
cycloneive_lcell_comb \ShiftRight0~47 (
// Equation(s):
// \ShiftRight0~47_combout  = (\ShiftRight0~45_combout ) # ((\port_b~7_combout  & \ShiftRight0~46_combout ))

	.dataa(gnd),
	.datab(port_b4),
	.datac(\ShiftRight0~45_combout ),
	.datad(\ShiftRight0~46_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~47_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~47 .lut_mask = 16'hFCF0;
defparam \ShiftRight0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N30
cycloneive_lcell_comb \ShiftRight0~49 (
// Equation(s):
// \ShiftRight0~49_combout  = (\port_b~4_combout  & (\rdat1[25]~47_combout )) # (!\port_b~4_combout  & ((\rdat1[23]~53_combout )))

	.dataa(rdat1_25),
	.datab(gnd),
	.datac(rdat1_23),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftRight0~49_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~49 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N0
cycloneive_lcell_comb \ShiftRight0~48 (
// Equation(s):
// \ShiftRight0~48_combout  = (!\port_b~7_combout  & ((\port_b~4_combout  & (\rdat1[24]~49_combout )) # (!\port_b~4_combout  & ((\rdat1[22]~51_combout )))))

	.dataa(port_b2),
	.datab(port_b4),
	.datac(rdat1_24),
	.datad(rdat1_22),
	.cin(gnd),
	.combout(\ShiftRight0~48_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~48 .lut_mask = 16'h3120;
defparam \ShiftRight0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N8
cycloneive_lcell_comb \ShiftRight0~50 (
// Equation(s):
// \ShiftRight0~50_combout  = (\ShiftRight0~48_combout ) # ((\port_b~7_combout  & \ShiftRight0~49_combout ))

	.dataa(gnd),
	.datab(port_b4),
	.datac(\ShiftRight0~49_combout ),
	.datad(\ShiftRight0~48_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~50_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~50 .lut_mask = 16'hFFC0;
defparam \ShiftRight0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N30
cycloneive_lcell_comb \ShiftRight0~51 (
// Equation(s):
// \ShiftRight0~51_combout  = (\port_b~10_combout  & (\ShiftRight0~47_combout )) # (!\port_b~10_combout  & ((\ShiftRight0~50_combout )))

	.dataa(gnd),
	.datab(port_b6),
	.datac(\ShiftRight0~47_combout ),
	.datad(\ShiftRight0~50_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~51_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~51 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N30
cycloneive_lcell_comb \ShiftLeft0~13 (
// Equation(s):
// \ShiftLeft0~13_combout  = (\port_b~9_combout ) # ((\port_b~4_combout ) # ((fuifrtReplace_2 & \port_b~0_combout )))

	.dataa(fuifrtReplace_2),
	.datab(port_b),
	.datac(port_b5),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftLeft0~13_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~13 .lut_mask = 16'hFFF8;
defparam \ShiftLeft0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N20
cycloneive_lcell_comb \ShiftRight0~53 (
// Equation(s):
// \ShiftRight0~53_combout  = (\port_b~14_combout  & (\ShiftRight0~52_combout  & ((!\ShiftLeft0~13_combout )))) # (!\port_b~14_combout  & (((\ShiftRight0~51_combout ))))

	.dataa(\ShiftRight0~52_combout ),
	.datab(port_b7),
	.datac(\ShiftRight0~51_combout ),
	.datad(\ShiftLeft0~13_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~53 .lut_mask = 16'h30B8;
defparam \ShiftRight0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N6
cycloneive_lcell_comb \myif.out[6]~19 (
// Equation(s):
// \myif.out[6]~19_combout  = (\myif.out[6]~18_combout  & (((\ShiftRight0~53_combout )) # (!\myif.out[5]~16_combout ))) # (!\myif.out[6]~18_combout  & (\myif.out[5]~16_combout  & (\ShiftRight0~38_combout )))

	.dataa(\myif.out[6]~18_combout ),
	.datab(\myif.out[5]~16_combout ),
	.datac(\ShiftRight0~38_combout ),
	.datad(\ShiftRight0~53_combout ),
	.cin(gnd),
	.combout(\myif.out[6]~19_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[6]~19 .lut_mask = 16'hEA62;
defparam \myif.out[6]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N0
cycloneive_lcell_comb \myif.out[6]~21 (
// Equation(s):
// \myif.out[6]~21_combout  = (idex_ifaluop_o_2 & ((\out~8_combout ) # ((!\myif.out[5]~20_combout )))) # (!idex_ifaluop_o_2 & (((\myif.out[5]~20_combout  & \myif.out[6]~19_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\out~8_combout ),
	.datac(\myif.out[5]~20_combout ),
	.datad(\myif.out[6]~19_combout ),
	.cin(gnd),
	.combout(\myif.out[6]~21_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[6]~21 .lut_mask = 16'hDA8A;
defparam \myif.out[6]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N10
cycloneive_lcell_comb \myif.out[6]~22 (
// Equation(s):
// \myif.out[6]~22_combout  = (idex_ifaluop_o_1 & ((\myif.out[6]~21_combout  & (!\out~8_combout )) # (!\myif.out[6]~21_combout  & ((\Add1~12_combout ))))) # (!idex_ifaluop_o_1 & (((\myif.out[6]~21_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(\out~8_combout ),
	.datac(\Add1~12_combout ),
	.datad(\myif.out[6]~21_combout ),
	.cin(gnd),
	.combout(\myif.out[6]~22_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[6]~22 .lut_mask = 16'h77A0;
defparam \myif.out[6]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N2
cycloneive_lcell_comb \out~77 (
// Equation(s):
// \out~77_combout  = (\rdat1[4]~6_combout ) # ((\port_b~17_combout ) # ((always03 & \mem_data~10_combout )))

	.dataa(always0),
	.datab(rdat1_4),
	.datac(mem_data),
	.datad(port_b8),
	.cin(gnd),
	.combout(\out~77_combout ),
	.cout());
// synopsys translate_off
defparam \out~77 .lut_mask = 16'hFFEC;
defparam \out~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N12
cycloneive_lcell_comb \myif.out[5]~17 (
// Equation(s):
// \myif.out[5]~17_combout  = (\port_b~17_combout ) # ((!\port_b~14_combout  & \port_b~10_combout ))

	.dataa(port_b7),
	.datab(port_b6),
	.datac(port_b8),
	.datad(gnd),
	.cin(gnd),
	.combout(\myif.out[5]~17_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[5]~17 .lut_mask = 16'hF4F4;
defparam \myif.out[5]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N22
cycloneive_lcell_comb \ShiftRight0~43 (
// Equation(s):
// \ShiftRight0~43_combout  = (\port_b~7_combout  & (\rdat1[7]~13_combout )) # (!\port_b~7_combout  & ((\rdat1[6]~15_combout )))

	.dataa(rdat1_7),
	.datab(gnd),
	.datac(rdat1_6),
	.datad(port_b4),
	.cin(gnd),
	.combout(\ShiftRight0~43_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~43 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N20
cycloneive_lcell_comb \ShiftRight0~60 (
// Equation(s):
// \ShiftRight0~60_combout  = (\port_b~4_combout  & ((\ShiftRight0~43_combout ))) # (!\port_b~4_combout  & (\ShiftRight0~59_combout ))

	.dataa(\ShiftRight0~59_combout ),
	.datab(port_b2),
	.datac(gnd),
	.datad(\ShiftRight0~43_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~60 .lut_mask = 16'hEE22;
defparam \ShiftRight0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N8
cycloneive_lcell_comb \ShiftRight0~55 (
// Equation(s):
// \ShiftRight0~55_combout  = (!\port_b~7_combout  & ((\port_b~4_combout  & (\rdat1[18]~59_combout )) # (!\port_b~4_combout  & ((\rdat1[16]~19_combout )))))

	.dataa(port_b2),
	.datab(port_b4),
	.datac(rdat1_18),
	.datad(rdat1_16),
	.cin(gnd),
	.combout(\ShiftRight0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~55 .lut_mask = 16'h3120;
defparam \ShiftRight0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N10
cycloneive_lcell_comb \ShiftRight0~56 (
// Equation(s):
// \ShiftRight0~56_combout  = (\ShiftRight0~55_combout ) # ((\port_b~7_combout  & \ShiftRight0~27_combout ))

	.dataa(gnd),
	.datab(port_b4),
	.datac(\ShiftRight0~55_combout ),
	.datad(\ShiftRight0~27_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~56 .lut_mask = 16'hFCF0;
defparam \ShiftRight0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N16
cycloneive_lcell_comb \ShiftRight0~58 (
// Equation(s):
// \ShiftRight0~58_combout  = (\port_b~10_combout  & ((\ShiftRight0~56_combout ))) # (!\port_b~10_combout  & (\ShiftRight0~57_combout ))

	.dataa(\ShiftRight0~57_combout ),
	.datab(port_b6),
	.datac(gnd),
	.datad(\ShiftRight0~56_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~58 .lut_mask = 16'hEE22;
defparam \ShiftRight0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N22
cycloneive_lcell_comb \myif.out[4]~27 (
// Equation(s):
// \myif.out[4]~27_combout  = (\myif.out[5]~17_combout  & (\myif.out[5]~16_combout )) # (!\myif.out[5]~17_combout  & ((\myif.out[5]~16_combout  & ((\ShiftRight0~58_combout ))) # (!\myif.out[5]~16_combout  & (\ShiftRight0~60_combout ))))

	.dataa(\myif.out[5]~17_combout ),
	.datab(\myif.out[5]~16_combout ),
	.datac(\ShiftRight0~60_combout ),
	.datad(\ShiftRight0~58_combout ),
	.cin(gnd),
	.combout(\myif.out[4]~27_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[4]~27 .lut_mask = 16'hDC98;
defparam \myif.out[4]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N26
cycloneive_lcell_comb \ShiftRight0~61 (
// Equation(s):
// \ShiftRight0~61_combout  = (!\port_b~7_combout  & ((\port_b~4_combout  & ((\rdat1[26]~43_combout ))) # (!\port_b~4_combout  & (\rdat1[24]~49_combout ))))

	.dataa(rdat1_24),
	.datab(rdat1_26),
	.datac(port_b4),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftRight0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~61 .lut_mask = 16'h0C0A;
defparam \ShiftRight0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N28
cycloneive_lcell_comb \ShiftRight0~62 (
// Equation(s):
// \ShiftRight0~62_combout  = (\ShiftRight0~61_combout ) # ((\port_b~7_combout  & \ShiftRight0~20_combout ))

	.dataa(gnd),
	.datab(port_b4),
	.datac(\ShiftRight0~61_combout ),
	.datad(\ShiftRight0~20_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~62 .lut_mask = 16'hFCF0;
defparam \ShiftRight0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N22
cycloneive_lcell_comb \ShiftRight0~63 (
// Equation(s):
// \ShiftRight0~63_combout  = (!\port_b~7_combout  & ((\port_b~4_combout  & ((\rdat1[22]~51_combout ))) # (!\port_b~4_combout  & (\rdat1[20]~57_combout ))))

	.dataa(rdat1_20),
	.datab(port_b4),
	.datac(port_b2),
	.datad(rdat1_22),
	.cin(gnd),
	.combout(\ShiftRight0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~63 .lut_mask = 16'h3202;
defparam \ShiftRight0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N16
cycloneive_lcell_comb \ShiftRight0~64 (
// Equation(s):
// \ShiftRight0~64_combout  = (\ShiftRight0~63_combout ) # ((\ShiftRight0~24_combout  & \port_b~7_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~24_combout ),
	.datac(\ShiftRight0~63_combout ),
	.datad(port_b4),
	.cin(gnd),
	.combout(\ShiftRight0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~64 .lut_mask = 16'hFCF0;
defparam \ShiftRight0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N0
cycloneive_lcell_comb \ShiftRight0~65 (
// Equation(s):
// \ShiftRight0~65_combout  = (\port_b~10_combout  & (\ShiftRight0~62_combout )) # (!\port_b~10_combout  & ((\ShiftRight0~64_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~62_combout ),
	.datac(port_b6),
	.datad(\ShiftRight0~64_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~65 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N2
cycloneive_lcell_comb \ShiftRight0~68 (
// Equation(s):
// \ShiftRight0~68_combout  = (\port_b~14_combout  & (\ShiftRight0~67_combout  & (!\port_b~10_combout ))) # (!\port_b~14_combout  & (((\ShiftRight0~65_combout ))))

	.dataa(\ShiftRight0~67_combout ),
	.datab(port_b6),
	.datac(port_b7),
	.datad(\ShiftRight0~65_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~68 .lut_mask = 16'h2F20;
defparam \ShiftRight0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N16
cycloneive_lcell_comb \myif.out[4]~28 (
// Equation(s):
// \myif.out[4]~28_combout  = (\myif.out[5]~17_combout  & ((\myif.out[4]~27_combout  & ((\ShiftRight0~68_combout ))) # (!\myif.out[4]~27_combout  & (\ShiftRight0~54_combout )))) # (!\myif.out[5]~17_combout  & (((\myif.out[4]~27_combout ))))

	.dataa(\ShiftRight0~54_combout ),
	.datab(\myif.out[5]~17_combout ),
	.datac(\myif.out[4]~27_combout ),
	.datad(\ShiftRight0~68_combout ),
	.cin(gnd),
	.combout(\myif.out[4]~28_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[4]~28 .lut_mask = 16'hF838;
defparam \myif.out[4]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N10
cycloneive_lcell_comb \myif.out[4]~29 (
// Equation(s):
// \myif.out[4]~29_combout  = (idex_ifaluop_o_2 & (((\out~77_combout )) # (!\myif.out[5]~20_combout ))) # (!idex_ifaluop_o_2 & (\myif.out[5]~20_combout  & ((\myif.out[4]~28_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\myif.out[5]~20_combout ),
	.datac(\out~77_combout ),
	.datad(\myif.out[4]~28_combout ),
	.cin(gnd),
	.combout(\myif.out[4]~29_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[4]~29 .lut_mask = 16'hE6A2;
defparam \myif.out[4]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N4
cycloneive_lcell_comb \myif.out[4]~30 (
// Equation(s):
// \myif.out[4]~30_combout  = (idex_ifaluop_o_1 & ((\myif.out[4]~29_combout  & ((!\out~77_combout ))) # (!\myif.out[4]~29_combout  & (\Add1~8_combout )))) # (!idex_ifaluop_o_1 & (((\myif.out[4]~29_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(\Add1~8_combout ),
	.datac(\out~77_combout ),
	.datad(\myif.out[4]~29_combout ),
	.cin(gnd),
	.combout(\myif.out[4]~30_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[4]~30 .lut_mask = 16'h5F88;
defparam \myif.out[4]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N16
cycloneive_lcell_comb \out~78 (
// Equation(s):
// \out~78_combout  = \port_b~17_combout  $ (((\rdat1[4]~6_combout ) # ((always03 & \mem_data~10_combout ))))

	.dataa(always0),
	.datab(rdat1_4),
	.datac(mem_data),
	.datad(port_b8),
	.cin(gnd),
	.combout(\out~78_combout ),
	.cout());
// synopsys translate_off
defparam \out~78 .lut_mask = 16'h13EC;
defparam \out~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N4
cycloneive_lcell_comb \ShiftLeft0~22 (
// Equation(s):
// \ShiftLeft0~22_combout  = (\port_b~4_combout  & ((\port_b~7_combout  & (\rdat1[1]~1_combout )) # (!\port_b~7_combout  & ((\rdat1[2]~5_combout )))))

	.dataa(rdat1_1),
	.datab(rdat1_2),
	.datac(port_b4),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftLeft0~22_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~22 .lut_mask = 16'hAC00;
defparam \ShiftLeft0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N14
cycloneive_lcell_comb \ShiftLeft0~23 (
// Equation(s):
// \ShiftLeft0~23_combout  = (\ShiftLeft0~22_combout ) # ((!\port_b~4_combout  & \ShiftLeft0~17_combout ))

	.dataa(port_b2),
	.datab(gnd),
	.datac(\ShiftLeft0~22_combout ),
	.datad(\ShiftLeft0~17_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~23_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~23 .lut_mask = 16'hF5F0;
defparam \ShiftLeft0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N20
cycloneive_lcell_comb \ShiftLeft0~21 (
// Equation(s):
// \ShiftLeft0~21_combout  = (!\port_b~7_combout  & (\rdat1[0]~3_combout  & !\port_b~4_combout ))

	.dataa(port_b4),
	.datab(rdat1_0),
	.datac(gnd),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftLeft0~21_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~21 .lut_mask = 16'h0044;
defparam \ShiftLeft0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N0
cycloneive_lcell_comb \ShiftLeft0~24 (
// Equation(s):
// \ShiftLeft0~24_combout  = (!\port_b~14_combout  & ((\port_b~10_combout  & ((\ShiftLeft0~21_combout ))) # (!\port_b~10_combout  & (\ShiftLeft0~23_combout ))))

	.dataa(port_b7),
	.datab(\ShiftLeft0~23_combout ),
	.datac(\ShiftLeft0~21_combout ),
	.datad(port_b6),
	.cin(gnd),
	.combout(\ShiftLeft0~24_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~24 .lut_mask = 16'h5044;
defparam \ShiftLeft0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N20
cycloneive_lcell_comb \myif.out[4]~31 (
// Equation(s):
// \myif.out[4]~31_combout  = (idex_ifaluop_o_2 & ((\out~79_combout ) # ((!\myif.out[13]~23_combout )))) # (!idex_ifaluop_o_2 & (((\ShiftLeft0~24_combout  & \myif.out[13]~23_combout ))))

	.dataa(\out~79_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\ShiftLeft0~24_combout ),
	.datad(\myif.out[13]~23_combout ),
	.cin(gnd),
	.combout(\myif.out[4]~31_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[4]~31 .lut_mask = 16'hB8CC;
defparam \myif.out[4]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N10
cycloneive_lcell_comb \myif.out[4]~32 (
// Equation(s):
// \myif.out[4]~32_combout  = (idex_ifaluop_o_1 & ((\myif.out[4]~31_combout  & (\out~78_combout )) # (!\myif.out[4]~31_combout  & ((\Add0~8_combout ))))) # (!idex_ifaluop_o_1 & (((\myif.out[4]~31_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(\out~78_combout ),
	.datac(\Add0~8_combout ),
	.datad(\myif.out[4]~31_combout ),
	.cin(gnd),
	.combout(\myif.out[4]~32_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[4]~32 .lut_mask = 16'hDDA0;
defparam \myif.out[4]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N14
cycloneive_lcell_comb \Add0~14 (
// Equation(s):
// \Add0~14_combout  = (\port_b~48_combout  & ((\rdat1[7]~13_combout  & (\Add0~13  & VCC)) # (!\rdat1[7]~13_combout  & (!\Add0~13 )))) # (!\port_b~48_combout  & ((\rdat1[7]~13_combout  & (!\Add0~13 )) # (!\rdat1[7]~13_combout  & ((\Add0~13 ) # (GND)))))
// \Add0~15  = CARRY((\port_b~48_combout  & (!\rdat1[7]~13_combout  & !\Add0~13 )) # (!\port_b~48_combout  & ((!\Add0~13 ) # (!\rdat1[7]~13_combout ))))

	.dataa(port_b38),
	.datab(rdat1_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
// synopsys translate_off
defparam \Add0~14 .lut_mask = 16'h9617;
defparam \Add0~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N20
cycloneive_lcell_comb \Add0~20 (
// Equation(s):
// \Add0~20_combout  = ((\rdat1[10]~31_combout  $ (\port_b~65_combout  $ (!\Add0~19 )))) # (GND)
// \Add0~21  = CARRY((\rdat1[10]~31_combout  & ((\port_b~65_combout ) # (!\Add0~19 ))) # (!\rdat1[10]~31_combout  & (\port_b~65_combout  & !\Add0~19 )))

	.dataa(rdat1_10),
	.datab(port_b55),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
// synopsys translate_off
defparam \Add0~20 .lut_mask = 16'h698E;
defparam \Add0~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N22
cycloneive_lcell_comb \Add0~22 (
// Equation(s):
// \Add0~22_combout  = (\rdat1[11]~29_combout  & ((\port_b~67_combout  & (\Add0~21  & VCC)) # (!\port_b~67_combout  & (!\Add0~21 )))) # (!\rdat1[11]~29_combout  & ((\port_b~67_combout  & (!\Add0~21 )) # (!\port_b~67_combout  & ((\Add0~21 ) # (GND)))))
// \Add0~23  = CARRY((\rdat1[11]~29_combout  & (!\port_b~67_combout  & !\Add0~21 )) # (!\rdat1[11]~29_combout  & ((!\Add0~21 ) # (!\port_b~67_combout ))))

	.dataa(rdat1_11),
	.datab(port_b57),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
// synopsys translate_off
defparam \Add0~22 .lut_mask = 16'h9617;
defparam \Add0~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N24
cycloneive_lcell_comb \Add0~24 (
// Equation(s):
// \Add0~24_combout  = ((\rdat1[12]~27_combout  $ (\port_b~72_combout  $ (!\Add0~23 )))) # (GND)
// \Add0~25  = CARRY((\rdat1[12]~27_combout  & ((\port_b~72_combout ) # (!\Add0~23 ))) # (!\rdat1[12]~27_combout  & (\port_b~72_combout  & !\Add0~23 )))

	.dataa(rdat1_12),
	.datab(port_b62),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
// synopsys translate_off
defparam \Add0~24 .lut_mask = 16'h698E;
defparam \Add0~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N30
cycloneive_lcell_comb \Add0~30 (
// Equation(s):
// \Add0~30_combout  = (\rdat1[15]~21_combout  & ((\port_b~63_combout  & (\Add0~29  & VCC)) # (!\port_b~63_combout  & (!\Add0~29 )))) # (!\rdat1[15]~21_combout  & ((\port_b~63_combout  & (!\Add0~29 )) # (!\port_b~63_combout  & ((\Add0~29 ) # (GND)))))
// \Add0~31  = CARRY((\rdat1[15]~21_combout  & (!\port_b~63_combout  & !\Add0~29 )) # (!\rdat1[15]~21_combout  & ((!\Add0~29 ) # (!\port_b~63_combout ))))

	.dataa(rdat1_15),
	.datab(port_b53),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~29 ),
	.combout(\Add0~30_combout ),
	.cout(\Add0~31 ));
// synopsys translate_off
defparam \Add0~30 .lut_mask = 16'h9617;
defparam \Add0~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N0
cycloneive_lcell_comb \Add0~32 (
// Equation(s):
// \Add0~32_combout  = ((\rdat1[16]~19_combout  $ (\port_b~22_combout  $ (!\Add0~31 )))) # (GND)
// \Add0~33  = CARRY((\rdat1[16]~19_combout  & ((\port_b~22_combout ) # (!\Add0~31 ))) # (!\rdat1[16]~19_combout  & (\port_b~22_combout  & !\Add0~31 )))

	.dataa(rdat1_16),
	.datab(port_b12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~31 ),
	.combout(\Add0~32_combout ),
	.cout(\Add0~33 ));
// synopsys translate_off
defparam \Add0~32 .lut_mask = 16'h698E;
defparam \Add0~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N2
cycloneive_lcell_comb \Add0~34 (
// Equation(s):
// \Add0~34_combout  = (\rdat1[17]~63_combout  & ((\port_b~24_combout  & (\Add0~33  & VCC)) # (!\port_b~24_combout  & (!\Add0~33 )))) # (!\rdat1[17]~63_combout  & ((\port_b~24_combout  & (!\Add0~33 )) # (!\port_b~24_combout  & ((\Add0~33 ) # (GND)))))
// \Add0~35  = CARRY((\rdat1[17]~63_combout  & (!\port_b~24_combout  & !\Add0~33 )) # (!\rdat1[17]~63_combout  & ((!\Add0~33 ) # (!\port_b~24_combout ))))

	.dataa(rdat1_17),
	.datab(port_b14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~33 ),
	.combout(\Add0~34_combout ),
	.cout(\Add0~35 ));
// synopsys translate_off
defparam \Add0~34 .lut_mask = 16'h9617;
defparam \Add0~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N4
cycloneive_lcell_comb \Add0~36 (
// Equation(s):
// \Add0~36_combout  = ((\rdat1[18]~59_combout  $ (\port_b~26_combout  $ (!\Add0~35 )))) # (GND)
// \Add0~37  = CARRY((\rdat1[18]~59_combout  & ((\port_b~26_combout ) # (!\Add0~35 ))) # (!\rdat1[18]~59_combout  & (\port_b~26_combout  & !\Add0~35 )))

	.dataa(rdat1_18),
	.datab(port_b16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~35 ),
	.combout(\Add0~36_combout ),
	.cout(\Add0~37 ));
// synopsys translate_off
defparam \Add0~36 .lut_mask = 16'h698E;
defparam \Add0~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N6
cycloneive_lcell_comb \Add0~38 (
// Equation(s):
// \Add0~38_combout  = (\rdat1[19]~61_combout  & ((\port_b~28_combout  & (\Add0~37  & VCC)) # (!\port_b~28_combout  & (!\Add0~37 )))) # (!\rdat1[19]~61_combout  & ((\port_b~28_combout  & (!\Add0~37 )) # (!\port_b~28_combout  & ((\Add0~37 ) # (GND)))))
// \Add0~39  = CARRY((\rdat1[19]~61_combout  & (!\port_b~28_combout  & !\Add0~37 )) # (!\rdat1[19]~61_combout  & ((!\Add0~37 ) # (!\port_b~28_combout ))))

	.dataa(rdat1_19),
	.datab(port_b18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~37 ),
	.combout(\Add0~38_combout ),
	.cout(\Add0~39 ));
// synopsys translate_off
defparam \Add0~38 .lut_mask = 16'h9617;
defparam \Add0~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N8
cycloneive_lcell_comb \Add0~40 (
// Equation(s):
// \Add0~40_combout  = ((\rdat1[20]~57_combout  $ (\port_b~30_combout  $ (!\Add0~39 )))) # (GND)
// \Add0~41  = CARRY((\rdat1[20]~57_combout  & ((\port_b~30_combout ) # (!\Add0~39 ))) # (!\rdat1[20]~57_combout  & (\port_b~30_combout  & !\Add0~39 )))

	.dataa(rdat1_20),
	.datab(port_b20),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~39 ),
	.combout(\Add0~40_combout ),
	.cout(\Add0~41 ));
// synopsys translate_off
defparam \Add0~40 .lut_mask = 16'h698E;
defparam \Add0~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N10
cycloneive_lcell_comb \Add0~42 (
// Equation(s):
// \Add0~42_combout  = (\rdat1[21]~55_combout  & ((\port_b~32_combout  & (\Add0~41  & VCC)) # (!\port_b~32_combout  & (!\Add0~41 )))) # (!\rdat1[21]~55_combout  & ((\port_b~32_combout  & (!\Add0~41 )) # (!\port_b~32_combout  & ((\Add0~41 ) # (GND)))))
// \Add0~43  = CARRY((\rdat1[21]~55_combout  & (!\port_b~32_combout  & !\Add0~41 )) # (!\rdat1[21]~55_combout  & ((!\Add0~41 ) # (!\port_b~32_combout ))))

	.dataa(rdat1_21),
	.datab(port_b22),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~41 ),
	.combout(\Add0~42_combout ),
	.cout(\Add0~43 ));
// synopsys translate_off
defparam \Add0~42 .lut_mask = 16'h9617;
defparam \Add0~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N12
cycloneive_lcell_comb \Add0~44 (
// Equation(s):
// \Add0~44_combout  = ((\rdat1[22]~51_combout  $ (\port_b~34_combout  $ (!\Add0~43 )))) # (GND)
// \Add0~45  = CARRY((\rdat1[22]~51_combout  & ((\port_b~34_combout ) # (!\Add0~43 ))) # (!\rdat1[22]~51_combout  & (\port_b~34_combout  & !\Add0~43 )))

	.dataa(rdat1_22),
	.datab(port_b24),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~43 ),
	.combout(\Add0~44_combout ),
	.cout(\Add0~45 ));
// synopsys translate_off
defparam \Add0~44 .lut_mask = 16'h698E;
defparam \Add0~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N16
cycloneive_lcell_comb \Add0~48 (
// Equation(s):
// \Add0~48_combout  = ((\rdat1[24]~49_combout  $ (\port_b~38_combout  $ (!\Add0~47 )))) # (GND)
// \Add0~49  = CARRY((\rdat1[24]~49_combout  & ((\port_b~38_combout ) # (!\Add0~47 ))) # (!\rdat1[24]~49_combout  & (\port_b~38_combout  & !\Add0~47 )))

	.dataa(rdat1_24),
	.datab(port_b28),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~47 ),
	.combout(\Add0~48_combout ),
	.cout(\Add0~49 ));
// synopsys translate_off
defparam \Add0~48 .lut_mask = 16'h698E;
defparam \Add0~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N10
cycloneive_lcell_comb \out~12 (
// Equation(s):
// \out~12_combout  = \rdat1[24]~49_combout  $ (((\port_b~37_combout ) # ((\port_b~0_combout  & fuifrtReplace_24))))

	.dataa(port_b),
	.datab(port_b27),
	.datac(fuifrtReplace_24),
	.datad(rdat1_24),
	.cin(gnd),
	.combout(\out~12_combout ),
	.cout());
// synopsys translate_off
defparam \out~12 .lut_mask = 16'h13EC;
defparam \out~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N8
cycloneive_lcell_comb \ShiftLeft0~34 (
// Equation(s):
// \ShiftLeft0~34_combout  = (!\port_b~7_combout  & ((\port_b~4_combout  & (\rdat1[22]~51_combout )) # (!\port_b~4_combout  & ((\rdat1[24]~49_combout )))))

	.dataa(rdat1_22),
	.datab(port_b4),
	.datac(port_b2),
	.datad(rdat1_24),
	.cin(gnd),
	.combout(\ShiftLeft0~34_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~34 .lut_mask = 16'h2320;
defparam \ShiftLeft0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N18
cycloneive_lcell_comb \ShiftLeft0~35 (
// Equation(s):
// \ShiftLeft0~35_combout  = (\port_b~4_combout  & ((\rdat1[21]~55_combout ))) # (!\port_b~4_combout  & (\rdat1[23]~53_combout ))

	.dataa(gnd),
	.datab(rdat1_23),
	.datac(port_b2),
	.datad(rdat1_21),
	.cin(gnd),
	.combout(\ShiftLeft0~35_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~35 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N24
cycloneive_lcell_comb \ShiftLeft0~36 (
// Equation(s):
// \ShiftLeft0~36_combout  = (\ShiftLeft0~34_combout ) # ((\port_b~7_combout  & \ShiftLeft0~35_combout ))

	.dataa(gnd),
	.datab(port_b4),
	.datac(\ShiftLeft0~34_combout ),
	.datad(\ShiftLeft0~35_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~36_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~36 .lut_mask = 16'hFCF0;
defparam \ShiftLeft0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N22
cycloneive_lcell_comb \myif.out[24]~36 (
// Equation(s):
// \myif.out[24]~36_combout  = (\myif.out[5]~17_combout  & ((\ShiftLeft0~33_combout ) # ((\myif.out[5]~16_combout )))) # (!\myif.out[5]~17_combout  & (((\ShiftLeft0~36_combout  & !\myif.out[5]~16_combout ))))

	.dataa(\ShiftLeft0~33_combout ),
	.datab(\ShiftLeft0~36_combout ),
	.datac(\myif.out[5]~17_combout ),
	.datad(\myif.out[5]~16_combout ),
	.cin(gnd),
	.combout(\myif.out[24]~36_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[24]~36 .lut_mask = 16'hF0AC;
defparam \myif.out[24]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N0
cycloneive_lcell_comb \ShiftLeft0~25 (
// Equation(s):
// \ShiftLeft0~25_combout  = (\port_b~7_combout  & ((\rdat1[9]~33_combout ))) # (!\port_b~7_combout  & (\rdat1[10]~31_combout ))

	.dataa(port_b4),
	.datab(gnd),
	.datac(rdat1_10),
	.datad(rdat1_9),
	.cin(gnd),
	.combout(\ShiftLeft0~25_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~25 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N16
cycloneive_lcell_comb \ShiftLeft0~26 (
// Equation(s):
// \ShiftLeft0~26_combout  = (\port_b~7_combout  & ((\rdat1[11]~29_combout ))) # (!\port_b~7_combout  & (\rdat1[12]~27_combout ))

	.dataa(port_b4),
	.datab(gnd),
	.datac(rdat1_12),
	.datad(rdat1_11),
	.cin(gnd),
	.combout(\ShiftLeft0~26_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~26 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N18
cycloneive_lcell_comb \ShiftLeft0~27 (
// Equation(s):
// \ShiftLeft0~27_combout  = (\port_b~4_combout  & (\ShiftLeft0~25_combout )) # (!\port_b~4_combout  & ((\ShiftLeft0~26_combout )))

	.dataa(port_b2),
	.datab(gnd),
	.datac(\ShiftLeft0~25_combout ),
	.datad(\ShiftLeft0~26_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~27_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~27 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N26
cycloneive_lcell_comb \ShiftLeft0~28 (
// Equation(s):
// \ShiftLeft0~28_combout  = (\port_b~7_combout  & ((\port_b~4_combout  & ((\rdat1[13]~25_combout ))) # (!\port_b~4_combout  & (\rdat1[15]~21_combout ))))

	.dataa(port_b2),
	.datab(port_b4),
	.datac(rdat1_15),
	.datad(rdat1_13),
	.cin(gnd),
	.combout(\ShiftLeft0~28_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~28 .lut_mask = 16'hC840;
defparam \ShiftLeft0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N8
cycloneive_lcell_comb \ShiftLeft0~30 (
// Equation(s):
// \ShiftLeft0~30_combout  = (\port_b~10_combout  & (((\ShiftLeft0~27_combout )))) # (!\port_b~10_combout  & ((\ShiftLeft0~29_combout ) # ((\ShiftLeft0~28_combout ))))

	.dataa(\ShiftLeft0~29_combout ),
	.datab(port_b6),
	.datac(\ShiftLeft0~27_combout ),
	.datad(\ShiftLeft0~28_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~30_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~30 .lut_mask = 16'hF3E2;
defparam \ShiftLeft0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N14
cycloneive_lcell_comb \ShiftLeft0~37 (
// Equation(s):
// \ShiftLeft0~37_combout  = (\port_b~7_combout  & (\rdat1[7]~13_combout )) # (!\port_b~7_combout  & ((\rdat1[8]~11_combout )))

	.dataa(rdat1_7),
	.datab(gnd),
	.datac(rdat1_8),
	.datad(port_b4),
	.cin(gnd),
	.combout(\ShiftLeft0~37_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~37 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N2
cycloneive_lcell_comb \ShiftLeft0~38 (
// Equation(s):
// \ShiftLeft0~38_combout  = (\port_b~4_combout  & (\ShiftLeft0~18_combout )) # (!\port_b~4_combout  & ((\ShiftLeft0~37_combout )))

	.dataa(port_b2),
	.datab(gnd),
	.datac(\ShiftLeft0~18_combout ),
	.datad(\ShiftLeft0~37_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~38_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~38 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N16
cycloneive_lcell_comb \ShiftLeft0~39 (
// Equation(s):
// \ShiftLeft0~39_combout  = (\port_b~10_combout  & (\ShiftLeft0~23_combout )) # (!\port_b~10_combout  & ((\ShiftLeft0~38_combout )))

	.dataa(gnd),
	.datab(port_b6),
	.datac(\ShiftLeft0~23_combout ),
	.datad(\ShiftLeft0~38_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~39_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~39 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N6
cycloneive_lcell_comb \ShiftLeft0~40 (
// Equation(s):
// \ShiftLeft0~40_combout  = (\port_b~14_combout  & (!\port_b~10_combout  & (\ShiftLeft0~21_combout ))) # (!\port_b~14_combout  & (((\ShiftLeft0~39_combout ))))

	.dataa(port_b6),
	.datab(\ShiftLeft0~21_combout ),
	.datac(port_b7),
	.datad(\ShiftLeft0~39_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~40_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~40 .lut_mask = 16'h4F40;
defparam \ShiftLeft0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N18
cycloneive_lcell_comb \myif.out[24]~37 (
// Equation(s):
// \myif.out[24]~37_combout  = (\myif.out[5]~16_combout  & ((\myif.out[24]~36_combout  & ((\ShiftLeft0~40_combout ))) # (!\myif.out[24]~36_combout  & (\ShiftLeft0~30_combout )))) # (!\myif.out[5]~16_combout  & (\myif.out[24]~36_combout ))

	.dataa(\myif.out[5]~16_combout ),
	.datab(\myif.out[24]~36_combout ),
	.datac(\ShiftLeft0~30_combout ),
	.datad(\ShiftLeft0~40_combout ),
	.cin(gnd),
	.combout(\myif.out[24]~37_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[24]~37 .lut_mask = 16'hEC64;
defparam \myif.out[24]~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N24
cycloneive_lcell_comb \myif.out[24]~38 (
// Equation(s):
// \myif.out[24]~38_combout  = (idex_ifaluop_o_2 & ((\out~13_combout ) # ((!\myif.out[5]~20_combout )))) # (!idex_ifaluop_o_2 & (((\myif.out[5]~20_combout  & \myif.out[24]~37_combout ))))

	.dataa(\out~13_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\myif.out[5]~20_combout ),
	.datad(\myif.out[24]~37_combout ),
	.cin(gnd),
	.combout(\myif.out[24]~38_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[24]~38 .lut_mask = 16'hBC8C;
defparam \myif.out[24]~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N22
cycloneive_lcell_comb \myif.out[24]~39 (
// Equation(s):
// \myif.out[24]~39_combout  = (idex_ifaluop_o_1 & ((\myif.out[24]~38_combout  & ((\out~12_combout ))) # (!\myif.out[24]~38_combout  & (\Add0~48_combout )))) # (!idex_ifaluop_o_1 & (((\myif.out[24]~38_combout ))))

	.dataa(\Add0~48_combout ),
	.datab(\out~12_combout ),
	.datac(idex_ifaluop_o_1),
	.datad(\myif.out[24]~38_combout ),
	.cin(gnd),
	.combout(\myif.out[24]~39_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[24]~39 .lut_mask = 16'hCFA0;
defparam \myif.out[24]~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N12
cycloneive_lcell_comb \out~11 (
// Equation(s):
// \out~11_combout  = (\port_b~37_combout ) # ((\rdat1[24]~49_combout ) # ((\port_b~0_combout  & fuifrtReplace_24)))

	.dataa(port_b),
	.datab(port_b27),
	.datac(fuifrtReplace_24),
	.datad(rdat1_24),
	.cin(gnd),
	.combout(\out~11_combout ),
	.cout());
// synopsys translate_off
defparam \out~11 .lut_mask = 16'hFFEC;
defparam \out~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N14
cycloneive_lcell_comb \Add1~14 (
// Equation(s):
// \Add1~14_combout  = (\rdat1[7]~13_combout  & ((\port_b~48_combout  & (!\Add1~13 )) # (!\port_b~48_combout  & (\Add1~13  & VCC)))) # (!\rdat1[7]~13_combout  & ((\port_b~48_combout  & ((\Add1~13 ) # (GND))) # (!\port_b~48_combout  & (!\Add1~13 ))))
// \Add1~15  = CARRY((\rdat1[7]~13_combout  & (\port_b~48_combout  & !\Add1~13 )) # (!\rdat1[7]~13_combout  & ((\port_b~48_combout ) # (!\Add1~13 ))))

	.dataa(rdat1_7),
	.datab(port_b38),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~13 ),
	.combout(\Add1~14_combout ),
	.cout(\Add1~15 ));
// synopsys translate_off
defparam \Add1~14 .lut_mask = 16'h694D;
defparam \Add1~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N16
cycloneive_lcell_comb \Add1~16 (
// Equation(s):
// \Add1~16_combout  = ((\rdat1[8]~11_combout  $ (\port_b~50_combout  $ (\Add1~15 )))) # (GND)
// \Add1~17  = CARRY((\rdat1[8]~11_combout  & ((!\Add1~15 ) # (!\port_b~50_combout ))) # (!\rdat1[8]~11_combout  & (!\port_b~50_combout  & !\Add1~15 )))

	.dataa(rdat1_8),
	.datab(port_b40),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~15 ),
	.combout(\Add1~16_combout ),
	.cout(\Add1~17 ));
// synopsys translate_off
defparam \Add1~16 .lut_mask = 16'h962B;
defparam \Add1~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N18
cycloneive_lcell_comb \Add1~18 (
// Equation(s):
// \Add1~18_combout  = (\rdat1[9]~33_combout  & ((\port_b~60_combout  & (!\Add1~17 )) # (!\port_b~60_combout  & (\Add1~17  & VCC)))) # (!\rdat1[9]~33_combout  & ((\port_b~60_combout  & ((\Add1~17 ) # (GND))) # (!\port_b~60_combout  & (!\Add1~17 ))))
// \Add1~19  = CARRY((\rdat1[9]~33_combout  & (\port_b~60_combout  & !\Add1~17 )) # (!\rdat1[9]~33_combout  & ((\port_b~60_combout ) # (!\Add1~17 ))))

	.dataa(rdat1_9),
	.datab(port_b50),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~17 ),
	.combout(\Add1~18_combout ),
	.cout(\Add1~19 ));
// synopsys translate_off
defparam \Add1~18 .lut_mask = 16'h694D;
defparam \Add1~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N20
cycloneive_lcell_comb \Add1~20 (
// Equation(s):
// \Add1~20_combout  = ((\port_b~65_combout  $ (\rdat1[10]~31_combout  $ (\Add1~19 )))) # (GND)
// \Add1~21  = CARRY((\port_b~65_combout  & (\rdat1[10]~31_combout  & !\Add1~19 )) # (!\port_b~65_combout  & ((\rdat1[10]~31_combout ) # (!\Add1~19 ))))

	.dataa(port_b55),
	.datab(rdat1_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~19 ),
	.combout(\Add1~20_combout ),
	.cout(\Add1~21 ));
// synopsys translate_off
defparam \Add1~20 .lut_mask = 16'h964D;
defparam \Add1~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N22
cycloneive_lcell_comb \Add1~22 (
// Equation(s):
// \Add1~22_combout  = (\port_b~67_combout  & ((\rdat1[11]~29_combout  & (!\Add1~21 )) # (!\rdat1[11]~29_combout  & ((\Add1~21 ) # (GND))))) # (!\port_b~67_combout  & ((\rdat1[11]~29_combout  & (\Add1~21  & VCC)) # (!\rdat1[11]~29_combout  & (!\Add1~21 ))))
// \Add1~23  = CARRY((\port_b~67_combout  & ((!\Add1~21 ) # (!\rdat1[11]~29_combout ))) # (!\port_b~67_combout  & (!\rdat1[11]~29_combout  & !\Add1~21 )))

	.dataa(port_b57),
	.datab(rdat1_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~21 ),
	.combout(\Add1~22_combout ),
	.cout(\Add1~23 ));
// synopsys translate_off
defparam \Add1~22 .lut_mask = 16'h692B;
defparam \Add1~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N24
cycloneive_lcell_comb \Add1~24 (
// Equation(s):
// \Add1~24_combout  = ((\port_b~72_combout  $ (\rdat1[12]~27_combout  $ (\Add1~23 )))) # (GND)
// \Add1~25  = CARRY((\port_b~72_combout  & (\rdat1[12]~27_combout  & !\Add1~23 )) # (!\port_b~72_combout  & ((\rdat1[12]~27_combout ) # (!\Add1~23 ))))

	.dataa(port_b62),
	.datab(rdat1_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~23 ),
	.combout(\Add1~24_combout ),
	.cout(\Add1~25 ));
// synopsys translate_off
defparam \Add1~24 .lut_mask = 16'h964D;
defparam \Add1~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N26
cycloneive_lcell_comb \Add1~26 (
// Equation(s):
// \Add1~26_combout  = (\rdat1[13]~25_combout  & ((\port_b~70_combout  & (!\Add1~25 )) # (!\port_b~70_combout  & (\Add1~25  & VCC)))) # (!\rdat1[13]~25_combout  & ((\port_b~70_combout  & ((\Add1~25 ) # (GND))) # (!\port_b~70_combout  & (!\Add1~25 ))))
// \Add1~27  = CARRY((\rdat1[13]~25_combout  & (\port_b~70_combout  & !\Add1~25 )) # (!\rdat1[13]~25_combout  & ((\port_b~70_combout ) # (!\Add1~25 ))))

	.dataa(rdat1_13),
	.datab(port_b60),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~25 ),
	.combout(\Add1~26_combout ),
	.cout(\Add1~27 ));
// synopsys translate_off
defparam \Add1~26 .lut_mask = 16'h694D;
defparam \Add1~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N28
cycloneive_lcell_comb \Add1~28 (
// Equation(s):
// \Add1~28_combout  = ((\rdat1[14]~23_combout  $ (\port_b~71_combout  $ (\Add1~27 )))) # (GND)
// \Add1~29  = CARRY((\rdat1[14]~23_combout  & ((!\Add1~27 ) # (!\port_b~71_combout ))) # (!\rdat1[14]~23_combout  & (!\port_b~71_combout  & !\Add1~27 )))

	.dataa(rdat1_14),
	.datab(port_b61),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~27 ),
	.combout(\Add1~28_combout ),
	.cout(\Add1~29 ));
// synopsys translate_off
defparam \Add1~28 .lut_mask = 16'h962B;
defparam \Add1~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N30
cycloneive_lcell_comb \Add1~30 (
// Equation(s):
// \Add1~30_combout  = (\port_b~63_combout  & ((\rdat1[15]~21_combout  & (!\Add1~29 )) # (!\rdat1[15]~21_combout  & ((\Add1~29 ) # (GND))))) # (!\port_b~63_combout  & ((\rdat1[15]~21_combout  & (\Add1~29  & VCC)) # (!\rdat1[15]~21_combout  & (!\Add1~29 ))))
// \Add1~31  = CARRY((\port_b~63_combout  & ((!\Add1~29 ) # (!\rdat1[15]~21_combout ))) # (!\port_b~63_combout  & (!\rdat1[15]~21_combout  & !\Add1~29 )))

	.dataa(port_b53),
	.datab(rdat1_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~29 ),
	.combout(\Add1~30_combout ),
	.cout(\Add1~31 ));
// synopsys translate_off
defparam \Add1~30 .lut_mask = 16'h692B;
defparam \Add1~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N2
cycloneive_lcell_comb \Add1~34 (
// Equation(s):
// \Add1~34_combout  = (\port_b~24_combout  & ((\rdat1[17]~63_combout  & (!\Add1~33 )) # (!\rdat1[17]~63_combout  & ((\Add1~33 ) # (GND))))) # (!\port_b~24_combout  & ((\rdat1[17]~63_combout  & (\Add1~33  & VCC)) # (!\rdat1[17]~63_combout  & (!\Add1~33 ))))
// \Add1~35  = CARRY((\port_b~24_combout  & ((!\Add1~33 ) # (!\rdat1[17]~63_combout ))) # (!\port_b~24_combout  & (!\rdat1[17]~63_combout  & !\Add1~33 )))

	.dataa(port_b14),
	.datab(rdat1_17),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~33 ),
	.combout(\Add1~34_combout ),
	.cout(\Add1~35 ));
// synopsys translate_off
defparam \Add1~34 .lut_mask = 16'h692B;
defparam \Add1~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N4
cycloneive_lcell_comb \Add1~36 (
// Equation(s):
// \Add1~36_combout  = ((\port_b~26_combout  $ (\rdat1[18]~59_combout  $ (\Add1~35 )))) # (GND)
// \Add1~37  = CARRY((\port_b~26_combout  & (\rdat1[18]~59_combout  & !\Add1~35 )) # (!\port_b~26_combout  & ((\rdat1[18]~59_combout ) # (!\Add1~35 ))))

	.dataa(port_b16),
	.datab(rdat1_18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~35 ),
	.combout(\Add1~36_combout ),
	.cout(\Add1~37 ));
// synopsys translate_off
defparam \Add1~36 .lut_mask = 16'h964D;
defparam \Add1~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N6
cycloneive_lcell_comb \Add1~38 (
// Equation(s):
// \Add1~38_combout  = (\rdat1[19]~61_combout  & ((\port_b~28_combout  & (!\Add1~37 )) # (!\port_b~28_combout  & (\Add1~37  & VCC)))) # (!\rdat1[19]~61_combout  & ((\port_b~28_combout  & ((\Add1~37 ) # (GND))) # (!\port_b~28_combout  & (!\Add1~37 ))))
// \Add1~39  = CARRY((\rdat1[19]~61_combout  & (\port_b~28_combout  & !\Add1~37 )) # (!\rdat1[19]~61_combout  & ((\port_b~28_combout ) # (!\Add1~37 ))))

	.dataa(rdat1_19),
	.datab(port_b18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~37 ),
	.combout(\Add1~38_combout ),
	.cout(\Add1~39 ));
// synopsys translate_off
defparam \Add1~38 .lut_mask = 16'h694D;
defparam \Add1~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N8
cycloneive_lcell_comb \Add1~40 (
// Equation(s):
// \Add1~40_combout  = ((\rdat1[20]~57_combout  $ (\port_b~30_combout  $ (\Add1~39 )))) # (GND)
// \Add1~41  = CARRY((\rdat1[20]~57_combout  & ((!\Add1~39 ) # (!\port_b~30_combout ))) # (!\rdat1[20]~57_combout  & (!\port_b~30_combout  & !\Add1~39 )))

	.dataa(rdat1_20),
	.datab(port_b20),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~39 ),
	.combout(\Add1~40_combout ),
	.cout(\Add1~41 ));
// synopsys translate_off
defparam \Add1~40 .lut_mask = 16'h962B;
defparam \Add1~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N10
cycloneive_lcell_comb \Add1~42 (
// Equation(s):
// \Add1~42_combout  = (\rdat1[21]~55_combout  & ((\port_b~32_combout  & (!\Add1~41 )) # (!\port_b~32_combout  & (\Add1~41  & VCC)))) # (!\rdat1[21]~55_combout  & ((\port_b~32_combout  & ((\Add1~41 ) # (GND))) # (!\port_b~32_combout  & (!\Add1~41 ))))
// \Add1~43  = CARRY((\rdat1[21]~55_combout  & (\port_b~32_combout  & !\Add1~41 )) # (!\rdat1[21]~55_combout  & ((\port_b~32_combout ) # (!\Add1~41 ))))

	.dataa(rdat1_21),
	.datab(port_b22),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~41 ),
	.combout(\Add1~42_combout ),
	.cout(\Add1~43 ));
// synopsys translate_off
defparam \Add1~42 .lut_mask = 16'h694D;
defparam \Add1~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N12
cycloneive_lcell_comb \Add1~44 (
// Equation(s):
// \Add1~44_combout  = ((\rdat1[22]~51_combout  $ (\port_b~34_combout  $ (\Add1~43 )))) # (GND)
// \Add1~45  = CARRY((\rdat1[22]~51_combout  & ((!\Add1~43 ) # (!\port_b~34_combout ))) # (!\rdat1[22]~51_combout  & (!\port_b~34_combout  & !\Add1~43 )))

	.dataa(rdat1_22),
	.datab(port_b24),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~43 ),
	.combout(\Add1~44_combout ),
	.cout(\Add1~45 ));
// synopsys translate_off
defparam \Add1~44 .lut_mask = 16'h962B;
defparam \Add1~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N14
cycloneive_lcell_comb \Add1~46 (
// Equation(s):
// \Add1~46_combout  = (\rdat1[23]~53_combout  & ((\port_b~36_combout  & (!\Add1~45 )) # (!\port_b~36_combout  & (\Add1~45  & VCC)))) # (!\rdat1[23]~53_combout  & ((\port_b~36_combout  & ((\Add1~45 ) # (GND))) # (!\port_b~36_combout  & (!\Add1~45 ))))
// \Add1~47  = CARRY((\rdat1[23]~53_combout  & (\port_b~36_combout  & !\Add1~45 )) # (!\rdat1[23]~53_combout  & ((\port_b~36_combout ) # (!\Add1~45 ))))

	.dataa(rdat1_23),
	.datab(port_b26),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~45 ),
	.combout(\Add1~46_combout ),
	.cout(\Add1~47 ));
// synopsys translate_off
defparam \Add1~46 .lut_mask = 16'h694D;
defparam \Add1~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N16
cycloneive_lcell_comb \Add1~48 (
// Equation(s):
// \Add1~48_combout  = ((\port_b~38_combout  $ (\rdat1[24]~49_combout  $ (\Add1~47 )))) # (GND)
// \Add1~49  = CARRY((\port_b~38_combout  & (\rdat1[24]~49_combout  & !\Add1~47 )) # (!\port_b~38_combout  & ((\rdat1[24]~49_combout ) # (!\Add1~47 ))))

	.dataa(port_b28),
	.datab(rdat1_24),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~47 ),
	.combout(\Add1~48_combout ),
	.cout(\Add1~49 ));
// synopsys translate_off
defparam \Add1~48 .lut_mask = 16'h964D;
defparam \Add1~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N22
cycloneive_lcell_comb \ShiftRight0~52 (
// Equation(s):
// \ShiftRight0~52_combout  = (\port_b~7_combout  & ((\rdat1[31]~35_combout ))) # (!\port_b~7_combout  & (\rdat1[30]~39_combout ))

	.dataa(port_b4),
	.datab(rdat1_30),
	.datac(gnd),
	.datad(rdat1_311),
	.cin(gnd),
	.combout(\ShiftRight0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~52 .lut_mask = 16'hEE44;
defparam \ShiftRight0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N2
cycloneive_lcell_comb \ShiftRight0~67 (
// Equation(s):
// \ShiftRight0~67_combout  = (\ShiftRight0~66_combout ) # ((\port_b~4_combout  & \ShiftRight0~52_combout ))

	.dataa(\ShiftRight0~66_combout ),
	.datab(port_b2),
	.datac(\ShiftRight0~52_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~67 .lut_mask = 16'hEAEA;
defparam \ShiftRight0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N24
cycloneive_lcell_comb \ShiftRight0~69 (
// Equation(s):
// \ShiftRight0~69_combout  = (!\port_b~14_combout  & ((\port_b~10_combout  & ((\ShiftRight0~67_combout ))) # (!\port_b~10_combout  & (\ShiftRight0~62_combout ))))

	.dataa(port_b7),
	.datab(\ShiftRight0~62_combout ),
	.datac(port_b6),
	.datad(\ShiftRight0~67_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~69 .lut_mask = 16'h5404;
defparam \ShiftRight0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N2
cycloneive_lcell_comb \myif.out[24]~34 (
// Equation(s):
// \myif.out[24]~34_combout  = (idex_ifaluop_o_2 & ((\out~11_combout ) # ((!\myif.out[13]~23_combout )))) # (!idex_ifaluop_o_2 & (((\ShiftRight0~69_combout  & \myif.out[13]~23_combout ))))

	.dataa(\out~11_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\ShiftRight0~69_combout ),
	.datad(\myif.out[13]~23_combout ),
	.cin(gnd),
	.combout(\myif.out[24]~34_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[24]~34 .lut_mask = 16'hB8CC;
defparam \myif.out[24]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N0
cycloneive_lcell_comb \myif.out[24]~35 (
// Equation(s):
// \myif.out[24]~35_combout  = (idex_ifaluop_o_1 & ((\myif.out[24]~34_combout  & (!\out~11_combout )) # (!\myif.out[24]~34_combout  & ((\Add1~48_combout ))))) # (!idex_ifaluop_o_1 & (((\myif.out[24]~34_combout ))))

	.dataa(\out~11_combout ),
	.datab(idex_ifaluop_o_1),
	.datac(\Add1~48_combout ),
	.datad(\myif.out[24]~34_combout ),
	.cin(gnd),
	.combout(\myif.out[24]~35_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[24]~35 .lut_mask = 16'h77C0;
defparam \myif.out[24]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N2
cycloneive_lcell_comb \out~14 (
// Equation(s):
// \out~14_combout  = (\port_b~41_combout ) # ((\rdat1[26]~43_combout ) # ((fuifrtReplace_26 & \port_b~0_combout )))

	.dataa(fuifrtReplace_26),
	.datab(port_b),
	.datac(port_b31),
	.datad(rdat1_26),
	.cin(gnd),
	.combout(\out~14_combout ),
	.cout());
// synopsys translate_off
defparam \out~14 .lut_mask = 16'hFFF8;
defparam \out~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N0
cycloneive_lcell_comb \ShiftRight0~70 (
// Equation(s):
// \ShiftRight0~70_combout  = (\port_b~10_combout  & (!\port_b~4_combout  & ((\ShiftRight0~52_combout )))) # (!\port_b~10_combout  & (((\ShiftRight0~47_combout ))))

	.dataa(port_b2),
	.datab(port_b6),
	.datac(\ShiftRight0~47_combout ),
	.datad(\ShiftRight0~52_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~70 .lut_mask = 16'h7430;
defparam \ShiftRight0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N30
cycloneive_lcell_comb \ShiftRight0~71 (
// Equation(s):
// \ShiftRight0~71_combout  = (!\port_b~14_combout  & \ShiftRight0~70_combout )

	.dataa(gnd),
	.datab(port_b7),
	.datac(gnd),
	.datad(\ShiftRight0~70_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~71 .lut_mask = 16'h3300;
defparam \ShiftRight0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N4
cycloneive_lcell_comb \myif.out[26]~41 (
// Equation(s):
// \myif.out[26]~41_combout  = (idex_ifaluop_o_2 & ((\out~14_combout ) # ((!\myif.out[13]~23_combout )))) # (!idex_ifaluop_o_2 & (((\ShiftRight0~71_combout  & \myif.out[13]~23_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\out~14_combout ),
	.datac(\ShiftRight0~71_combout ),
	.datad(\myif.out[13]~23_combout ),
	.cin(gnd),
	.combout(\myif.out[26]~41_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[26]~41 .lut_mask = 16'hD8AA;
defparam \myif.out[26]~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N18
cycloneive_lcell_comb \Add1~50 (
// Equation(s):
// \Add1~50_combout  = (\port_b~40_combout  & ((\rdat1[25]~47_combout  & (!\Add1~49 )) # (!\rdat1[25]~47_combout  & ((\Add1~49 ) # (GND))))) # (!\port_b~40_combout  & ((\rdat1[25]~47_combout  & (\Add1~49  & VCC)) # (!\rdat1[25]~47_combout  & (!\Add1~49 ))))
// \Add1~51  = CARRY((\port_b~40_combout  & ((!\Add1~49 ) # (!\rdat1[25]~47_combout ))) # (!\port_b~40_combout  & (!\rdat1[25]~47_combout  & !\Add1~49 )))

	.dataa(port_b30),
	.datab(rdat1_25),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~49 ),
	.combout(\Add1~50_combout ),
	.cout(\Add1~51 ));
// synopsys translate_off
defparam \Add1~50 .lut_mask = 16'h692B;
defparam \Add1~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N20
cycloneive_lcell_comb \Add1~52 (
// Equation(s):
// \Add1~52_combout  = ((\rdat1[26]~43_combout  $ (\port_b~42_combout  $ (\Add1~51 )))) # (GND)
// \Add1~53  = CARRY((\rdat1[26]~43_combout  & ((!\Add1~51 ) # (!\port_b~42_combout ))) # (!\rdat1[26]~43_combout  & (!\port_b~42_combout  & !\Add1~51 )))

	.dataa(rdat1_26),
	.datab(port_b32),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~51 ),
	.combout(\Add1~52_combout ),
	.cout(\Add1~53 ));
// synopsys translate_off
defparam \Add1~52 .lut_mask = 16'h962B;
defparam \Add1~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N26
cycloneive_lcell_comb \myif.out[26]~42 (
// Equation(s):
// \myif.out[26]~42_combout  = (idex_ifaluop_o_1 & ((\myif.out[26]~41_combout  & (!\out~14_combout )) # (!\myif.out[26]~41_combout  & ((\Add1~52_combout ))))) # (!idex_ifaluop_o_1 & (((\myif.out[26]~41_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(\out~14_combout ),
	.datac(\myif.out[26]~41_combout ),
	.datad(\Add1~52_combout ),
	.cin(gnd),
	.combout(\myif.out[26]~42_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[26]~42 .lut_mask = 16'h7A70;
defparam \myif.out[26]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N30
cycloneive_lcell_comb \out~15 (
// Equation(s):
// \out~15_combout  = \rdat1[26]~43_combout  $ (((\port_b~41_combout ) # ((\port_b~0_combout  & fuifrtReplace_26))))

	.dataa(rdat1_26),
	.datab(port_b),
	.datac(port_b31),
	.datad(fuifrtReplace_26),
	.cin(gnd),
	.combout(\out~15_combout ),
	.cout());
// synopsys translate_off
defparam \out~15 .lut_mask = 16'h565A;
defparam \out~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N28
cycloneive_lcell_comb \out~16 (
// Equation(s):
// \out~16_combout  = (\rdat1[26]~43_combout  & ((\port_b~41_combout ) # ((fuifrtReplace_26 & \port_b~0_combout ))))

	.dataa(fuifrtReplace_26),
	.datab(rdat1_26),
	.datac(port_b31),
	.datad(port_b),
	.cin(gnd),
	.combout(\out~16_combout ),
	.cout());
// synopsys translate_off
defparam \out~16 .lut_mask = 16'hC8C0;
defparam \out~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N8
cycloneive_lcell_comb \ShiftLeft0~15 (
// Equation(s):
// \ShiftLeft0~15_combout  = (!\port_b~7_combout  & ((\port_b~4_combout  & (\rdat1[0]~3_combout )) # (!\port_b~4_combout  & ((\rdat1[2]~5_combout )))))

	.dataa(rdat1_0),
	.datab(rdat1_2),
	.datac(port_b4),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftLeft0~15_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~15 .lut_mask = 16'h0A0C;
defparam \ShiftLeft0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N22
cycloneive_lcell_comb \ShiftLeft0~16 (
// Equation(s):
// \ShiftLeft0~16_combout  = (\ShiftLeft0~15_combout ) # ((!\port_b~4_combout  & (\port_b~7_combout  & \rdat1[1]~1_combout )))

	.dataa(port_b2),
	.datab(port_b4),
	.datac(\ShiftLeft0~15_combout ),
	.datad(rdat1_1),
	.cin(gnd),
	.combout(\ShiftLeft0~16_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~16 .lut_mask = 16'hF4F0;
defparam \ShiftLeft0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N12
cycloneive_lcell_comb \ShiftLeft0~52 (
// Equation(s):
// \ShiftLeft0~52_combout  = (\port_b~4_combout  & ((\ShiftLeft0~37_combout ))) # (!\port_b~4_combout  & (\ShiftLeft0~25_combout ))

	.dataa(port_b2),
	.datab(\ShiftLeft0~25_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~37_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~52 .lut_mask = 16'hEE44;
defparam \ShiftLeft0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N10
cycloneive_lcell_comb \ShiftLeft0~53 (
// Equation(s):
// \ShiftLeft0~53_combout  = (\port_b~10_combout  & (\ShiftLeft0~19_combout )) # (!\port_b~10_combout  & ((\ShiftLeft0~52_combout )))

	.dataa(gnd),
	.datab(port_b6),
	.datac(\ShiftLeft0~19_combout ),
	.datad(\ShiftLeft0~52_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~53 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N16
cycloneive_lcell_comb \ShiftLeft0~54 (
// Equation(s):
// \ShiftLeft0~54_combout  = (\port_b~14_combout  & (!\port_b~10_combout  & (\ShiftLeft0~16_combout ))) # (!\port_b~14_combout  & (((\ShiftLeft0~53_combout ))))

	.dataa(port_b7),
	.datab(port_b6),
	.datac(\ShiftLeft0~16_combout ),
	.datad(\ShiftLeft0~53_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~54 .lut_mask = 16'h7520;
defparam \ShiftLeft0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N24
cycloneive_lcell_comb \ShiftLeft0~44 (
// Equation(s):
// \ShiftLeft0~44_combout  = (!\port_b~4_combout  & ((\port_b~7_combout  & (\rdat1[13]~25_combout )) # (!\port_b~7_combout  & ((\rdat1[14]~23_combout )))))

	.dataa(port_b4),
	.datab(rdat1_13),
	.datac(rdat1_14),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftLeft0~44_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~44 .lut_mask = 16'h00D8;
defparam \ShiftLeft0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N2
cycloneive_lcell_comb \ShiftLeft0~45 (
// Equation(s):
// \ShiftLeft0~45_combout  = (\ShiftLeft0~44_combout ) # ((\port_b~4_combout  & \ShiftLeft0~26_combout ))

	.dataa(port_b2),
	.datab(gnd),
	.datac(\ShiftLeft0~26_combout ),
	.datad(\ShiftLeft0~44_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~45_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~45 .lut_mask = 16'hFFA0;
defparam \ShiftLeft0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N26
cycloneive_lcell_comb \ShiftLeft0~46 (
// Equation(s):
// \ShiftLeft0~46_combout  = (\port_b~7_combout  & ((\port_b~4_combout  & (\rdat1[15]~21_combout )) # (!\port_b~4_combout  & ((\rdat1[17]~63_combout )))))

	.dataa(port_b2),
	.datab(rdat1_15),
	.datac(port_b4),
	.datad(rdat1_17),
	.cin(gnd),
	.combout(\ShiftLeft0~46_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~46 .lut_mask = 16'hD080;
defparam \ShiftLeft0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N20
cycloneive_lcell_comb \ShiftLeft0~47 (
// Equation(s):
// \ShiftLeft0~47_combout  = (!\port_b~7_combout  & ((\port_b~4_combout  & ((\rdat1[16]~19_combout ))) # (!\port_b~4_combout  & (\rdat1[18]~59_combout ))))

	.dataa(port_b2),
	.datab(rdat1_18),
	.datac(port_b4),
	.datad(rdat1_16),
	.cin(gnd),
	.combout(\ShiftLeft0~47_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~47 .lut_mask = 16'h0E04;
defparam \ShiftLeft0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N20
cycloneive_lcell_comb \ShiftLeft0~48 (
// Equation(s):
// \ShiftLeft0~48_combout  = (\port_b~10_combout  & (\ShiftLeft0~45_combout )) # (!\port_b~10_combout  & (((\ShiftLeft0~46_combout ) # (\ShiftLeft0~47_combout ))))

	.dataa(port_b6),
	.datab(\ShiftLeft0~45_combout ),
	.datac(\ShiftLeft0~46_combout ),
	.datad(\ShiftLeft0~47_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~48_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~48 .lut_mask = 16'hDDD8;
defparam \ShiftLeft0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N6
cycloneive_lcell_comb \myif.out[26]~43 (
// Equation(s):
// \myif.out[26]~43_combout  = (\myif.out[5]~16_combout  & (((\myif.out[5]~17_combout ) # (\ShiftLeft0~48_combout )))) # (!\myif.out[5]~16_combout  & (\ShiftLeft0~51_combout  & (!\myif.out[5]~17_combout )))

	.dataa(\ShiftLeft0~51_combout ),
	.datab(\myif.out[5]~16_combout ),
	.datac(\myif.out[5]~17_combout ),
	.datad(\ShiftLeft0~48_combout ),
	.cin(gnd),
	.combout(\myif.out[26]~43_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[26]~43 .lut_mask = 16'hCEC2;
defparam \myif.out[26]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N22
cycloneive_lcell_comb \myif.out[26]~44 (
// Equation(s):
// \myif.out[26]~44_combout  = (\myif.out[5]~17_combout  & ((\myif.out[26]~43_combout  & ((\ShiftLeft0~54_combout ))) # (!\myif.out[26]~43_combout  & (\ShiftLeft0~43_combout )))) # (!\myif.out[5]~17_combout  & (((\myif.out[26]~43_combout ))))

	.dataa(\ShiftLeft0~43_combout ),
	.datab(\ShiftLeft0~54_combout ),
	.datac(\myif.out[5]~17_combout ),
	.datad(\myif.out[26]~43_combout ),
	.cin(gnd),
	.combout(\myif.out[26]~44_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[26]~44 .lut_mask = 16'hCFA0;
defparam \myif.out[26]~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N14
cycloneive_lcell_comb \myif.out[26]~45 (
// Equation(s):
// \myif.out[26]~45_combout  = (idex_ifaluop_o_2 & ((\out~16_combout ) # ((!\myif.out[5]~20_combout )))) # (!idex_ifaluop_o_2 & (((\myif.out[26]~44_combout  & \myif.out[5]~20_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\out~16_combout ),
	.datac(\myif.out[26]~44_combout ),
	.datad(\myif.out[5]~20_combout ),
	.cin(gnd),
	.combout(\myif.out[26]~45_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[26]~45 .lut_mask = 16'hD8AA;
defparam \myif.out[26]~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N18
cycloneive_lcell_comb \Add0~50 (
// Equation(s):
// \Add0~50_combout  = (\port_b~40_combout  & ((\rdat1[25]~47_combout  & (\Add0~49  & VCC)) # (!\rdat1[25]~47_combout  & (!\Add0~49 )))) # (!\port_b~40_combout  & ((\rdat1[25]~47_combout  & (!\Add0~49 )) # (!\rdat1[25]~47_combout  & ((\Add0~49 ) # (GND)))))
// \Add0~51  = CARRY((\port_b~40_combout  & (!\rdat1[25]~47_combout  & !\Add0~49 )) # (!\port_b~40_combout  & ((!\Add0~49 ) # (!\rdat1[25]~47_combout ))))

	.dataa(port_b30),
	.datab(rdat1_25),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~49 ),
	.combout(\Add0~50_combout ),
	.cout(\Add0~51 ));
// synopsys translate_off
defparam \Add0~50 .lut_mask = 16'h9617;
defparam \Add0~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N20
cycloneive_lcell_comb \Add0~52 (
// Equation(s):
// \Add0~52_combout  = ((\rdat1[26]~43_combout  $ (\port_b~42_combout  $ (!\Add0~51 )))) # (GND)
// \Add0~53  = CARRY((\rdat1[26]~43_combout  & ((\port_b~42_combout ) # (!\Add0~51 ))) # (!\rdat1[26]~43_combout  & (\port_b~42_combout  & !\Add0~51 )))

	.dataa(rdat1_26),
	.datab(port_b32),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~51 ),
	.combout(\Add0~52_combout ),
	.cout(\Add0~53 ));
// synopsys translate_off
defparam \Add0~52 .lut_mask = 16'h698E;
defparam \Add0~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N8
cycloneive_lcell_comb \myif.out[26]~46 (
// Equation(s):
// \myif.out[26]~46_combout  = (idex_ifaluop_o_1 & ((\myif.out[26]~45_combout  & (\out~15_combout )) # (!\myif.out[26]~45_combout  & ((\Add0~52_combout ))))) # (!idex_ifaluop_o_1 & (((\myif.out[26]~45_combout ))))

	.dataa(\out~15_combout ),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[26]~45_combout ),
	.datad(\Add0~52_combout ),
	.cin(gnd),
	.combout(\myif.out[26]~46_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[26]~46 .lut_mask = 16'hBCB0;
defparam \myif.out[26]~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N8
cycloneive_lcell_comb \out~17 (
// Equation(s):
// \out~17_combout  = (\port_b~39_combout ) # ((\rdat1[25]~47_combout ) # ((\port_b~0_combout  & fuifrtReplace_25)))

	.dataa(port_b29),
	.datab(port_b),
	.datac(rdat1_25),
	.datad(fuifrtReplace_25),
	.cin(gnd),
	.combout(\out~17_combout ),
	.cout());
// synopsys translate_off
defparam \out~17 .lut_mask = 16'hFEFA;
defparam \out~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N0
cycloneive_lcell_comb \ShiftRight0~17 (
// Equation(s):
// \ShiftRight0~17_combout  = (!\port_b~7_combout  & ((\port_b~4_combout  & (\rdat1[31]~35_combout )) # (!\port_b~4_combout  & ((\rdat1[29]~37_combout )))))

	.dataa(port_b4),
	.datab(rdat1_311),
	.datac(port_b2),
	.datad(rdat1_29),
	.cin(gnd),
	.combout(\ShiftRight0~17_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~17 .lut_mask = 16'h4540;
defparam \ShiftRight0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N22
cycloneive_lcell_comb \ShiftRight0~18 (
// Equation(s):
// \ShiftRight0~18_combout  = (\ShiftRight0~17_combout ) # ((\port_b~7_combout  & (!\port_b~4_combout  & \rdat1[30]~39_combout )))

	.dataa(port_b4),
	.datab(port_b2),
	.datac(rdat1_30),
	.datad(\ShiftRight0~17_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~18_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~18 .lut_mask = 16'hFF20;
defparam \ShiftRight0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N16
cycloneive_lcell_comb \ShiftRight0~72 (
// Equation(s):
// \ShiftRight0~72_combout  = (!\port_b~14_combout  & ((\port_b~10_combout  & ((\ShiftRight0~18_combout ))) # (!\port_b~10_combout  & (\ShiftRight0~21_combout ))))

	.dataa(\ShiftRight0~21_combout ),
	.datab(port_b7),
	.datac(\ShiftRight0~18_combout ),
	.datad(port_b6),
	.cin(gnd),
	.combout(\ShiftRight0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~72 .lut_mask = 16'h3022;
defparam \ShiftRight0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N30
cycloneive_lcell_comb \myif.out[25]~48 (
// Equation(s):
// \myif.out[25]~48_combout  = (idex_ifaluop_o_2 & ((\out~17_combout ) # ((!\myif.out[13]~23_combout )))) # (!idex_ifaluop_o_2 & (((\ShiftRight0~72_combout  & \myif.out[13]~23_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\out~17_combout ),
	.datac(\ShiftRight0~72_combout ),
	.datad(\myif.out[13]~23_combout ),
	.cin(gnd),
	.combout(\myif.out[25]~48_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[25]~48 .lut_mask = 16'hD8AA;
defparam \myif.out[25]~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N8
cycloneive_lcell_comb \myif.out[25]~49 (
// Equation(s):
// \myif.out[25]~49_combout  = (idex_ifaluop_o_1 & ((\myif.out[25]~48_combout  & (!\out~17_combout )) # (!\myif.out[25]~48_combout  & ((\Add1~50_combout ))))) # (!idex_ifaluop_o_1 & (((\myif.out[25]~48_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(\out~17_combout ),
	.datac(\myif.out[25]~48_combout ),
	.datad(\Add1~50_combout ),
	.cin(gnd),
	.combout(\myif.out[25]~49_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[25]~49 .lut_mask = 16'h7A70;
defparam \myif.out[25]~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N12
cycloneive_lcell_comb \out~18 (
// Equation(s):
// \out~18_combout  = \rdat1[25]~47_combout  $ (((\port_b~39_combout ) # ((\port_b~0_combout  & fuifrtReplace_25))))

	.dataa(port_b29),
	.datab(port_b),
	.datac(rdat1_25),
	.datad(fuifrtReplace_25),
	.cin(gnd),
	.combout(\out~18_combout ),
	.cout());
// synopsys translate_off
defparam \out~18 .lut_mask = 16'h1E5A;
defparam \out~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N20
cycloneive_lcell_comb \out~19 (
// Equation(s):
// \out~19_combout  = (\rdat1[25]~47_combout  & ((\port_b~39_combout ) # ((\port_b~0_combout  & fuifrtReplace_25))))

	.dataa(port_b),
	.datab(rdat1_25),
	.datac(port_b29),
	.datad(fuifrtReplace_25),
	.cin(gnd),
	.combout(\out~19_combout ),
	.cout());
// synopsys translate_off
defparam \out~19 .lut_mask = 16'hC8C0;
defparam \out~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N22
cycloneive_lcell_comb \ShiftLeft0~64 (
// Equation(s):
// \ShiftLeft0~64_combout  = (\port_b~7_combout  & (((\port_b~4_combout )))) # (!\port_b~7_combout  & ((\port_b~4_combout  & ((\rdat1[23]~53_combout ))) # (!\port_b~4_combout  & (\rdat1[25]~47_combout ))))

	.dataa(rdat1_25),
	.datab(port_b4),
	.datac(rdat1_23),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftLeft0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~64 .lut_mask = 16'hFC22;
defparam \ShiftLeft0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N24
cycloneive_lcell_comb \ShiftLeft0~65 (
// Equation(s):
// \ShiftLeft0~65_combout  = (\port_b~7_combout  & ((\ShiftLeft0~64_combout  & ((\rdat1[22]~51_combout ))) # (!\ShiftLeft0~64_combout  & (\rdat1[24]~49_combout )))) # (!\port_b~7_combout  & (((\ShiftLeft0~64_combout ))))

	.dataa(rdat1_24),
	.datab(port_b4),
	.datac(\ShiftLeft0~64_combout ),
	.datad(rdat1_22),
	.cin(gnd),
	.combout(\ShiftLeft0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~65 .lut_mask = 16'hF838;
defparam \ShiftLeft0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N18
cycloneive_lcell_comb \myif.out[25]~50 (
// Equation(s):
// \myif.out[25]~50_combout  = (\myif.out[5]~17_combout  & ((\ShiftLeft0~63_combout ) # ((\myif.out[5]~16_combout )))) # (!\myif.out[5]~17_combout  & (((\ShiftLeft0~65_combout  & !\myif.out[5]~16_combout ))))

	.dataa(\ShiftLeft0~63_combout ),
	.datab(\myif.out[5]~17_combout ),
	.datac(\ShiftLeft0~65_combout ),
	.datad(\myif.out[5]~16_combout ),
	.cin(gnd),
	.combout(\myif.out[25]~50_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[25]~50 .lut_mask = 16'hCCB8;
defparam \myif.out[25]~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N4
cycloneive_lcell_comb \ShiftLeft0~55 (
// Equation(s):
// \ShiftLeft0~55_combout  = (\port_b~7_combout  & (\rdat1[10]~31_combout )) # (!\port_b~7_combout  & ((\rdat1[11]~29_combout )))

	.dataa(gnd),
	.datab(rdat1_10),
	.datac(port_b4),
	.datad(rdat1_11),
	.cin(gnd),
	.combout(\ShiftLeft0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~55 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N26
cycloneive_lcell_comb \ShiftLeft0~56 (
// Equation(s):
// \ShiftLeft0~56_combout  = (\port_b~7_combout  & (\rdat1[12]~27_combout )) # (!\port_b~7_combout  & ((\rdat1[13]~25_combout )))

	.dataa(port_b4),
	.datab(gnd),
	.datac(rdat1_12),
	.datad(rdat1_13),
	.cin(gnd),
	.combout(\ShiftLeft0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~56 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N8
cycloneive_lcell_comb \ShiftLeft0~57 (
// Equation(s):
// \ShiftLeft0~57_combout  = (\port_b~4_combout  & (\ShiftLeft0~55_combout )) # (!\port_b~4_combout  & ((\ShiftLeft0~56_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~55_combout ),
	.datac(\ShiftLeft0~56_combout ),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftLeft0~57_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~57 .lut_mask = 16'hCCF0;
defparam \ShiftLeft0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N22
cycloneive_lcell_comb \ShiftLeft0~58 (
// Equation(s):
// \ShiftLeft0~58_combout  = (!\port_b~4_combout  & ((\port_b~7_combout  & ((\rdat1[16]~19_combout ))) # (!\port_b~7_combout  & (\rdat1[17]~63_combout ))))

	.dataa(port_b2),
	.datab(rdat1_17),
	.datac(port_b4),
	.datad(rdat1_16),
	.cin(gnd),
	.combout(\ShiftLeft0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~58 .lut_mask = 16'h5404;
defparam \ShiftLeft0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N0
cycloneive_lcell_comb \ShiftLeft0~59 (
// Equation(s):
// \ShiftLeft0~59_combout  = (\port_b~7_combout  & ((\rdat1[14]~23_combout ))) # (!\port_b~7_combout  & (\rdat1[15]~21_combout ))

	.dataa(gnd),
	.datab(port_b4),
	.datac(rdat1_15),
	.datad(rdat1_14),
	.cin(gnd),
	.combout(\ShiftLeft0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~59 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N10
cycloneive_lcell_comb \ShiftLeft0~60 (
// Equation(s):
// \ShiftLeft0~60_combout  = (\ShiftLeft0~58_combout ) # ((\port_b~4_combout  & \ShiftLeft0~59_combout ))

	.dataa(port_b2),
	.datab(gnd),
	.datac(\ShiftLeft0~58_combout ),
	.datad(\ShiftLeft0~59_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~60 .lut_mask = 16'hFAF0;
defparam \ShiftLeft0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N8
cycloneive_lcell_comb \ShiftLeft0~61 (
// Equation(s):
// \ShiftLeft0~61_combout  = (\port_b~10_combout  & (\ShiftLeft0~57_combout )) # (!\port_b~10_combout  & ((\ShiftLeft0~60_combout )))

	.dataa(port_b6),
	.datab(gnd),
	.datac(\ShiftLeft0~57_combout ),
	.datad(\ShiftLeft0~60_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~61 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N4
cycloneive_lcell_comb \ShiftLeft0~67 (
// Equation(s):
// \ShiftLeft0~67_combout  = (\port_b~7_combout  & (\rdat1[4]~7_combout )) # (!\port_b~7_combout  & ((\rdat1[5]~17_combout )))

	.dataa(port_b4),
	.datab(gnd),
	.datac(rdat1_41),
	.datad(rdat1_5),
	.cin(gnd),
	.combout(\ShiftLeft0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~67 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N2
cycloneive_lcell_comb \ShiftLeft0~68 (
// Equation(s):
// \ShiftLeft0~68_combout  = (\port_b~4_combout  & (\ShiftLeft0~66_combout )) # (!\port_b~4_combout  & ((\ShiftLeft0~67_combout )))

	.dataa(\ShiftLeft0~66_combout ),
	.datab(port_b2),
	.datac(\ShiftLeft0~67_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~68 .lut_mask = 16'hB8B8;
defparam \ShiftLeft0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N6
cycloneive_lcell_comb \ShiftLeft0~70 (
// Equation(s):
// \ShiftLeft0~70_combout  = (\port_b~7_combout  & ((\rdat1[8]~11_combout ))) # (!\port_b~7_combout  & (\rdat1[9]~33_combout ))

	.dataa(port_b4),
	.datab(gnd),
	.datac(rdat1_9),
	.datad(rdat1_8),
	.cin(gnd),
	.combout(\ShiftLeft0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~70 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N16
cycloneive_lcell_comb \ShiftLeft0~71 (
// Equation(s):
// \ShiftLeft0~71_combout  = (\port_b~4_combout  & (\ShiftLeft0~69_combout )) # (!\port_b~4_combout  & ((\ShiftLeft0~70_combout )))

	.dataa(\ShiftLeft0~69_combout ),
	.datab(gnd),
	.datac(port_b2),
	.datad(\ShiftLeft0~70_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~71 .lut_mask = 16'hAFA0;
defparam \ShiftLeft0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N30
cycloneive_lcell_comb \ShiftLeft0~72 (
// Equation(s):
// \ShiftLeft0~72_combout  = (\port_b~10_combout  & (\ShiftLeft0~68_combout )) # (!\port_b~10_combout  & ((\ShiftLeft0~71_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~68_combout ),
	.datac(port_b6),
	.datad(\ShiftLeft0~71_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~72 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N28
cycloneive_lcell_comb \ShiftLeft0~73 (
// Equation(s):
// \ShiftLeft0~73_combout  = (\port_b~14_combout  & (\ShiftLeft0~12_combout  & ((!\ShiftLeft0~13_combout )))) # (!\port_b~14_combout  & (((\ShiftLeft0~72_combout ))))

	.dataa(\ShiftLeft0~12_combout ),
	.datab(port_b7),
	.datac(\ShiftLeft0~72_combout ),
	.datad(\ShiftLeft0~13_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~73 .lut_mask = 16'h30B8;
defparam \ShiftLeft0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N30
cycloneive_lcell_comb \myif.out[25]~51 (
// Equation(s):
// \myif.out[25]~51_combout  = (\myif.out[5]~16_combout  & ((\myif.out[25]~50_combout  & ((\ShiftLeft0~73_combout ))) # (!\myif.out[25]~50_combout  & (\ShiftLeft0~61_combout )))) # (!\myif.out[5]~16_combout  & (\myif.out[25]~50_combout ))

	.dataa(\myif.out[5]~16_combout ),
	.datab(\myif.out[25]~50_combout ),
	.datac(\ShiftLeft0~61_combout ),
	.datad(\ShiftLeft0~73_combout ),
	.cin(gnd),
	.combout(\myif.out[25]~51_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[25]~51 .lut_mask = 16'hEC64;
defparam \myif.out[25]~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N6
cycloneive_lcell_comb \myif.out[25]~52 (
// Equation(s):
// \myif.out[25]~52_combout  = (\myif.out[5]~20_combout  & ((idex_ifaluop_o_2 & (\out~19_combout )) # (!idex_ifaluop_o_2 & ((\myif.out[25]~51_combout ))))) # (!\myif.out[5]~20_combout  & (idex_ifaluop_o_2))

	.dataa(\myif.out[5]~20_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\out~19_combout ),
	.datad(\myif.out[25]~51_combout ),
	.cin(gnd),
	.combout(\myif.out[25]~52_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[25]~52 .lut_mask = 16'hE6C4;
defparam \myif.out[25]~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N16
cycloneive_lcell_comb \myif.out[25]~53 (
// Equation(s):
// \myif.out[25]~53_combout  = (idex_ifaluop_o_1 & ((\myif.out[25]~52_combout  & ((\out~18_combout ))) # (!\myif.out[25]~52_combout  & (\Add0~50_combout )))) # (!idex_ifaluop_o_1 & (((\myif.out[25]~52_combout ))))

	.dataa(\Add0~50_combout ),
	.datab(\out~18_combout ),
	.datac(idex_ifaluop_o_1),
	.datad(\myif.out[25]~52_combout ),
	.cin(gnd),
	.combout(\myif.out[25]~53_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[25]~53 .lut_mask = 16'hCFA0;
defparam \myif.out[25]~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N4
cycloneive_lcell_comb \out~21 (
// Equation(s):
// \out~21_combout  = \rdat1[27]~45_combout  $ (((\port_b~51_combout ) # ((fuifrtReplace_27 & \port_b~0_combout ))))

	.dataa(rdat1_27),
	.datab(fuifrtReplace_27),
	.datac(port_b),
	.datad(port_b41),
	.cin(gnd),
	.combout(\out~21_combout ),
	.cout());
// synopsys translate_off
defparam \out~21 .lut_mask = 16'h556A;
defparam \out~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N26
cycloneive_lcell_comb \out~22 (
// Equation(s):
// \out~22_combout  = (\rdat1[27]~45_combout  & ((\port_b~51_combout ) # ((\port_b~0_combout  & fuifrtReplace_27))))

	.dataa(rdat1_27),
	.datab(port_b41),
	.datac(port_b),
	.datad(fuifrtReplace_27),
	.cin(gnd),
	.combout(\out~22_combout ),
	.cout());
// synopsys translate_off
defparam \out~22 .lut_mask = 16'hA888;
defparam \out~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N24
cycloneive_lcell_comb \ShiftLeft0~12 (
// Equation(s):
// \ShiftLeft0~12_combout  = (\port_b~7_combout  & (\rdat1[0]~3_combout )) # (!\port_b~7_combout  & ((\rdat1[1]~1_combout )))

	.dataa(port_b4),
	.datab(rdat1_0),
	.datac(gnd),
	.datad(rdat1_1),
	.cin(gnd),
	.combout(\ShiftLeft0~12_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~12 .lut_mask = 16'hDD88;
defparam \ShiftLeft0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N20
cycloneive_lcell_comb \ShiftLeft0~66 (
// Equation(s):
// \ShiftLeft0~66_combout  = (\port_b~7_combout  & ((\rdat1[2]~5_combout ))) # (!\port_b~7_combout  & (\rdat1[3]~9_combout ))

	.dataa(gnd),
	.datab(rdat1_31),
	.datac(rdat1_2),
	.datad(port_b4),
	.cin(gnd),
	.combout(\ShiftLeft0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~66 .lut_mask = 16'hF0CC;
defparam \ShiftLeft0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N14
cycloneive_lcell_comb \ShiftLeft0~85 (
// Equation(s):
// \ShiftLeft0~85_combout  = (\port_b~4_combout  & (\ShiftLeft0~12_combout )) # (!\port_b~4_combout  & ((\ShiftLeft0~66_combout )))

	.dataa(port_b2),
	.datab(gnd),
	.datac(\ShiftLeft0~12_combout ),
	.datad(\ShiftLeft0~66_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~85_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~85 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N4
cycloneive_lcell_comb \ShiftLeft0~69 (
// Equation(s):
// \ShiftLeft0~69_combout  = (\port_b~7_combout  & ((\rdat1[6]~15_combout ))) # (!\port_b~7_combout  & (\rdat1[7]~13_combout ))

	.dataa(rdat1_7),
	.datab(gnd),
	.datac(rdat1_6),
	.datad(port_b4),
	.cin(gnd),
	.combout(\ShiftLeft0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~69 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N20
cycloneive_lcell_comb \ShiftLeft0~82 (
// Equation(s):
// \ShiftLeft0~82_combout  = (\port_b~4_combout  & (\ShiftLeft0~67_combout )) # (!\port_b~4_combout  & ((\ShiftLeft0~69_combout )))

	.dataa(gnd),
	.datab(port_b2),
	.datac(\ShiftLeft0~67_combout ),
	.datad(\ShiftLeft0~69_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~82 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N0
cycloneive_lcell_comb \ShiftLeft0~83 (
// Equation(s):
// \ShiftLeft0~83_combout  = (\port_b~4_combout  & ((\ShiftLeft0~70_combout ))) # (!\port_b~4_combout  & (\ShiftLeft0~55_combout ))

	.dataa(port_b2),
	.datab(gnd),
	.datac(\ShiftLeft0~55_combout ),
	.datad(\ShiftLeft0~70_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~83 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N10
cycloneive_lcell_comb \ShiftLeft0~84 (
// Equation(s):
// \ShiftLeft0~84_combout  = (\port_b~10_combout  & (\ShiftLeft0~82_combout )) # (!\port_b~10_combout  & ((\ShiftLeft0~83_combout )))

	.dataa(port_b6),
	.datab(gnd),
	.datac(\ShiftLeft0~82_combout ),
	.datad(\ShiftLeft0~83_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~84 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N24
cycloneive_lcell_comb \ShiftLeft0~86 (
// Equation(s):
// \ShiftLeft0~86_combout  = (\port_b~14_combout  & (!\port_b~10_combout  & (\ShiftLeft0~85_combout ))) # (!\port_b~14_combout  & (((\ShiftLeft0~84_combout ))))

	.dataa(port_b6),
	.datab(port_b7),
	.datac(\ShiftLeft0~85_combout ),
	.datad(\ShiftLeft0~84_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~86 .lut_mask = 16'h7340;
defparam \ShiftLeft0~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N20
cycloneive_lcell_comb \ShiftLeft0~75 (
// Equation(s):
// \ShiftLeft0~75_combout  = (\port_b~4_combout  & (\ShiftLeft0~56_combout )) # (!\port_b~4_combout  & ((\ShiftLeft0~59_combout )))

	.dataa(port_b2),
	.datab(gnd),
	.datac(\ShiftLeft0~56_combout ),
	.datad(\ShiftLeft0~59_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~75 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N14
cycloneive_lcell_comb \ShiftLeft0~76 (
// Equation(s):
// \ShiftLeft0~76_combout  = (\port_b~7_combout  & ((\port_b~4_combout  & ((\rdat1[16]~19_combout ))) # (!\port_b~4_combout  & (\rdat1[18]~59_combout ))))

	.dataa(rdat1_18),
	.datab(port_b4),
	.datac(port_b2),
	.datad(rdat1_16),
	.cin(gnd),
	.combout(\ShiftLeft0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~76 .lut_mask = 16'hC808;
defparam \ShiftLeft0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N16
cycloneive_lcell_comb \ShiftLeft0~32 (
// Equation(s):
// \ShiftLeft0~32_combout  = (\port_b~4_combout  & (\rdat1[17]~63_combout )) # (!\port_b~4_combout  & ((\rdat1[19]~61_combout )))

	.dataa(gnd),
	.datab(port_b2),
	.datac(rdat1_17),
	.datad(rdat1_19),
	.cin(gnd),
	.combout(\ShiftLeft0~32_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~32 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N20
cycloneive_lcell_comb \ShiftLeft0~77 (
// Equation(s):
// \ShiftLeft0~77_combout  = (\ShiftLeft0~76_combout ) # ((!\port_b~7_combout  & \ShiftLeft0~32_combout ))

	.dataa(gnd),
	.datab(port_b4),
	.datac(\ShiftLeft0~76_combout ),
	.datad(\ShiftLeft0~32_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~77 .lut_mask = 16'hF3F0;
defparam \ShiftLeft0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N28
cycloneive_lcell_comb \ShiftLeft0~78 (
// Equation(s):
// \ShiftLeft0~78_combout  = (\port_b~10_combout  & (\ShiftLeft0~75_combout )) # (!\port_b~10_combout  & ((\ShiftLeft0~77_combout )))

	.dataa(gnd),
	.datab(port_b6),
	.datac(\ShiftLeft0~75_combout ),
	.datad(\ShiftLeft0~77_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~78 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N20
cycloneive_lcell_comb \myif.out[27]~57 (
// Equation(s):
// \myif.out[27]~57_combout  = (\myif.out[5]~17_combout  & (((\myif.out[5]~16_combout )))) # (!\myif.out[5]~17_combout  & ((\myif.out[5]~16_combout  & ((\ShiftLeft0~78_combout ))) # (!\myif.out[5]~16_combout  & (\ShiftLeft0~81_combout ))))

	.dataa(\ShiftLeft0~81_combout ),
	.datab(\myif.out[5]~17_combout ),
	.datac(\myif.out[5]~16_combout ),
	.datad(\ShiftLeft0~78_combout ),
	.cin(gnd),
	.combout(\myif.out[27]~57_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[27]~57 .lut_mask = 16'hF2C2;
defparam \myif.out[27]~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N6
cycloneive_lcell_comb \myif.out[27]~58 (
// Equation(s):
// \myif.out[27]~58_combout  = (\myif.out[5]~17_combout  & ((\myif.out[27]~57_combout  & ((\ShiftLeft0~86_combout ))) # (!\myif.out[27]~57_combout  & (\ShiftLeft0~74_combout )))) # (!\myif.out[5]~17_combout  & (((\myif.out[27]~57_combout ))))

	.dataa(\ShiftLeft0~74_combout ),
	.datab(\myif.out[5]~17_combout ),
	.datac(\ShiftLeft0~86_combout ),
	.datad(\myif.out[27]~57_combout ),
	.cin(gnd),
	.combout(\myif.out[27]~58_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[27]~58 .lut_mask = 16'hF388;
defparam \myif.out[27]~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N16
cycloneive_lcell_comb \myif.out[27]~59 (
// Equation(s):
// \myif.out[27]~59_combout  = (idex_ifaluop_o_2 & ((\out~22_combout ) # ((!\myif.out[5]~20_combout )))) # (!idex_ifaluop_o_2 & (((\myif.out[5]~20_combout  & \myif.out[27]~58_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\out~22_combout ),
	.datac(\myif.out[5]~20_combout ),
	.datad(\myif.out[27]~58_combout ),
	.cin(gnd),
	.combout(\myif.out[27]~59_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[27]~59 .lut_mask = 16'hDA8A;
defparam \myif.out[27]~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N22
cycloneive_lcell_comb \Add0~54 (
// Equation(s):
// \Add0~54_combout  = (\rdat1[27]~45_combout  & ((\port_b~52_combout  & (\Add0~53  & VCC)) # (!\port_b~52_combout  & (!\Add0~53 )))) # (!\rdat1[27]~45_combout  & ((\port_b~52_combout  & (!\Add0~53 )) # (!\port_b~52_combout  & ((\Add0~53 ) # (GND)))))
// \Add0~55  = CARRY((\rdat1[27]~45_combout  & (!\port_b~52_combout  & !\Add0~53 )) # (!\rdat1[27]~45_combout  & ((!\Add0~53 ) # (!\port_b~52_combout ))))

	.dataa(rdat1_27),
	.datab(port_b42),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~53 ),
	.combout(\Add0~54_combout ),
	.cout(\Add0~55 ));
// synopsys translate_off
defparam \Add0~54 .lut_mask = 16'h9617;
defparam \Add0~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N30
cycloneive_lcell_comb \myif.out[27]~60 (
// Equation(s):
// \myif.out[27]~60_combout  = (idex_ifaluop_o_1 & ((\myif.out[27]~59_combout  & (\out~21_combout )) # (!\myif.out[27]~59_combout  & ((\Add0~54_combout ))))) # (!idex_ifaluop_o_1 & (((\myif.out[27]~59_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(\out~21_combout ),
	.datac(\myif.out[27]~59_combout ),
	.datad(\Add0~54_combout ),
	.cin(gnd),
	.combout(\myif.out[27]~60_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[27]~60 .lut_mask = 16'hDAD0;
defparam \myif.out[27]~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N18
cycloneive_lcell_comb \out~20 (
// Equation(s):
// \out~20_combout  = (\port_b~51_combout ) # ((\rdat1[27]~45_combout ) # ((\port_b~0_combout  & fuifrtReplace_27)))

	.dataa(port_b41),
	.datab(port_b),
	.datac(rdat1_27),
	.datad(fuifrtReplace_27),
	.cin(gnd),
	.combout(\out~20_combout ),
	.cout());
// synopsys translate_off
defparam \out~20 .lut_mask = 16'hFEFA;
defparam \out~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N22
cycloneive_lcell_comb \Add1~54 (
// Equation(s):
// \Add1~54_combout  = (\rdat1[27]~45_combout  & ((\port_b~52_combout  & (!\Add1~53 )) # (!\port_b~52_combout  & (\Add1~53  & VCC)))) # (!\rdat1[27]~45_combout  & ((\port_b~52_combout  & ((\Add1~53 ) # (GND))) # (!\port_b~52_combout  & (!\Add1~53 ))))
// \Add1~55  = CARRY((\rdat1[27]~45_combout  & (\port_b~52_combout  & !\Add1~53 )) # (!\rdat1[27]~45_combout  & ((\port_b~52_combout ) # (!\Add1~53 ))))

	.dataa(rdat1_27),
	.datab(port_b42),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~53 ),
	.combout(\Add1~54_combout ),
	.cout(\Add1~55 ));
// synopsys translate_off
defparam \Add1~54 .lut_mask = 16'h694D;
defparam \Add1~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N26
cycloneive_lcell_comb \ShiftRight0~74 (
// Equation(s):
// \ShiftRight0~74_combout  = (\port_b~7_combout  & ((\port_b~4_combout  & (\rdat1[30]~39_combout )) # (!\port_b~4_combout  & ((\rdat1[28]~41_combout )))))

	.dataa(rdat1_30),
	.datab(rdat1_28),
	.datac(port_b4),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftRight0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~74 .lut_mask = 16'hA0C0;
defparam \ShiftRight0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N20
cycloneive_lcell_comb \ShiftRight0~75 (
// Equation(s):
// \ShiftRight0~75_combout  = (\ShiftRight0~74_combout ) # ((!\port_b~7_combout  & \ShiftRight0~46_combout ))

	.dataa(gnd),
	.datab(port_b4),
	.datac(\ShiftRight0~74_combout ),
	.datad(\ShiftRight0~46_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~75 .lut_mask = 16'hF3F0;
defparam \ShiftRight0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N10
cycloneive_lcell_comb \ShiftRight0~76 (
// Equation(s):
// \ShiftRight0~76_combout  = (!\port_b~14_combout  & ((\port_b~10_combout  & (\ShiftRight0~73_combout )) # (!\port_b~10_combout  & ((\ShiftRight0~75_combout )))))

	.dataa(\ShiftRight0~73_combout ),
	.datab(port_b6),
	.datac(port_b7),
	.datad(\ShiftRight0~75_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~76 .lut_mask = 16'h0B08;
defparam \ShiftRight0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N12
cycloneive_lcell_comb \myif.out[27]~55 (
// Equation(s):
// \myif.out[27]~55_combout  = (idex_ifaluop_o_2 & ((\out~20_combout ) # ((!\myif.out[13]~23_combout )))) # (!idex_ifaluop_o_2 & (((\ShiftRight0~76_combout  & \myif.out[13]~23_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\out~20_combout ),
	.datac(\ShiftRight0~76_combout ),
	.datad(\myif.out[13]~23_combout ),
	.cin(gnd),
	.combout(\myif.out[27]~55_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[27]~55 .lut_mask = 16'hD8AA;
defparam \myif.out[27]~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N6
cycloneive_lcell_comb \myif.out[27]~56 (
// Equation(s):
// \myif.out[27]~56_combout  = (idex_ifaluop_o_1 & ((\myif.out[27]~55_combout  & (!\out~20_combout )) # (!\myif.out[27]~55_combout  & ((\Add1~54_combout ))))) # (!idex_ifaluop_o_1 & (((\myif.out[27]~55_combout ))))

	.dataa(\out~20_combout ),
	.datab(\Add1~54_combout ),
	.datac(idex_ifaluop_o_1),
	.datad(\myif.out[27]~55_combout ),
	.cin(gnd),
	.combout(\myif.out[27]~56_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[27]~56 .lut_mask = 16'h5FC0;
defparam \myif.out[27]~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N10
cycloneive_lcell_comb \out~24 (
// Equation(s):
// \out~24_combout  = \rdat1[5]~17_combout  $ (((\port_b~43_combout ) # ((fuifrtReplace_5 & \port_b~0_combout ))))

	.dataa(port_b33),
	.datab(fuifrtReplace_5),
	.datac(port_b),
	.datad(rdat1_5),
	.cin(gnd),
	.combout(\out~24_combout ),
	.cout());
// synopsys translate_off
defparam \out~24 .lut_mask = 16'h15EA;
defparam \out~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N8
cycloneive_lcell_comb \ShiftLeft0~87 (
// Equation(s):
// \ShiftLeft0~87_combout  = (\port_b~10_combout  & (\ShiftLeft0~12_combout  & (!\port_b~4_combout ))) # (!\port_b~10_combout  & (((\ShiftLeft0~68_combout ))))

	.dataa(\ShiftLeft0~12_combout ),
	.datab(port_b6),
	.datac(port_b2),
	.datad(\ShiftLeft0~68_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~87_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~87 .lut_mask = 16'h3B08;
defparam \ShiftLeft0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N14
cycloneive_lcell_comb \ShiftLeft0~88 (
// Equation(s):
// \ShiftLeft0~88_combout  = (!\port_b~14_combout  & \ShiftLeft0~87_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(port_b7),
	.datad(\ShiftLeft0~87_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~88_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~88 .lut_mask = 16'h0F00;
defparam \ShiftLeft0~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N14
cycloneive_lcell_comb \out~25 (
// Equation(s):
// \out~25_combout  = (\rdat1[5]~17_combout  & ((\port_b~43_combout ) # ((\port_b~0_combout  & fuifrtReplace_5))))

	.dataa(rdat1_5),
	.datab(port_b33),
	.datac(port_b),
	.datad(fuifrtReplace_5),
	.cin(gnd),
	.combout(\out~25_combout ),
	.cout());
// synopsys translate_off
defparam \out~25 .lut_mask = 16'hA888;
defparam \out~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N24
cycloneive_lcell_comb \myif.out[5]~66 (
// Equation(s):
// \myif.out[5]~66_combout  = (idex_ifaluop_o_2 & (((\out~25_combout ) # (!\myif.out[13]~23_combout )))) # (!idex_ifaluop_o_2 & (\ShiftLeft0~88_combout  & ((\myif.out[13]~23_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\ShiftLeft0~88_combout ),
	.datac(\out~25_combout ),
	.datad(\myif.out[13]~23_combout ),
	.cin(gnd),
	.combout(\myif.out[5]~66_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[5]~66 .lut_mask = 16'hE4AA;
defparam \myif.out[5]~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N4
cycloneive_lcell_comb \myif.out[5]~67 (
// Equation(s):
// \myif.out[5]~67_combout  = (idex_ifaluop_o_1 & ((\myif.out[5]~66_combout  & (\out~24_combout )) # (!\myif.out[5]~66_combout  & ((\Add0~10_combout ))))) # (!idex_ifaluop_o_1 & (((\myif.out[5]~66_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(\out~24_combout ),
	.datac(\myif.out[5]~66_combout ),
	.datad(\Add0~10_combout ),
	.cin(gnd),
	.combout(\myif.out[5]~67_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[5]~67 .lut_mask = 16'hDAD0;
defparam \myif.out[5]~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N30
cycloneive_lcell_comb \out~23 (
// Equation(s):
// \out~23_combout  = (\rdat1[5]~17_combout ) # ((\port_b~43_combout ) # ((\port_b~0_combout  & fuifrtReplace_5)))

	.dataa(rdat1_5),
	.datab(port_b33),
	.datac(port_b),
	.datad(fuifrtReplace_5),
	.cin(gnd),
	.combout(\out~23_combout ),
	.cout());
// synopsys translate_off
defparam \out~23 .lut_mask = 16'hFEEE;
defparam \out~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N4
cycloneive_lcell_comb \myif.out[5]~62 (
// Equation(s):
// \myif.out[5]~62_combout  = (\myif.out[5]~17_combout  & ((\myif.out[5]~16_combout ) # ((\ShiftRight0~14_combout )))) # (!\myif.out[5]~17_combout  & (!\myif.out[5]~16_combout  & (\ShiftRight0~7_combout )))

	.dataa(\myif.out[5]~17_combout ),
	.datab(\myif.out[5]~16_combout ),
	.datac(\ShiftRight0~7_combout ),
	.datad(\ShiftRight0~14_combout ),
	.cin(gnd),
	.combout(\myif.out[5]~62_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[5]~62 .lut_mask = 16'hBA98;
defparam \myif.out[5]~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N22
cycloneive_lcell_comb \ShiftRight0~77 (
// Equation(s):
// \ShiftRight0~77_combout  = (\port_b~10_combout  & (\ShiftRight0~28_combout )) # (!\port_b~10_combout  & ((\ShiftRight0~11_combout )))

	.dataa(port_b6),
	.datab(gnd),
	.datac(\ShiftRight0~28_combout ),
	.datad(\ShiftRight0~11_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~77 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N20
cycloneive_lcell_comb \ShiftRight0~78 (
// Equation(s):
// \ShiftRight0~78_combout  = (\port_b~10_combout  & (\ShiftRight0~21_combout )) # (!\port_b~10_combout  & ((\ShiftRight0~25_combout )))

	.dataa(gnd),
	.datab(port_b6),
	.datac(\ShiftRight0~21_combout ),
	.datad(\ShiftRight0~25_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~78 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N6
cycloneive_lcell_comb \ShiftRight0~79 (
// Equation(s):
// \ShiftRight0~79_combout  = (\port_b~14_combout  & (!\port_b~10_combout  & (\ShiftRight0~18_combout ))) # (!\port_b~14_combout  & (((\ShiftRight0~78_combout ))))

	.dataa(port_b6),
	.datab(port_b7),
	.datac(\ShiftRight0~18_combout ),
	.datad(\ShiftRight0~78_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~79 .lut_mask = 16'h7340;
defparam \ShiftRight0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N0
cycloneive_lcell_comb \myif.out[5]~63 (
// Equation(s):
// \myif.out[5]~63_combout  = (\myif.out[5]~16_combout  & ((\myif.out[5]~62_combout  & ((\ShiftRight0~79_combout ))) # (!\myif.out[5]~62_combout  & (\ShiftRight0~77_combout )))) # (!\myif.out[5]~16_combout  & (\myif.out[5]~62_combout ))

	.dataa(\myif.out[5]~16_combout ),
	.datab(\myif.out[5]~62_combout ),
	.datac(\ShiftRight0~77_combout ),
	.datad(\ShiftRight0~79_combout ),
	.cin(gnd),
	.combout(\myif.out[5]~63_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[5]~63 .lut_mask = 16'hEC64;
defparam \myif.out[5]~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N20
cycloneive_lcell_comb \myif.out[5]~64 (
// Equation(s):
// \myif.out[5]~64_combout  = (\myif.out[5]~20_combout  & ((idex_ifaluop_o_2 & (\out~23_combout )) # (!idex_ifaluop_o_2 & ((\myif.out[5]~63_combout ))))) # (!\myif.out[5]~20_combout  & (idex_ifaluop_o_2))

	.dataa(\myif.out[5]~20_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\out~23_combout ),
	.datad(\myif.out[5]~63_combout ),
	.cin(gnd),
	.combout(\myif.out[5]~64_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[5]~64 .lut_mask = 16'hE6C4;
defparam \myif.out[5]~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N26
cycloneive_lcell_comb \myif.out[5]~65 (
// Equation(s):
// \myif.out[5]~65_combout  = (idex_ifaluop_o_1 & ((\myif.out[5]~64_combout  & ((!\out~23_combout ))) # (!\myif.out[5]~64_combout  & (\Add1~10_combout )))) # (!idex_ifaluop_o_1 & (((\myif.out[5]~64_combout ))))

	.dataa(\Add1~10_combout ),
	.datab(\out~23_combout ),
	.datac(idex_ifaluop_o_1),
	.datad(\myif.out[5]~64_combout ),
	.cin(gnd),
	.combout(\myif.out[5]~65_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[5]~65 .lut_mask = 16'h3FA0;
defparam \myif.out[5]~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N0
cycloneive_lcell_comb \ShiftLeft0~89 (
// Equation(s):
// \ShiftLeft0~89_combout  = (!\port_b~14_combout  & ((\port_b~10_combout  & (\ShiftLeft0~85_combout )) # (!\port_b~10_combout  & ((\ShiftLeft0~82_combout )))))

	.dataa(port_b7),
	.datab(\ShiftLeft0~85_combout ),
	.datac(port_b6),
	.datad(\ShiftLeft0~82_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~89_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~89 .lut_mask = 16'h4540;
defparam \ShiftLeft0~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N26
cycloneive_lcell_comb \myif.out[7]~75 (
// Equation(s):
// \myif.out[7]~75_combout  = (idex_ifaluop_o_2 & ((\port_b~47_combout ) # ((\port_b~0_combout  & fuifrtReplace_7))))

	.dataa(port_b),
	.datab(idex_ifaluop_o_2),
	.datac(port_b37),
	.datad(fuifrtReplace_7),
	.cin(gnd),
	.combout(\myif.out[7]~75_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[7]~75 .lut_mask = 16'hC8C0;
defparam \myif.out[7]~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N0
cycloneive_lcell_comb \myif.out[7]~76 (
// Equation(s):
// \myif.out[7]~76_combout  = (idex_ifaluop_o_1 & (\Add0~14_combout  & ((!\myif.out[7]~75_combout ) # (!\rdat1[7]~13_combout )))) # (!idex_ifaluop_o_1 & (\rdat1[7]~13_combout  & ((\myif.out[7]~75_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(rdat1_7),
	.datac(\Add0~14_combout ),
	.datad(\myif.out[7]~75_combout ),
	.cin(gnd),
	.combout(\myif.out[7]~76_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[7]~76 .lut_mask = 16'h64A0;
defparam \myif.out[7]~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N22
cycloneive_lcell_comb \myif.out[7]~77 (
// Equation(s):
// \myif.out[7]~77_combout  = (\ShiftLeft0~89_combout  & ((idex_ifaluop_o_2 & ((\myif.out[7]~76_combout ))) # (!idex_ifaluop_o_2 & (\myif.out[7]~74_combout )))) # (!\ShiftLeft0~89_combout  & (((\myif.out[7]~76_combout ))))

	.dataa(\myif.out[7]~74_combout ),
	.datab(\ShiftLeft0~89_combout ),
	.datac(idex_ifaluop_o_2),
	.datad(\myif.out[7]~76_combout ),
	.cin(gnd),
	.combout(\myif.out[7]~77_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[7]~77 .lut_mask = 16'hFB08;
defparam \myif.out[7]~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N6
cycloneive_lcell_comb \myif.out[7]~78 (
// Equation(s):
// \myif.out[7]~78_combout  = \rdat1[7]~13_combout  $ (((\port_b~47_combout ) # ((fuifrtReplace_7 & \port_b~0_combout ))))

	.dataa(port_b37),
	.datab(fuifrtReplace_7),
	.datac(port_b),
	.datad(rdat1_7),
	.cin(gnd),
	.combout(\myif.out[7]~78_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[7]~78 .lut_mask = 16'h15EA;
defparam \myif.out[7]~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N20
cycloneive_lcell_comb \myif.out[7]~79 (
// Equation(s):
// \myif.out[7]~79_combout  = (idex_ifaluop_o_2 & (((\myif.out[7]~78_combout )) # (!idex_ifaluop_o_1))) # (!idex_ifaluop_o_2 & (((\myif.out[7]~76_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(idex_ifaluop_o_2),
	.datac(\myif.out[7]~78_combout ),
	.datad(\myif.out[7]~76_combout ),
	.cin(gnd),
	.combout(\myif.out[7]~79_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[7]~79 .lut_mask = 16'hF7C4;
defparam \myif.out[7]~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N26
cycloneive_lcell_comb \myif.out[7]~80 (
// Equation(s):
// \myif.out[7]~80_combout  = (\myif.out[13]~23_combout  & (\myif.out[7]~77_combout )) # (!\myif.out[13]~23_combout  & ((\myif.out[7]~79_combout )))

	.dataa(gnd),
	.datab(\myif.out[13]~23_combout ),
	.datac(\myif.out[7]~77_combout ),
	.datad(\myif.out[7]~79_combout ),
	.cin(gnd),
	.combout(\myif.out[7]~80_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[7]~80 .lut_mask = 16'hF3C0;
defparam \myif.out[7]~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N20
cycloneive_lcell_comb \out~26 (
// Equation(s):
// \out~26_combout  = (\port_b~47_combout ) # ((\rdat1[7]~13_combout ) # ((fuifrtReplace_7 & \port_b~0_combout )))

	.dataa(port_b37),
	.datab(fuifrtReplace_7),
	.datac(port_b),
	.datad(rdat1_7),
	.cin(gnd),
	.combout(\out~26_combout ),
	.cout());
// synopsys translate_off
defparam \out~26 .lut_mask = 16'hFFEA;
defparam \out~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N28
cycloneive_lcell_comb \ShiftRight0~80 (
// Equation(s):
// \ShiftRight0~80_combout  = (\port_b~4_combout  & (\ShiftRight0~10_combout )) # (!\port_b~4_combout  & ((\ShiftRight0~12_combout )))

	.dataa(gnd),
	.datab(port_b2),
	.datac(\ShiftRight0~10_combout ),
	.datad(\ShiftRight0~12_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~80 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N30
cycloneive_lcell_comb \ShiftRight0~86 (
// Equation(s):
// \ShiftRight0~86_combout  = (\port_b~4_combout  & (\ShiftRight0~13_combout )) # (!\port_b~4_combout  & ((\ShiftRight0~5_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~13_combout ),
	.datac(port_b2),
	.datad(\ShiftRight0~5_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~86 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N26
cycloneive_lcell_comb \ShiftRight0~81 (
// Equation(s):
// \ShiftRight0~81_combout  = (\port_b~7_combout  & ((\port_b~4_combout  & ((\rdat1[22]~51_combout ))) # (!\port_b~4_combout  & (\rdat1[20]~57_combout ))))

	.dataa(rdat1_20),
	.datab(port_b4),
	.datac(port_b2),
	.datad(rdat1_22),
	.cin(gnd),
	.combout(\ShiftRight0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~81 .lut_mask = 16'hC808;
defparam \ShiftRight0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N12
cycloneive_lcell_comb \ShiftRight0~33 (
// Equation(s):
// \ShiftRight0~33_combout  = (\port_b~4_combout  & (\rdat1[21]~55_combout )) # (!\port_b~4_combout  & ((\rdat1[19]~61_combout )))

	.dataa(gnd),
	.datab(rdat1_21),
	.datac(port_b2),
	.datad(rdat1_19),
	.cin(gnd),
	.combout(\ShiftRight0~33_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~33 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N8
cycloneive_lcell_comb \ShiftRight0~82 (
// Equation(s):
// \ShiftRight0~82_combout  = (\ShiftRight0~81_combout ) # ((!\port_b~7_combout  & \ShiftRight0~33_combout ))

	.dataa(gnd),
	.datab(port_b4),
	.datac(\ShiftRight0~81_combout ),
	.datad(\ShiftRight0~33_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~82 .lut_mask = 16'hF3F0;
defparam \ShiftRight0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N12
cycloneive_lcell_comb \ShiftRight0~83 (
// Equation(s):
// \ShiftRight0~83_combout  = (!\port_b~7_combout  & ((\port_b~4_combout  & ((\rdat1[17]~63_combout ))) # (!\port_b~4_combout  & (\rdat1[15]~21_combout ))))

	.dataa(rdat1_15),
	.datab(port_b4),
	.datac(rdat1_17),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftRight0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~83 .lut_mask = 16'h3022;
defparam \ShiftRight0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N2
cycloneive_lcell_comb \ShiftRight0~84 (
// Equation(s):
// \ShiftRight0~84_combout  = (\port_b~7_combout  & ((\port_b~4_combout  & ((\rdat1[18]~59_combout ))) # (!\port_b~4_combout  & (\rdat1[16]~19_combout ))))

	.dataa(port_b2),
	.datab(rdat1_16),
	.datac(rdat1_18),
	.datad(port_b4),
	.cin(gnd),
	.combout(\ShiftRight0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~84 .lut_mask = 16'hE400;
defparam \ShiftRight0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N18
cycloneive_lcell_comb \ShiftRight0~85 (
// Equation(s):
// \ShiftRight0~85_combout  = (\port_b~10_combout  & (\ShiftRight0~82_combout )) # (!\port_b~10_combout  & (((\ShiftRight0~83_combout ) # (\ShiftRight0~84_combout ))))

	.dataa(port_b6),
	.datab(\ShiftRight0~82_combout ),
	.datac(\ShiftRight0~83_combout ),
	.datad(\ShiftRight0~84_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~85_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~85 .lut_mask = 16'hDDD8;
defparam \ShiftRight0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N20
cycloneive_lcell_comb \myif.out[7]~69 (
// Equation(s):
// \myif.out[7]~69_combout  = (\myif.out[5]~16_combout  & ((\myif.out[5]~17_combout ) # ((\ShiftRight0~85_combout )))) # (!\myif.out[5]~16_combout  & (!\myif.out[5]~17_combout  & (\ShiftRight0~86_combout )))

	.dataa(\myif.out[5]~16_combout ),
	.datab(\myif.out[5]~17_combout ),
	.datac(\ShiftRight0~86_combout ),
	.datad(\ShiftRight0~85_combout ),
	.cin(gnd),
	.combout(\myif.out[7]~69_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[7]~69 .lut_mask = 16'hBA98;
defparam \myif.out[7]~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N6
cycloneive_lcell_comb \myif.out[7]~70 (
// Equation(s):
// \myif.out[7]~70_combout  = (\myif.out[5]~17_combout  & ((\myif.out[7]~69_combout  & (\ShiftRight0~90_combout )) # (!\myif.out[7]~69_combout  & ((\ShiftRight0~80_combout ))))) # (!\myif.out[5]~17_combout  & (((\myif.out[7]~69_combout ))))

	.dataa(\ShiftRight0~90_combout ),
	.datab(\ShiftRight0~80_combout ),
	.datac(\myif.out[5]~17_combout ),
	.datad(\myif.out[7]~69_combout ),
	.cin(gnd),
	.combout(\myif.out[7]~70_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[7]~70 .lut_mask = 16'hAFC0;
defparam \myif.out[7]~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N16
cycloneive_lcell_comb \myif.out[7]~71 (
// Equation(s):
// \myif.out[7]~71_combout  = (idex_ifaluop_o_2 & ((\out~26_combout ) # ((!\myif.out[5]~20_combout )))) # (!idex_ifaluop_o_2 & (((\myif.out[7]~70_combout  & \myif.out[5]~20_combout ))))

	.dataa(\out~26_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\myif.out[7]~70_combout ),
	.datad(\myif.out[5]~20_combout ),
	.cin(gnd),
	.combout(\myif.out[7]~71_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[7]~71 .lut_mask = 16'hB8CC;
defparam \myif.out[7]~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N18
cycloneive_lcell_comb \myif.out[7]~72 (
// Equation(s):
// \myif.out[7]~72_combout  = (idex_ifaluop_o_1 & ((\myif.out[7]~71_combout  & ((!\out~26_combout ))) # (!\myif.out[7]~71_combout  & (\Add1~14_combout )))) # (!idex_ifaluop_o_1 & (((\myif.out[7]~71_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(\Add1~14_combout ),
	.datac(\out~26_combout ),
	.datad(\myif.out[7]~71_combout ),
	.cin(gnd),
	.combout(\myif.out[7]~72_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[7]~72 .lut_mask = 16'h5F88;
defparam \myif.out[7]~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N4
cycloneive_lcell_comb \out~27 (
// Equation(s):
// \out~27_combout  = (\port_b~69_combout ) # ((\rdat1[13]~25_combout ) # ((\port_b~0_combout  & fuifrtReplace_13)))

	.dataa(port_b),
	.datab(fuifrtReplace_13),
	.datac(port_b59),
	.datad(rdat1_13),
	.cin(gnd),
	.combout(\out~27_combout ),
	.cout());
// synopsys translate_off
defparam \out~27 .lut_mask = 16'hFFF8;
defparam \out~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N8
cycloneive_lcell_comb \myif.out[13]~87 (
// Equation(s):
// \myif.out[13]~87_combout  = (idex_ifaluop_o_0 & ((idex_ifaluop_o_2) # (!idex_ifaluop_o_1)))

	.dataa(gnd),
	.datab(idex_ifaluop_o_0),
	.datac(idex_ifaluop_o_2),
	.datad(idex_ifaluop_o_1),
	.cin(gnd),
	.combout(\myif.out[13]~87_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[13]~87 .lut_mask = 16'hC0CC;
defparam \myif.out[13]~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N12
cycloneive_lcell_comb \myif.out[13]~82 (
// Equation(s):
// \myif.out[13]~82_combout  = (idex_ifaluop_o_2) # ((\port_b~17_combout ) # (\ShiftLeft0~11_combout ))

	.dataa(gnd),
	.datab(idex_ifaluop_o_2),
	.datac(port_b8),
	.datad(\ShiftLeft0~11_combout ),
	.cin(gnd),
	.combout(\myif.out[13]~82_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[13]~82 .lut_mask = 16'hFFFC;
defparam \myif.out[13]~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N26
cycloneive_lcell_comb \myif.out[13]~83 (
// Equation(s):
// \myif.out[13]~83_combout  = (idex_ifaluop_o_2) # ((\port_b~17_combout  & !\ShiftLeft0~11_combout ))

	.dataa(port_b8),
	.datab(gnd),
	.datac(idex_ifaluop_o_2),
	.datad(\ShiftLeft0~11_combout ),
	.cin(gnd),
	.combout(\myif.out[13]~83_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[13]~83 .lut_mask = 16'hF0FA;
defparam \myif.out[13]~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N30
cycloneive_lcell_comb \myif.out[13]~84 (
// Equation(s):
// \myif.out[13]~84_combout  = (idex_ifaluop_o_2) # ((\port_b~14_combout  & (!\port_b~17_combout  & !\ShiftLeft0~11_combout )))

	.dataa(port_b7),
	.datab(idex_ifaluop_o_2),
	.datac(port_b8),
	.datad(\ShiftLeft0~11_combout ),
	.cin(gnd),
	.combout(\myif.out[13]~84_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[13]~84 .lut_mask = 16'hCCCE;
defparam \myif.out[13]~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N26
cycloneive_lcell_comb \myif.out[13]~85 (
// Equation(s):
// \myif.out[13]~85_combout  = (\myif.out[13]~83_combout  & ((\myif.out[13]~84_combout  & ((\out~27_combout ))) # (!\myif.out[13]~84_combout  & (\ShiftRight0~91_combout )))) # (!\myif.out[13]~83_combout  & (((\myif.out[13]~84_combout ))))

	.dataa(\ShiftRight0~91_combout ),
	.datab(\myif.out[13]~83_combout ),
	.datac(\out~27_combout ),
	.datad(\myif.out[13]~84_combout ),
	.cin(gnd),
	.combout(\myif.out[13]~85_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[13]~85 .lut_mask = 16'hF388;
defparam \myif.out[13]~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N20
cycloneive_lcell_comb \myif.out[13]~86 (
// Equation(s):
// \myif.out[13]~86_combout  = (\myif.out[13]~82_combout  & (((\myif.out[13]~85_combout )))) # (!\myif.out[13]~82_combout  & ((\myif.out[13]~85_combout  & ((\ShiftRight0~78_combout ))) # (!\myif.out[13]~85_combout  & (\ShiftRight0~77_combout ))))

	.dataa(\myif.out[13]~82_combout ),
	.datab(\ShiftRight0~77_combout ),
	.datac(\myif.out[13]~85_combout ),
	.datad(\ShiftRight0~78_combout ),
	.cin(gnd),
	.combout(\myif.out[13]~86_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[13]~86 .lut_mask = 16'hF4A4;
defparam \myif.out[13]~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N14
cycloneive_lcell_comb \myif.out[13]~88 (
// Equation(s):
// \myif.out[13]~88_combout  = (idex_ifaluop_o_1 & idex_ifaluop_o_0)

	.dataa(gnd),
	.datab(idex_ifaluop_o_1),
	.datac(gnd),
	.datad(idex_ifaluop_o_0),
	.cin(gnd),
	.combout(\myif.out[13]~88_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[13]~88 .lut_mask = 16'hCC00;
defparam \myif.out[13]~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N22
cycloneive_lcell_comb \out~28 (
// Equation(s):
// \out~28_combout  = \rdat1[13]~25_combout  $ (((\port_b~69_combout ) # ((\port_b~0_combout  & fuifrtReplace_13))))

	.dataa(port_b),
	.datab(fuifrtReplace_13),
	.datac(port_b59),
	.datad(rdat1_13),
	.cin(gnd),
	.combout(\out~28_combout ),
	.cout());
// synopsys translate_off
defparam \out~28 .lut_mask = 16'h07F8;
defparam \out~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N2
cycloneive_lcell_comb \out~29 (
// Equation(s):
// \out~29_combout  = (\rdat1[13]~25_combout  & ((\port_b~69_combout ) # ((fuifrtReplace_13 & \port_b~0_combout ))))

	.dataa(fuifrtReplace_13),
	.datab(port_b),
	.datac(port_b59),
	.datad(rdat1_13),
	.cin(gnd),
	.combout(\out~29_combout ),
	.cout());
// synopsys translate_off
defparam \out~29 .lut_mask = 16'hF800;
defparam \out~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N20
cycloneive_lcell_comb \ShiftLeft0~90 (
// Equation(s):
// \ShiftLeft0~90_combout  = (\port_b~10_combout  & ((\ShiftLeft0~71_combout ))) # (!\port_b~10_combout  & (\ShiftLeft0~57_combout ))

	.dataa(gnd),
	.datab(port_b6),
	.datac(\ShiftLeft0~57_combout ),
	.datad(\ShiftLeft0~71_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~90_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~90 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N14
cycloneive_lcell_comb \ShiftLeft0~91 (
// Equation(s):
// \ShiftLeft0~91_combout  = (\port_b~14_combout  & (\ShiftLeft0~87_combout )) # (!\port_b~14_combout  & ((\ShiftLeft0~90_combout )))

	.dataa(port_b7),
	.datab(gnd),
	.datac(\ShiftLeft0~87_combout ),
	.datad(\ShiftLeft0~90_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~91_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~91 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N2
cycloneive_lcell_comb \myif.out[13]~89 (
// Equation(s):
// \myif.out[13]~89_combout  = (idex_ifaluop_o_2 & (((\out~29_combout )) # (!\myif.out[13]~23_combout ))) # (!idex_ifaluop_o_2 & (\myif.out[13]~23_combout  & ((\ShiftLeft0~91_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\myif.out[13]~23_combout ),
	.datac(\out~29_combout ),
	.datad(\ShiftLeft0~91_combout ),
	.cin(gnd),
	.combout(\myif.out[13]~89_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[13]~89 .lut_mask = 16'hE6A2;
defparam \myif.out[13]~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N20
cycloneive_lcell_comb \myif.out[13]~90 (
// Equation(s):
// \myif.out[13]~90_combout  = (idex_ifaluop_o_1 & ((\myif.out[13]~89_combout  & ((\out~28_combout ))) # (!\myif.out[13]~89_combout  & (\Add0~26_combout )))) # (!idex_ifaluop_o_1 & (((\myif.out[13]~89_combout ))))

	.dataa(\Add0~26_combout ),
	.datab(idex_ifaluop_o_1),
	.datac(\out~28_combout ),
	.datad(\myif.out[13]~89_combout ),
	.cin(gnd),
	.combout(\myif.out[13]~90_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[13]~90 .lut_mask = 16'hF388;
defparam \myif.out[13]~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N18
cycloneive_lcell_comb \myif.out[13]~91 (
// Equation(s):
// \myif.out[13]~91_combout  = (\myif.out[13]~88_combout  & ((\Add1~26_combout ) # ((\myif.out[13]~87_combout )))) # (!\myif.out[13]~88_combout  & (((!\myif.out[13]~87_combout  & \myif.out[13]~90_combout ))))

	.dataa(\myif.out[13]~88_combout ),
	.datab(\Add1~26_combout ),
	.datac(\myif.out[13]~87_combout ),
	.datad(\myif.out[13]~90_combout ),
	.cin(gnd),
	.combout(\myif.out[13]~91_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[13]~91 .lut_mask = 16'hADA8;
defparam \myif.out[13]~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N30
cycloneive_lcell_comb \out~30 (
// Equation(s):
// \out~30_combout  = (\rdat1[9]~33_combout ) # ((\port_b~59_combout ) # ((fuifrtReplace_9 & \port_b~0_combout )))

	.dataa(fuifrtReplace_9),
	.datab(rdat1_9),
	.datac(port_b),
	.datad(port_b49),
	.cin(gnd),
	.combout(\out~30_combout ),
	.cout());
// synopsys translate_off
defparam \out~30 .lut_mask = 16'hFFEC;
defparam \out~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N30
cycloneive_lcell_comb \myif.out[9]~93 (
// Equation(s):
// \myif.out[9]~93_combout  = (\myif.out[13]~84_combout  & ((\out~30_combout ) # ((!\myif.out[13]~83_combout )))) # (!\myif.out[13]~84_combout  & (((\ShiftRight0~72_combout  & \myif.out[13]~83_combout ))))

	.dataa(\myif.out[13]~84_combout ),
	.datab(\out~30_combout ),
	.datac(\ShiftRight0~72_combout ),
	.datad(\myif.out[13]~83_combout ),
	.cin(gnd),
	.combout(\myif.out[9]~93_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[9]~93 .lut_mask = 16'hD8AA;
defparam \myif.out[9]~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N8
cycloneive_lcell_comb \myif.out[9]~94 (
// Equation(s):
// \myif.out[9]~94_combout  = (\myif.out[13]~82_combout  & (((\myif.out[9]~93_combout )))) # (!\myif.out[13]~82_combout  & ((\myif.out[9]~93_combout  & ((\ShiftRight0~29_combout ))) # (!\myif.out[9]~93_combout  & (\ShiftRight0~15_combout ))))

	.dataa(\myif.out[13]~82_combout ),
	.datab(\ShiftRight0~15_combout ),
	.datac(\myif.out[9]~93_combout ),
	.datad(\ShiftRight0~29_combout ),
	.cin(gnd),
	.combout(\myif.out[9]~94_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[9]~94 .lut_mask = 16'hF4A4;
defparam \myif.out[9]~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N12
cycloneive_lcell_comb \out~32 (
// Equation(s):
// \out~32_combout  = (\rdat1[9]~33_combout  & ((\port_b~59_combout ) # ((fuifrtReplace_9 & \port_b~0_combout ))))

	.dataa(port_b49),
	.datab(fuifrtReplace_9),
	.datac(rdat1_9),
	.datad(port_b),
	.cin(gnd),
	.combout(\out~32_combout ),
	.cout());
// synopsys translate_off
defparam \out~32 .lut_mask = 16'hE0A0;
defparam \out~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N14
cycloneive_lcell_comb \myif.out[9]~95 (
// Equation(s):
// \myif.out[9]~95_combout  = (idex_ifaluop_o_2 & (((\out~32_combout )) # (!\myif.out[13]~23_combout ))) # (!idex_ifaluop_o_2 & (\myif.out[13]~23_combout  & ((\ShiftLeft0~73_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\myif.out[13]~23_combout ),
	.datac(\out~32_combout ),
	.datad(\ShiftLeft0~73_combout ),
	.cin(gnd),
	.combout(\myif.out[9]~95_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[9]~95 .lut_mask = 16'hE6A2;
defparam \myif.out[9]~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N8
cycloneive_lcell_comb \out~31 (
// Equation(s):
// \out~31_combout  = \rdat1[9]~33_combout  $ (((\port_b~59_combout ) # ((fuifrtReplace_9 & \port_b~0_combout ))))

	.dataa(fuifrtReplace_9),
	.datab(rdat1_9),
	.datac(port_b),
	.datad(port_b49),
	.cin(gnd),
	.combout(\out~31_combout ),
	.cout());
// synopsys translate_off
defparam \out~31 .lut_mask = 16'h336C;
defparam \out~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N0
cycloneive_lcell_comb \myif.out[9]~96 (
// Equation(s):
// \myif.out[9]~96_combout  = (idex_ifaluop_o_1 & ((\myif.out[9]~95_combout  & ((\out~31_combout ))) # (!\myif.out[9]~95_combout  & (\Add0~18_combout )))) # (!idex_ifaluop_o_1 & (((\myif.out[9]~95_combout ))))

	.dataa(\Add0~18_combout ),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[9]~95_combout ),
	.datad(\out~31_combout ),
	.cin(gnd),
	.combout(\myif.out[9]~96_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[9]~96 .lut_mask = 16'hF838;
defparam \myif.out[9]~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N10
cycloneive_lcell_comb \myif.out[9]~97 (
// Equation(s):
// \myif.out[9]~97_combout  = (\myif.out[13]~88_combout  & (\myif.out[13]~87_combout )) # (!\myif.out[13]~88_combout  & ((\myif.out[13]~87_combout  & (\myif.out[9]~94_combout )) # (!\myif.out[13]~87_combout  & ((\myif.out[9]~96_combout )))))

	.dataa(\myif.out[13]~88_combout ),
	.datab(\myif.out[13]~87_combout ),
	.datac(\myif.out[9]~94_combout ),
	.datad(\myif.out[9]~96_combout ),
	.cin(gnd),
	.combout(\myif.out[9]~97_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[9]~97 .lut_mask = 16'hD9C8;
defparam \myif.out[9]~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N14
cycloneive_lcell_comb \ShiftRight0~40 (
// Equation(s):
// \ShiftRight0~40_combout  = (\port_b~7_combout  & ((\rdat1[11]~29_combout ))) # (!\port_b~7_combout  & (\rdat1[10]~31_combout ))

	.dataa(port_b4),
	.datab(rdat1_10),
	.datac(gnd),
	.datad(rdat1_11),
	.cin(gnd),
	.combout(\ShiftRight0~40_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~40 .lut_mask = 16'hEE44;
defparam \ShiftRight0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N18
cycloneive_lcell_comb \ShiftRight0~42 (
// Equation(s):
// \ShiftRight0~42_combout  = (\port_b~7_combout  & ((\rdat1[9]~33_combout ))) # (!\port_b~7_combout  & (\rdat1[8]~11_combout ))

	.dataa(port_b4),
	.datab(gnd),
	.datac(rdat1_8),
	.datad(rdat1_9),
	.cin(gnd),
	.combout(\ShiftRight0~42_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~42 .lut_mask = 16'hFA50;
defparam \ShiftRight0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N12
cycloneive_lcell_comb \ShiftRight0~54 (
// Equation(s):
// \ShiftRight0~54_combout  = (\port_b~4_combout  & (\ShiftRight0~40_combout )) # (!\port_b~4_combout  & ((\ShiftRight0~42_combout )))

	.dataa(gnd),
	.datab(port_b2),
	.datac(\ShiftRight0~40_combout ),
	.datad(\ShiftRight0~42_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~54 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N20
cycloneive_lcell_comb \ShiftRight0~92 (
// Equation(s):
// \ShiftRight0~92_combout  = (\port_b~10_combout  & (\ShiftRight0~57_combout )) # (!\port_b~10_combout  & ((\ShiftRight0~54_combout )))

	.dataa(\ShiftRight0~57_combout ),
	.datab(gnd),
	.datac(port_b6),
	.datad(\ShiftRight0~54_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~92_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~92 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N30
cycloneive_lcell_comb \ShiftRight0~93 (
// Equation(s):
// \ShiftRight0~93_combout  = (\port_b~10_combout  & (\ShiftRight0~64_combout )) # (!\port_b~10_combout  & ((\ShiftRight0~56_combout )))

	.dataa(gnd),
	.datab(port_b6),
	.datac(\ShiftRight0~64_combout ),
	.datad(\ShiftRight0~56_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~93_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~93 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N24
cycloneive_lcell_comb \myif.out[8]~99 (
// Equation(s):
// \myif.out[8]~99_combout  = (\myif.out[13]~83_combout  & ((\myif.out[13]~84_combout  & (\out~33_combout )) # (!\myif.out[13]~84_combout  & ((\ShiftRight0~69_combout ))))) # (!\myif.out[13]~83_combout  & (((\myif.out[13]~84_combout ))))

	.dataa(\out~33_combout ),
	.datab(\myif.out[13]~83_combout ),
	.datac(\myif.out[13]~84_combout ),
	.datad(\ShiftRight0~69_combout ),
	.cin(gnd),
	.combout(\myif.out[8]~99_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[8]~99 .lut_mask = 16'hBCB0;
defparam \myif.out[8]~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N6
cycloneive_lcell_comb \myif.out[8]~100 (
// Equation(s):
// \myif.out[8]~100_combout  = (\myif.out[13]~82_combout  & (((\myif.out[8]~99_combout )))) # (!\myif.out[13]~82_combout  & ((\myif.out[8]~99_combout  & ((\ShiftRight0~93_combout ))) # (!\myif.out[8]~99_combout  & (\ShiftRight0~92_combout ))))

	.dataa(\ShiftRight0~92_combout ),
	.datab(\myif.out[13]~82_combout ),
	.datac(\ShiftRight0~93_combout ),
	.datad(\myif.out[8]~99_combout ),
	.cin(gnd),
	.combout(\myif.out[8]~100_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[8]~100 .lut_mask = 16'hFC22;
defparam \myif.out[8]~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N8
cycloneive_lcell_comb \out~35 (
// Equation(s):
// \out~35_combout  = (\rdat1[8]~11_combout  & ((\port_b~49_combout ) # ((fuifrtReplace_8 & \port_b~0_combout ))))

	.dataa(fuifrtReplace_8),
	.datab(port_b39),
	.datac(port_b),
	.datad(rdat1_8),
	.cin(gnd),
	.combout(\out~35_combout ),
	.cout());
// synopsys translate_off
defparam \out~35 .lut_mask = 16'hEC00;
defparam \out~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N22
cycloneive_lcell_comb \myif.out[8]~101 (
// Equation(s):
// \myif.out[8]~101_combout  = (idex_ifaluop_o_2 & ((\out~35_combout ) # ((!\myif.out[13]~23_combout )))) # (!idex_ifaluop_o_2 & (((\ShiftLeft0~40_combout  & \myif.out[13]~23_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\out~35_combout ),
	.datac(\ShiftLeft0~40_combout ),
	.datad(\myif.out[13]~23_combout ),
	.cin(gnd),
	.combout(\myif.out[8]~101_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[8]~101 .lut_mask = 16'hD8AA;
defparam \myif.out[8]~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N0
cycloneive_lcell_comb \out~34 (
// Equation(s):
// \out~34_combout  = \rdat1[8]~11_combout  $ (((\port_b~49_combout ) # ((\port_b~0_combout  & fuifrtReplace_8))))

	.dataa(rdat1_8),
	.datab(port_b),
	.datac(fuifrtReplace_8),
	.datad(port_b39),
	.cin(gnd),
	.combout(\out~34_combout ),
	.cout());
// synopsys translate_off
defparam \out~34 .lut_mask = 16'h556A;
defparam \out~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N28
cycloneive_lcell_comb \myif.out[8]~102 (
// Equation(s):
// \myif.out[8]~102_combout  = (idex_ifaluop_o_1 & ((\myif.out[8]~101_combout  & ((\out~34_combout ))) # (!\myif.out[8]~101_combout  & (\Add0~16_combout )))) # (!idex_ifaluop_o_1 & (((\myif.out[8]~101_combout ))))

	.dataa(\Add0~16_combout ),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[8]~101_combout ),
	.datad(\out~34_combout ),
	.cin(gnd),
	.combout(\myif.out[8]~102_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[8]~102 .lut_mask = 16'hF838;
defparam \myif.out[8]~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N26
cycloneive_lcell_comb \myif.out[8]~103 (
// Equation(s):
// \myif.out[8]~103_combout  = (\myif.out[13]~88_combout  & ((\myif.out[13]~87_combout ) # ((\Add1~16_combout )))) # (!\myif.out[13]~88_combout  & (!\myif.out[13]~87_combout  & ((\myif.out[8]~102_combout ))))

	.dataa(\myif.out[13]~88_combout ),
	.datab(\myif.out[13]~87_combout ),
	.datac(\Add1~16_combout ),
	.datad(\myif.out[8]~102_combout ),
	.cin(gnd),
	.combout(\myif.out[8]~103_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[8]~103 .lut_mask = 16'hB9A8;
defparam \myif.out[8]~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N10
cycloneive_lcell_comb \out~33 (
// Equation(s):
// \out~33_combout  = (\port_b~49_combout ) # ((\rdat1[8]~11_combout ) # ((\port_b~0_combout  & fuifrtReplace_8)))

	.dataa(port_b),
	.datab(fuifrtReplace_8),
	.datac(port_b39),
	.datad(rdat1_8),
	.cin(gnd),
	.combout(\out~33_combout ),
	.cout());
// synopsys translate_off
defparam \out~33 .lut_mask = 16'hFFF8;
defparam \out~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N6
cycloneive_lcell_comb \out~36 (
// Equation(s):
// \out~36_combout  = (\port_b~61_combout ) # ((\rdat1[14]~23_combout ) # ((\port_b~0_combout  & fuifrtReplace_14)))

	.dataa(port_b),
	.datab(port_b51),
	.datac(rdat1_14),
	.datad(fuifrtReplace_14),
	.cin(gnd),
	.combout(\out~36_combout ),
	.cout());
// synopsys translate_off
defparam \out~36 .lut_mask = 16'hFEFC;
defparam \out~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N12
cycloneive_lcell_comb \out~37 (
// Equation(s):
// \out~37_combout  = \rdat1[14]~23_combout  $ (((\port_b~61_combout ) # ((\port_b~0_combout  & fuifrtReplace_14))))

	.dataa(port_b),
	.datab(port_b51),
	.datac(rdat1_14),
	.datad(fuifrtReplace_14),
	.cin(gnd),
	.combout(\out~37_combout ),
	.cout());
// synopsys translate_off
defparam \out~37 .lut_mask = 16'h1E3C;
defparam \out~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N26
cycloneive_lcell_comb \out~38 (
// Equation(s):
// \out~38_combout  = (\rdat1[14]~23_combout  & ((\port_b~61_combout ) # ((\port_b~0_combout  & fuifrtReplace_14))))

	.dataa(port_b),
	.datab(port_b51),
	.datac(rdat1_14),
	.datad(fuifrtReplace_14),
	.cin(gnd),
	.combout(\out~38_combout ),
	.cout());
// synopsys translate_off
defparam \out~38 .lut_mask = 16'hE0C0;
defparam \out~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N28
cycloneive_lcell_comb \ShiftLeft0~92 (
// Equation(s):
// \ShiftLeft0~92_combout  = (\port_b~10_combout  & (\ShiftLeft0~16_combout )) # (!\port_b~10_combout  & ((\ShiftLeft0~19_combout )))

	.dataa(gnd),
	.datab(port_b6),
	.datac(\ShiftLeft0~16_combout ),
	.datad(\ShiftLeft0~19_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~92_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~92 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N18
cycloneive_lcell_comb \ShiftLeft0~93 (
// Equation(s):
// \ShiftLeft0~93_combout  = (\port_b~10_combout  & ((\ShiftLeft0~52_combout ))) # (!\port_b~10_combout  & (\ShiftLeft0~45_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~45_combout ),
	.datac(port_b6),
	.datad(\ShiftLeft0~52_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~93_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~93 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N28
cycloneive_lcell_comb \ShiftLeft0~94 (
// Equation(s):
// \ShiftLeft0~94_combout  = (\port_b~14_combout  & (\ShiftLeft0~92_combout )) # (!\port_b~14_combout  & ((\ShiftLeft0~93_combout )))

	.dataa(gnd),
	.datab(port_b7),
	.datac(\ShiftLeft0~92_combout ),
	.datad(\ShiftLeft0~93_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~94_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~94 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N2
cycloneive_lcell_comb \myif.out[14]~107 (
// Equation(s):
// \myif.out[14]~107_combout  = (\myif.out[13]~23_combout  & ((idex_ifaluop_o_2 & (\out~38_combout )) # (!idex_ifaluop_o_2 & ((\ShiftLeft0~94_combout ))))) # (!\myif.out[13]~23_combout  & (idex_ifaluop_o_2))

	.dataa(\myif.out[13]~23_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\out~38_combout ),
	.datad(\ShiftLeft0~94_combout ),
	.cin(gnd),
	.combout(\myif.out[14]~107_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[14]~107 .lut_mask = 16'hE6C4;
defparam \myif.out[14]~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N16
cycloneive_lcell_comb \myif.out[14]~108 (
// Equation(s):
// \myif.out[14]~108_combout  = (idex_ifaluop_o_1 & ((\myif.out[14]~107_combout  & ((\out~37_combout ))) # (!\myif.out[14]~107_combout  & (\Add0~28_combout )))) # (!idex_ifaluop_o_1 & (((\myif.out[14]~107_combout ))))

	.dataa(\Add0~28_combout ),
	.datab(idex_ifaluop_o_1),
	.datac(\out~37_combout ),
	.datad(\myif.out[14]~107_combout ),
	.cin(gnd),
	.combout(\myif.out[14]~108_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[14]~108 .lut_mask = 16'hF388;
defparam \myif.out[14]~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N24
cycloneive_lcell_comb \ShiftRight0~94 (
// Equation(s):
// \ShiftRight0~94_combout  = (!\port_b~14_combout  & (\ShiftRight0~52_combout  & !\ShiftLeft0~13_combout ))

	.dataa(port_b7),
	.datab(gnd),
	.datac(\ShiftRight0~52_combout ),
	.datad(\ShiftLeft0~13_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~94_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~94 .lut_mask = 16'h0050;
defparam \ShiftRight0~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N4
cycloneive_lcell_comb \myif.out[14]~105 (
// Equation(s):
// \myif.out[14]~105_combout  = (\myif.out[13]~83_combout  & ((\myif.out[13]~84_combout  & (\out~36_combout )) # (!\myif.out[13]~84_combout  & ((\ShiftRight0~94_combout ))))) # (!\myif.out[13]~83_combout  & (((\myif.out[13]~84_combout ))))

	.dataa(\out~36_combout ),
	.datab(\ShiftRight0~94_combout ),
	.datac(\myif.out[13]~83_combout ),
	.datad(\myif.out[13]~84_combout ),
	.cin(gnd),
	.combout(\myif.out[14]~105_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[14]~105 .lut_mask = 16'hAFC0;
defparam \myif.out[14]~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N6
cycloneive_lcell_comb \myif.out[14]~106 (
// Equation(s):
// \myif.out[14]~106_combout  = (\myif.out[13]~82_combout  & (\myif.out[14]~105_combout )) # (!\myif.out[13]~82_combout  & ((\myif.out[14]~105_combout  & (\ShiftRight0~51_combout )) # (!\myif.out[14]~105_combout  & ((\ShiftRight0~38_combout )))))

	.dataa(\myif.out[13]~82_combout ),
	.datab(\myif.out[14]~105_combout ),
	.datac(\ShiftRight0~51_combout ),
	.datad(\ShiftRight0~38_combout ),
	.cin(gnd),
	.combout(\myif.out[14]~106_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[14]~106 .lut_mask = 16'hD9C8;
defparam \myif.out[14]~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N0
cycloneive_lcell_comb \myif.out[14]~109 (
// Equation(s):
// \myif.out[14]~109_combout  = (\myif.out[13]~87_combout  & ((\myif.out[13]~88_combout ) # ((\myif.out[14]~106_combout )))) # (!\myif.out[13]~87_combout  & (!\myif.out[13]~88_combout  & (\myif.out[14]~108_combout )))

	.dataa(\myif.out[13]~87_combout ),
	.datab(\myif.out[13]~88_combout ),
	.datac(\myif.out[14]~108_combout ),
	.datad(\myif.out[14]~106_combout ),
	.cin(gnd),
	.combout(\myif.out[14]~109_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[14]~109 .lut_mask = 16'hBA98;
defparam \myif.out[14]~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N8
cycloneive_lcell_comb \out~39 (
// Equation(s):
// \out~39_combout  = (\port_b~68_combout ) # ((\rdat1[12]~27_combout ) # ((\port_b~0_combout  & fuifrtReplace_12)))

	.dataa(port_b),
	.datab(port_b58),
	.datac(rdat1_12),
	.datad(fuifrtReplace_12),
	.cin(gnd),
	.combout(\out~39_combout ),
	.cout());
// synopsys translate_off
defparam \out~39 .lut_mask = 16'hFEFC;
defparam \out~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N26
cycloneive_lcell_comb \out~40 (
// Equation(s):
// \out~40_combout  = \rdat1[12]~27_combout  $ (((\port_b~68_combout ) # ((\port_b~0_combout  & fuifrtReplace_12))))

	.dataa(port_b),
	.datab(port_b58),
	.datac(rdat1_12),
	.datad(fuifrtReplace_12),
	.cin(gnd),
	.combout(\out~40_combout ),
	.cout());
// synopsys translate_off
defparam \out~40 .lut_mask = 16'h1E3C;
defparam \out~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N6
cycloneive_lcell_comb \ShiftLeft0~96 (
// Equation(s):
// \ShiftLeft0~96_combout  = (\port_b~10_combout  & ((\ShiftLeft0~38_combout ))) # (!\port_b~10_combout  & (\ShiftLeft0~27_combout ))

	.dataa(gnd),
	.datab(port_b6),
	.datac(\ShiftLeft0~27_combout ),
	.datad(\ShiftLeft0~38_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~96_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~96 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N12
cycloneive_lcell_comb \ShiftLeft0~97 (
// Equation(s):
// \ShiftLeft0~97_combout  = (\port_b~14_combout  & (\ShiftLeft0~95_combout )) # (!\port_b~14_combout  & ((\ShiftLeft0~96_combout )))

	.dataa(\ShiftLeft0~95_combout ),
	.datab(port_b7),
	.datac(gnd),
	.datad(\ShiftLeft0~96_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~97_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~97 .lut_mask = 16'hBB88;
defparam \ShiftLeft0~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N16
cycloneive_lcell_comb \out~41 (
// Equation(s):
// \out~41_combout  = (\rdat1[12]~27_combout  & ((\port_b~68_combout ) # ((\port_b~0_combout  & fuifrtReplace_12))))

	.dataa(port_b),
	.datab(port_b58),
	.datac(rdat1_12),
	.datad(fuifrtReplace_12),
	.cin(gnd),
	.combout(\out~41_combout ),
	.cout());
// synopsys translate_off
defparam \out~41 .lut_mask = 16'hE0C0;
defparam \out~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N12
cycloneive_lcell_comb \myif.out[12]~113 (
// Equation(s):
// \myif.out[12]~113_combout  = (idex_ifaluop_o_2 & (((\out~41_combout )) # (!\myif.out[13]~23_combout ))) # (!idex_ifaluop_o_2 & (\myif.out[13]~23_combout  & (\ShiftLeft0~97_combout )))

	.dataa(idex_ifaluop_o_2),
	.datab(\myif.out[13]~23_combout ),
	.datac(\ShiftLeft0~97_combout ),
	.datad(\out~41_combout ),
	.cin(gnd),
	.combout(\myif.out[12]~113_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[12]~113 .lut_mask = 16'hEA62;
defparam \myif.out[12]~113 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N10
cycloneive_lcell_comb \myif.out[12]~114 (
// Equation(s):
// \myif.out[12]~114_combout  = (idex_ifaluop_o_1 & ((\myif.out[12]~113_combout  & ((\out~40_combout ))) # (!\myif.out[12]~113_combout  & (\Add0~24_combout )))) # (!idex_ifaluop_o_1 & (((\myif.out[12]~113_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(\Add0~24_combout ),
	.datac(\out~40_combout ),
	.datad(\myif.out[12]~113_combout ),
	.cin(gnd),
	.combout(\myif.out[12]~114_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[12]~114 .lut_mask = 16'hF588;
defparam \myif.out[12]~114 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N4
cycloneive_lcell_comb \myif.out[12]~115 (
// Equation(s):
// \myif.out[12]~115_combout  = (\myif.out[13]~87_combout  & (((\myif.out[13]~88_combout )))) # (!\myif.out[13]~87_combout  & ((\myif.out[13]~88_combout  & (\Add1~24_combout )) # (!\myif.out[13]~88_combout  & ((\myif.out[12]~114_combout )))))

	.dataa(\myif.out[13]~87_combout ),
	.datab(\Add1~24_combout ),
	.datac(\myif.out[13]~88_combout ),
	.datad(\myif.out[12]~114_combout ),
	.cin(gnd),
	.combout(\myif.out[12]~115_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[12]~115 .lut_mask = 16'hE5E0;
defparam \myif.out[12]~115 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N24
cycloneive_lcell_comb \myif.out[12]~111 (
// Equation(s):
// \myif.out[12]~111_combout  = (\myif.out[13]~84_combout  & (((\out~39_combout ) # (!\myif.out[13]~83_combout )))) # (!\myif.out[13]~84_combout  & (\ShiftRight0~95_combout  & ((\myif.out[13]~83_combout ))))

	.dataa(\ShiftRight0~95_combout ),
	.datab(\out~39_combout ),
	.datac(\myif.out[13]~84_combout ),
	.datad(\myif.out[13]~83_combout ),
	.cin(gnd),
	.combout(\myif.out[12]~111_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[12]~111 .lut_mask = 16'hCAF0;
defparam \myif.out[12]~111 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N6
cycloneive_lcell_comb \myif.out[12]~112 (
// Equation(s):
// \myif.out[12]~112_combout  = (\myif.out[13]~82_combout  & (((\myif.out[12]~111_combout )))) # (!\myif.out[13]~82_combout  & ((\myif.out[12]~111_combout  & (\ShiftRight0~65_combout )) # (!\myif.out[12]~111_combout  & ((\ShiftRight0~58_combout )))))

	.dataa(\myif.out[13]~82_combout ),
	.datab(\ShiftRight0~65_combout ),
	.datac(\ShiftRight0~58_combout ),
	.datad(\myif.out[12]~111_combout ),
	.cin(gnd),
	.combout(\myif.out[12]~112_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[12]~112 .lut_mask = 16'hEE50;
defparam \myif.out[12]~112 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N28
cycloneive_lcell_comb \out~42 (
// Equation(s):
// \out~42_combout  = (\port_b~62_combout ) # ((\rdat1[15]~21_combout ) # ((\port_b~0_combout  & fuifrtReplace_15)))

	.dataa(port_b),
	.datab(port_b52),
	.datac(rdat1_15),
	.datad(fuifrtReplace_15),
	.cin(gnd),
	.combout(\out~42_combout ),
	.cout());
// synopsys translate_off
defparam \out~42 .lut_mask = 16'hFEFC;
defparam \out~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N18
cycloneive_lcell_comb \ShiftRight0~87 (
// Equation(s):
// \ShiftRight0~87_combout  = (\port_b~7_combout  & ((\port_b~4_combout  & ((\rdat1[26]~43_combout ))) # (!\port_b~4_combout  & (\rdat1[24]~49_combout ))))

	.dataa(rdat1_24),
	.datab(rdat1_26),
	.datac(port_b4),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftRight0~87_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~87 .lut_mask = 16'hC0A0;
defparam \ShiftRight0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N16
cycloneive_lcell_comb \ShiftRight0~88 (
// Equation(s):
// \ShiftRight0~88_combout  = (\ShiftRight0~87_combout ) # ((!\port_b~7_combout  & \ShiftRight0~49_combout ))

	.dataa(gnd),
	.datab(port_b4),
	.datac(\ShiftRight0~49_combout ),
	.datad(\ShiftRight0~87_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~88_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~88 .lut_mask = 16'hFF30;
defparam \ShiftRight0~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N24
cycloneive_lcell_comb \ShiftRight0~89 (
// Equation(s):
// \ShiftRight0~89_combout  = (\port_b~10_combout  & ((\ShiftRight0~75_combout ))) # (!\port_b~10_combout  & (\ShiftRight0~88_combout ))

	.dataa(gnd),
	.datab(port_b6),
	.datac(\ShiftRight0~88_combout ),
	.datad(\ShiftRight0~75_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~89_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~89 .lut_mask = 16'hFC30;
defparam \ShiftRight0~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N12
cycloneive_lcell_comb \ShiftRight0~73 (
// Equation(s):
// \ShiftRight0~73_combout  = (!\port_b~7_combout  & (\rdat1[31]~35_combout  & !\port_b~4_combout ))

	.dataa(gnd),
	.datab(port_b4),
	.datac(rdat1_311),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftRight0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~73 .lut_mask = 16'h0030;
defparam \ShiftRight0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N16
cycloneive_lcell_comb \ShiftRight0~96 (
// Equation(s):
// \ShiftRight0~96_combout  = (!\port_b~10_combout  & (!\port_b~14_combout  & \ShiftRight0~73_combout ))

	.dataa(gnd),
	.datab(port_b6),
	.datac(port_b7),
	.datad(\ShiftRight0~73_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~96_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~96 .lut_mask = 16'h0300;
defparam \ShiftRight0~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N6
cycloneive_lcell_comb \myif.out[15]~117 (
// Equation(s):
// \myif.out[15]~117_combout  = (\myif.out[13]~84_combout  & ((\out~42_combout ) # ((!\myif.out[13]~83_combout )))) # (!\myif.out[13]~84_combout  & (((\ShiftRight0~96_combout  & \myif.out[13]~83_combout ))))

	.dataa(\out~42_combout ),
	.datab(\ShiftRight0~96_combout ),
	.datac(\myif.out[13]~84_combout ),
	.datad(\myif.out[13]~83_combout ),
	.cin(gnd),
	.combout(\myif.out[15]~117_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[15]~117 .lut_mask = 16'hACF0;
defparam \myif.out[15]~117 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N8
cycloneive_lcell_comb \myif.out[15]~118 (
// Equation(s):
// \myif.out[15]~118_combout  = (\myif.out[13]~82_combout  & (((\myif.out[15]~117_combout )))) # (!\myif.out[13]~82_combout  & ((\myif.out[15]~117_combout  & ((\ShiftRight0~89_combout ))) # (!\myif.out[15]~117_combout  & (\ShiftRight0~85_combout ))))

	.dataa(\ShiftRight0~85_combout ),
	.datab(\ShiftRight0~89_combout ),
	.datac(\myif.out[13]~82_combout ),
	.datad(\myif.out[15]~117_combout ),
	.cin(gnd),
	.combout(\myif.out[15]~118_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[15]~118 .lut_mask = 16'hFC0A;
defparam \myif.out[15]~118 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N2
cycloneive_lcell_comb \out~43 (
// Equation(s):
// \out~43_combout  = \rdat1[15]~21_combout  $ (((\port_b~62_combout ) # ((fuifrtReplace_15 & \port_b~0_combout ))))

	.dataa(fuifrtReplace_15),
	.datab(rdat1_15),
	.datac(port_b52),
	.datad(port_b),
	.cin(gnd),
	.combout(\out~43_combout ),
	.cout());
// synopsys translate_off
defparam \out~43 .lut_mask = 16'h363C;
defparam \out~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N14
cycloneive_lcell_comb \ShiftLeft0~98 (
// Equation(s):
// \ShiftLeft0~98_combout  = (\port_b~10_combout  & ((\ShiftLeft0~85_combout ))) # (!\port_b~10_combout  & (\ShiftLeft0~82_combout ))

	.dataa(\ShiftLeft0~82_combout ),
	.datab(gnd),
	.datac(\ShiftLeft0~85_combout ),
	.datad(port_b6),
	.cin(gnd),
	.combout(\ShiftLeft0~98_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~98 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N12
cycloneive_lcell_comb \ShiftLeft0~99 (
// Equation(s):
// \ShiftLeft0~99_combout  = (\port_b~10_combout  & (\ShiftLeft0~83_combout )) # (!\port_b~10_combout  & ((\ShiftLeft0~75_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~83_combout ),
	.datac(port_b6),
	.datad(\ShiftLeft0~75_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~99_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~99 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N2
cycloneive_lcell_comb \ShiftLeft0~100 (
// Equation(s):
// \ShiftLeft0~100_combout  = (\port_b~14_combout  & (\ShiftLeft0~98_combout )) # (!\port_b~14_combout  & ((\ShiftLeft0~99_combout )))

	.dataa(gnd),
	.datab(port_b7),
	.datac(\ShiftLeft0~98_combout ),
	.datad(\ShiftLeft0~99_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~100_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~100 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N10
cycloneive_lcell_comb \myif.out[15]~119 (
// Equation(s):
// \myif.out[15]~119_combout  = (idex_ifaluop_o_2 & ((\out~44_combout ) # ((!\myif.out[13]~23_combout )))) # (!idex_ifaluop_o_2 & (((\myif.out[13]~23_combout  & \ShiftLeft0~100_combout ))))

	.dataa(\out~44_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\myif.out[13]~23_combout ),
	.datad(\ShiftLeft0~100_combout ),
	.cin(gnd),
	.combout(\myif.out[15]~119_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[15]~119 .lut_mask = 16'hBC8C;
defparam \myif.out[15]~119 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N28
cycloneive_lcell_comb \myif.out[15]~120 (
// Equation(s):
// \myif.out[15]~120_combout  = (idex_ifaluop_o_1 & ((\myif.out[15]~119_combout  & (\out~43_combout )) # (!\myif.out[15]~119_combout  & ((\Add0~30_combout ))))) # (!idex_ifaluop_o_1 & (((\myif.out[15]~119_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(\out~43_combout ),
	.datac(\Add0~30_combout ),
	.datad(\myif.out[15]~119_combout ),
	.cin(gnd),
	.combout(\myif.out[15]~120_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[15]~120 .lut_mask = 16'hDDA0;
defparam \myif.out[15]~120 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N2
cycloneive_lcell_comb \myif.out[15]~121 (
// Equation(s):
// \myif.out[15]~121_combout  = (\myif.out[13]~87_combout  & ((\myif.out[13]~88_combout ) # ((\myif.out[15]~118_combout )))) # (!\myif.out[13]~87_combout  & (!\myif.out[13]~88_combout  & ((\myif.out[15]~120_combout ))))

	.dataa(\myif.out[13]~87_combout ),
	.datab(\myif.out[13]~88_combout ),
	.datac(\myif.out[15]~118_combout ),
	.datad(\myif.out[15]~120_combout ),
	.cin(gnd),
	.combout(\myif.out[15]~121_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[15]~121 .lut_mask = 16'hB9A8;
defparam \myif.out[15]~121 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N20
cycloneive_lcell_comb \out~45 (
// Equation(s):
// \out~45_combout  = (\rdat1[10]~31_combout ) # ((\port_b~64_combout ) # ((\port_b~0_combout  & fuifrtReplace_10)))

	.dataa(port_b),
	.datab(rdat1_10),
	.datac(port_b54),
	.datad(fuifrtReplace_10),
	.cin(gnd),
	.combout(\out~45_combout ),
	.cout());
// synopsys translate_off
defparam \out~45 .lut_mask = 16'hFEFC;
defparam \out~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N28
cycloneive_lcell_comb \ShiftRight0~98 (
// Equation(s):
// \ShiftRight0~98_combout  = (\port_b~10_combout  & ((\ShiftRight0~50_combout ))) # (!\port_b~10_combout  & (\ShiftRight0~34_combout ))

	.dataa(\ShiftRight0~34_combout ),
	.datab(port_b6),
	.datac(gnd),
	.datad(\ShiftRight0~50_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~98_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~98 .lut_mask = 16'hEE22;
defparam \ShiftRight0~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N0
cycloneive_lcell_comb \ShiftRight0~39 (
// Equation(s):
// \ShiftRight0~39_combout  = (\port_b~7_combout  & (\rdat1[13]~25_combout )) # (!\port_b~7_combout  & ((\rdat1[12]~27_combout )))

	.dataa(rdat1_13),
	.datab(gnd),
	.datac(rdat1_12),
	.datad(port_b4),
	.cin(gnd),
	.combout(\ShiftRight0~39_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~39 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N4
cycloneive_lcell_comb \ShiftRight0~41 (
// Equation(s):
// \ShiftRight0~41_combout  = (\port_b~4_combout  & ((\ShiftRight0~39_combout ))) # (!\port_b~4_combout  & (\ShiftRight0~40_combout ))

	.dataa(gnd),
	.datab(port_b2),
	.datac(\ShiftRight0~40_combout ),
	.datad(\ShiftRight0~39_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~41_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~41 .lut_mask = 16'hFC30;
defparam \ShiftRight0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N10
cycloneive_lcell_comb \ShiftRight0~97 (
// Equation(s):
// \ShiftRight0~97_combout  = (\port_b~10_combout  & ((\ShiftRight0~37_combout ))) # (!\port_b~10_combout  & (\ShiftRight0~41_combout ))

	.dataa(gnd),
	.datab(port_b6),
	.datac(\ShiftRight0~41_combout ),
	.datad(\ShiftRight0~37_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~97_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~97 .lut_mask = 16'hFC30;
defparam \ShiftRight0~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N0
cycloneive_lcell_comb \myif.out[10]~123 (
// Equation(s):
// \myif.out[10]~123_combout  = (\myif.out[13]~83_combout  & ((\myif.out[13]~84_combout  & ((\out~45_combout ))) # (!\myif.out[13]~84_combout  & (\ShiftRight0~71_combout )))) # (!\myif.out[13]~83_combout  & (((\myif.out[13]~84_combout ))))

	.dataa(\ShiftRight0~71_combout ),
	.datab(\out~45_combout ),
	.datac(\myif.out[13]~83_combout ),
	.datad(\myif.out[13]~84_combout ),
	.cin(gnd),
	.combout(\myif.out[10]~123_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[10]~123 .lut_mask = 16'hCFA0;
defparam \myif.out[10]~123 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N22
cycloneive_lcell_comb \myif.out[10]~124 (
// Equation(s):
// \myif.out[10]~124_combout  = (\myif.out[13]~82_combout  & (((\myif.out[10]~123_combout )))) # (!\myif.out[13]~82_combout  & ((\myif.out[10]~123_combout  & (\ShiftRight0~98_combout )) # (!\myif.out[10]~123_combout  & ((\ShiftRight0~97_combout )))))

	.dataa(\ShiftRight0~98_combout ),
	.datab(\myif.out[13]~82_combout ),
	.datac(\ShiftRight0~97_combout ),
	.datad(\myif.out[10]~123_combout ),
	.cin(gnd),
	.combout(\myif.out[10]~124_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[10]~124 .lut_mask = 16'hEE30;
defparam \myif.out[10]~124 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N14
cycloneive_lcell_comb \out~46 (
// Equation(s):
// \out~46_combout  = \rdat1[10]~31_combout  $ (((\port_b~64_combout ) # ((\port_b~0_combout  & fuifrtReplace_10))))

	.dataa(port_b),
	.datab(rdat1_10),
	.datac(port_b54),
	.datad(fuifrtReplace_10),
	.cin(gnd),
	.combout(\out~46_combout ),
	.cout());
// synopsys translate_off
defparam \out~46 .lut_mask = 16'h363C;
defparam \out~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N4
cycloneive_lcell_comb \out~47 (
// Equation(s):
// \out~47_combout  = (\rdat1[10]~31_combout  & ((\port_b~64_combout ) # ((\port_b~0_combout  & fuifrtReplace_10))))

	.dataa(port_b),
	.datab(rdat1_10),
	.datac(port_b54),
	.datad(fuifrtReplace_10),
	.cin(gnd),
	.combout(\out~47_combout ),
	.cout());
// synopsys translate_off
defparam \out~47 .lut_mask = 16'hC8C0;
defparam \out~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N10
cycloneive_lcell_comb \myif.out[10]~125 (
// Equation(s):
// \myif.out[10]~125_combout  = (idex_ifaluop_o_2 & ((\out~47_combout ) # ((!\myif.out[13]~23_combout )))) # (!idex_ifaluop_o_2 & (((\ShiftLeft0~54_combout  & \myif.out[13]~23_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\out~47_combout ),
	.datac(\ShiftLeft0~54_combout ),
	.datad(\myif.out[13]~23_combout ),
	.cin(gnd),
	.combout(\myif.out[10]~125_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[10]~125 .lut_mask = 16'hD8AA;
defparam \myif.out[10]~125 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N24
cycloneive_lcell_comb \myif.out[10]~126 (
// Equation(s):
// \myif.out[10]~126_combout  = (idex_ifaluop_o_1 & ((\myif.out[10]~125_combout  & (\out~46_combout )) # (!\myif.out[10]~125_combout  & ((\Add0~20_combout ))))) # (!idex_ifaluop_o_1 & (((\myif.out[10]~125_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(\out~46_combout ),
	.datac(\Add0~20_combout ),
	.datad(\myif.out[10]~125_combout ),
	.cin(gnd),
	.combout(\myif.out[10]~126_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[10]~126 .lut_mask = 16'hDDA0;
defparam \myif.out[10]~126 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N24
cycloneive_lcell_comb \myif.out[10]~127 (
// Equation(s):
// \myif.out[10]~127_combout  = (\myif.out[13]~87_combout  & (((\myif.out[13]~88_combout )))) # (!\myif.out[13]~87_combout  & ((\myif.out[13]~88_combout  & (\Add1~20_combout )) # (!\myif.out[13]~88_combout  & ((\myif.out[10]~126_combout )))))

	.dataa(\Add1~20_combout ),
	.datab(\myif.out[13]~87_combout ),
	.datac(\myif.out[13]~88_combout ),
	.datad(\myif.out[10]~126_combout ),
	.cin(gnd),
	.combout(\myif.out[10]~127_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[10]~127 .lut_mask = 16'hE3E0;
defparam \myif.out[10]~127 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N30
cycloneive_lcell_comb \out~48 (
// Equation(s):
// \out~48_combout  = (\rdat1[11]~29_combout ) # ((\port_b~66_combout ) # ((\port_b~0_combout  & fuifrtReplace_11)))

	.dataa(rdat1_11),
	.datab(port_b56),
	.datac(port_b),
	.datad(fuifrtReplace_11),
	.cin(gnd),
	.combout(\out~48_combout ),
	.cout());
// synopsys translate_off
defparam \out~48 .lut_mask = 16'hFEEE;
defparam \out~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N2
cycloneive_lcell_comb \ShiftRight0~100 (
// Equation(s):
// \ShiftRight0~100_combout  = (\port_b~10_combout  & (\ShiftRight0~88_combout )) # (!\port_b~10_combout  & ((\ShiftRight0~82_combout )))

	.dataa(gnd),
	.datab(port_b6),
	.datac(\ShiftRight0~88_combout ),
	.datad(\ShiftRight0~82_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~100_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~100 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N12
cycloneive_lcell_comb \myif.out[11]~129 (
// Equation(s):
// \myif.out[11]~129_combout  = (\myif.out[13]~83_combout  & ((\myif.out[13]~84_combout  & ((\out~48_combout ))) # (!\myif.out[13]~84_combout  & (\ShiftRight0~76_combout )))) # (!\myif.out[13]~83_combout  & (((\myif.out[13]~84_combout ))))

	.dataa(\ShiftRight0~76_combout ),
	.datab(\out~48_combout ),
	.datac(\myif.out[13]~83_combout ),
	.datad(\myif.out[13]~84_combout ),
	.cin(gnd),
	.combout(\myif.out[11]~129_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[11]~129 .lut_mask = 16'hCFA0;
defparam \myif.out[11]~129 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N26
cycloneive_lcell_comb \myif.out[11]~130 (
// Equation(s):
// \myif.out[11]~130_combout  = (\myif.out[13]~82_combout  & (((\myif.out[11]~129_combout )))) # (!\myif.out[13]~82_combout  & ((\myif.out[11]~129_combout  & ((\ShiftRight0~100_combout ))) # (!\myif.out[11]~129_combout  & (\ShiftRight0~99_combout ))))

	.dataa(\ShiftRight0~99_combout ),
	.datab(\ShiftRight0~100_combout ),
	.datac(\myif.out[13]~82_combout ),
	.datad(\myif.out[11]~129_combout ),
	.cin(gnd),
	.combout(\myif.out[11]~130_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[11]~130 .lut_mask = 16'hFC0A;
defparam \myif.out[11]~130 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N28
cycloneive_lcell_comb \out~50 (
// Equation(s):
// \out~50_combout  = (\rdat1[11]~29_combout  & ((\port_b~66_combout ) # ((\port_b~0_combout  & fuifrtReplace_11))))

	.dataa(port_b),
	.datab(port_b56),
	.datac(fuifrtReplace_11),
	.datad(rdat1_11),
	.cin(gnd),
	.combout(\out~50_combout ),
	.cout());
// synopsys translate_off
defparam \out~50 .lut_mask = 16'hEC00;
defparam \out~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N14
cycloneive_lcell_comb \myif.out[11]~131 (
// Equation(s):
// \myif.out[11]~131_combout  = (\myif.out[13]~23_combout  & ((idex_ifaluop_o_2 & (\out~50_combout )) # (!idex_ifaluop_o_2 & ((\ShiftLeft0~86_combout ))))) # (!\myif.out[13]~23_combout  & (idex_ifaluop_o_2))

	.dataa(\myif.out[13]~23_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\out~50_combout ),
	.datad(\ShiftLeft0~86_combout ),
	.cin(gnd),
	.combout(\myif.out[11]~131_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[11]~131 .lut_mask = 16'hE6C4;
defparam \myif.out[11]~131 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N20
cycloneive_lcell_comb \myif.out[11]~132 (
// Equation(s):
// \myif.out[11]~132_combout  = (idex_ifaluop_o_1 & ((\myif.out[11]~131_combout  & (\out~49_combout )) # (!\myif.out[11]~131_combout  & ((\Add0~22_combout ))))) # (!idex_ifaluop_o_1 & (((\myif.out[11]~131_combout ))))

	.dataa(\out~49_combout ),
	.datab(idex_ifaluop_o_1),
	.datac(\Add0~22_combout ),
	.datad(\myif.out[11]~131_combout ),
	.cin(gnd),
	.combout(\myif.out[11]~132_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[11]~132 .lut_mask = 16'hBBC0;
defparam \myif.out[11]~132 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N6
cycloneive_lcell_comb \myif.out[11]~133 (
// Equation(s):
// \myif.out[11]~133_combout  = (\myif.out[13]~88_combout  & (\myif.out[13]~87_combout )) # (!\myif.out[13]~88_combout  & ((\myif.out[13]~87_combout  & (\myif.out[11]~130_combout )) # (!\myif.out[13]~87_combout  & ((\myif.out[11]~132_combout )))))

	.dataa(\myif.out[13]~88_combout ),
	.datab(\myif.out[13]~87_combout ),
	.datac(\myif.out[11]~130_combout ),
	.datad(\myif.out[11]~132_combout ),
	.cin(gnd),
	.combout(\myif.out[11]~133_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[11]~133 .lut_mask = 16'hD9C8;
defparam \myif.out[11]~133 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N14
cycloneive_lcell_comb \myif.out[23]~135 (
// Equation(s):
// \myif.out[23]~135_combout  = (idex_ifaluop_o_1 & !idex_ifaluop_o_0)

	.dataa(gnd),
	.datab(gnd),
	.datac(idex_ifaluop_o_1),
	.datad(idex_ifaluop_o_0),
	.cin(gnd),
	.combout(\myif.out[23]~135_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~135 .lut_mask = 16'h00F0;
defparam \myif.out[23]~135 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N28
cycloneive_lcell_comb \out~51 (
// Equation(s):
// \out~51_combout  = (\rdat1[23]~53_combout  & ((\port_b~35_combout ) # ((fuifrtReplace_23 & \port_b~0_combout ))))

	.dataa(fuifrtReplace_23),
	.datab(port_b),
	.datac(rdat1_23),
	.datad(port_b25),
	.cin(gnd),
	.combout(\out~51_combout ),
	.cout());
// synopsys translate_off
defparam \out~51 .lut_mask = 16'hF080;
defparam \out~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N12
cycloneive_lcell_comb \myif.out[23]~136 (
// Equation(s):
// \myif.out[23]~136_combout  = (\myif.out[13]~83_combout  & ((\myif.out[13]~84_combout  & (\out~51_combout )) # (!\myif.out[13]~84_combout  & ((\ShiftLeft0~89_combout ))))) # (!\myif.out[13]~83_combout  & (((\myif.out[13]~84_combout ))))

	.dataa(\myif.out[13]~83_combout ),
	.datab(\out~51_combout ),
	.datac(\myif.out[13]~84_combout ),
	.datad(\ShiftLeft0~89_combout ),
	.cin(gnd),
	.combout(\myif.out[23]~136_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~136 .lut_mask = 16'hDAD0;
defparam \myif.out[23]~136 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N6
cycloneive_lcell_comb \ShiftLeft0~42 (
// Equation(s):
// \ShiftLeft0~42_combout  = (\port_b~4_combout  & (\rdat1[20]~57_combout )) # (!\port_b~4_combout  & ((\rdat1[22]~51_combout )))

	.dataa(port_b2),
	.datab(gnd),
	.datac(rdat1_20),
	.datad(rdat1_22),
	.cin(gnd),
	.combout(\ShiftLeft0~42_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~42 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N28
cycloneive_lcell_comb \ShiftLeft0~74 (
// Equation(s):
// \ShiftLeft0~74_combout  = (\port_b~7_combout  & (\ShiftLeft0~42_combout )) # (!\port_b~7_combout  & ((\ShiftLeft0~35_combout )))

	.dataa(gnd),
	.datab(port_b4),
	.datac(\ShiftLeft0~42_combout ),
	.datad(\ShiftLeft0~35_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~74 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N10
cycloneive_lcell_comb \ShiftLeft0~101 (
// Equation(s):
// \ShiftLeft0~101_combout  = (\port_b~10_combout  & (\ShiftLeft0~77_combout )) # (!\port_b~10_combout  & ((\ShiftLeft0~74_combout )))

	.dataa(\ShiftLeft0~77_combout ),
	.datab(port_b6),
	.datac(gnd),
	.datad(\ShiftLeft0~74_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~101_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~101 .lut_mask = 16'hBB88;
defparam \ShiftLeft0~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N30
cycloneive_lcell_comb \myif.out[23]~137 (
// Equation(s):
// \myif.out[23]~137_combout  = (\myif.out[23]~136_combout  & ((\ShiftLeft0~99_combout ) # ((\myif.out[13]~82_combout )))) # (!\myif.out[23]~136_combout  & (((!\myif.out[13]~82_combout  & \ShiftLeft0~101_combout ))))

	.dataa(\myif.out[23]~136_combout ),
	.datab(\ShiftLeft0~99_combout ),
	.datac(\myif.out[13]~82_combout ),
	.datad(\ShiftLeft0~101_combout ),
	.cin(gnd),
	.combout(\myif.out[23]~137_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~137 .lut_mask = 16'hADA8;
defparam \myif.out[23]~137 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N18
cycloneive_lcell_comb \myif.out[23]~150 (
// Equation(s):
// \myif.out[23]~150_combout  = (idex_ifaluop_o_0) # ((idex_ifaluop_o_2 & idex_ifaluop_o_1))

	.dataa(idex_ifaluop_o_2),
	.datab(gnd),
	.datac(idex_ifaluop_o_0),
	.datad(idex_ifaluop_o_1),
	.cin(gnd),
	.combout(\myif.out[23]~150_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~150 .lut_mask = 16'hFAF0;
defparam \myif.out[23]~150 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N14
cycloneive_lcell_comb \myif.out[23]~138 (
// Equation(s):
// \myif.out[23]~138_combout  = \rdat1[23]~53_combout  $ (((\port_b~35_combout ) # ((fuifrtReplace_23 & \port_b~0_combout ))))

	.dataa(fuifrtReplace_23),
	.datab(port_b),
	.datac(rdat1_23),
	.datad(port_b25),
	.cin(gnd),
	.combout(\myif.out[23]~138_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~138 .lut_mask = 16'h0F78;
defparam \myif.out[23]~138 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N18
cycloneive_lcell_comb \myif.out[23]~140 (
// Equation(s):
// \myif.out[23]~140_combout  = (idex_ifaluop_o_1 & (((\Add1~46_combout )))) # (!idex_ifaluop_o_1 & ((\rdat1[23]~53_combout ) # ((\myif.out[23]~138_combout ))))

	.dataa(rdat1_23),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[23]~138_combout ),
	.datad(\Add1~46_combout ),
	.cin(gnd),
	.combout(\myif.out[23]~140_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~140 .lut_mask = 16'hFE32;
defparam \myif.out[23]~140 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N12
cycloneive_lcell_comb \myif.out[23]~141 (
// Equation(s):
// \myif.out[23]~141_combout  = (\myif.out[23]~135_combout  & (\Add0~46_combout )) # (!\myif.out[23]~135_combout  & (((idex_ifaluop_o_2) # (\myif.out[23]~140_combout ))))

	.dataa(\Add0~46_combout ),
	.datab(\myif.out[23]~135_combout ),
	.datac(idex_ifaluop_o_2),
	.datad(\myif.out[23]~140_combout ),
	.cin(gnd),
	.combout(\myif.out[23]~141_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~141 .lut_mask = 16'hBBB8;
defparam \myif.out[23]~141 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N8
cycloneive_lcell_comb \myif.out[23]~151 (
// Equation(s):
// \myif.out[23]~151_combout  = (\myif.out[23]~150_combout  & ((\myif.out[23]~138_combout ) # ((!\myif.out[23]~135_combout )))) # (!\myif.out[23]~150_combout  & (((\myif.out[23]~135_combout  & \myif.out[23]~141_combout ))))

	.dataa(\myif.out[23]~150_combout ),
	.datab(\myif.out[23]~138_combout ),
	.datac(\myif.out[23]~135_combout ),
	.datad(\myif.out[23]~141_combout ),
	.cin(gnd),
	.combout(\myif.out[23]~151_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~151 .lut_mask = 16'hDA8A;
defparam \myif.out[23]~151 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N0
cycloneive_lcell_comb \myif.out[23]~139 (
// Equation(s):
// \myif.out[23]~139_combout  = (idex_ifaluop_o_2 & (((!\rdat1[23]~53_combout  & !\myif.out[23]~138_combout )) # (!idex_ifaluop_o_1))) # (!idex_ifaluop_o_2 & (((idex_ifaluop_o_1))))

	.dataa(rdat1_23),
	.datab(idex_ifaluop_o_2),
	.datac(\myif.out[23]~138_combout ),
	.datad(idex_ifaluop_o_1),
	.cin(gnd),
	.combout(\myif.out[23]~139_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~139 .lut_mask = 16'h37CC;
defparam \myif.out[23]~139 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N10
cycloneive_lcell_comb \myif.out[23]~147 (
// Equation(s):
// \myif.out[23]~147_combout  = (\myif.out[23]~142_combout  & (!idex_ifaluop_o_1)) # (!\myif.out[23]~142_combout  & ((idex_ifaluop_o_1 & (!\rdat1[23]~53_combout  & \Add1~46_combout )) # (!idex_ifaluop_o_1 & (\rdat1[23]~53_combout ))))

	.dataa(\myif.out[23]~142_combout ),
	.datab(idex_ifaluop_o_1),
	.datac(rdat1_23),
	.datad(\Add1~46_combout ),
	.cin(gnd),
	.combout(\myif.out[23]~147_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~147 .lut_mask = 16'h3632;
defparam \myif.out[23]~147 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N22
cycloneive_lcell_comb \myif.out[23]~142 (
// Equation(s):
// \myif.out[23]~142_combout  = (\port_b~35_combout ) # ((\port_b~0_combout  & fuifrtReplace_23))

	.dataa(port_b),
	.datab(gnd),
	.datac(fuifrtReplace_23),
	.datad(port_b25),
	.cin(gnd),
	.combout(\myif.out[23]~142_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~142 .lut_mask = 16'hFFA0;
defparam \myif.out[23]~142 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N20
cycloneive_lcell_comb \myif.out[23]~143 (
// Equation(s):
// \myif.out[23]~143_combout  = (\rdat1[23]~53_combout  & (idex_ifaluop_o_1 $ (((!idex_ifaluop_o_2))))) # (!\rdat1[23]~53_combout  & ((idex_ifaluop_o_1 $ (!idex_ifaluop_o_2)) # (!\myif.out[23]~142_combout )))

	.dataa(rdat1_23),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[23]~142_combout ),
	.datad(idex_ifaluop_o_2),
	.cin(gnd),
	.combout(\myif.out[23]~143_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~143 .lut_mask = 16'hCD37;
defparam \myif.out[23]~143 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N22
cycloneive_lcell_comb \ShiftRight0~90 (
// Equation(s):
// \ShiftRight0~90_combout  = (\port_b~14_combout  & (\ShiftRight0~73_combout  & (!\port_b~10_combout ))) # (!\port_b~14_combout  & (((\ShiftRight0~89_combout ))))

	.dataa(\ShiftRight0~73_combout ),
	.datab(port_b6),
	.datac(port_b7),
	.datad(\ShiftRight0~89_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~90_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~90 .lut_mask = 16'h2F20;
defparam \ShiftRight0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N26
cycloneive_lcell_comb \myif.out[23]~144 (
// Equation(s):
// \myif.out[23]~144_combout  = (\rdat1[23]~53_combout ) # ((\port_b~35_combout ) # ((\port_b~0_combout  & fuifrtReplace_23)))

	.dataa(rdat1_23),
	.datab(port_b),
	.datac(fuifrtReplace_23),
	.datad(port_b25),
	.cin(gnd),
	.combout(\myif.out[23]~144_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~144 .lut_mask = 16'hFFEA;
defparam \myif.out[23]~144 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N16
cycloneive_lcell_comb \myif.out[23]~145 (
// Equation(s):
// \myif.out[23]~145_combout  = (idex_ifaluop_o_1 & (\Add1~46_combout  & ((!\myif.out[23]~144_combout ) # (!idex_ifaluop_o_2)))) # (!idex_ifaluop_o_1 & (idex_ifaluop_o_2 & (\myif.out[23]~144_combout )))

	.dataa(idex_ifaluop_o_2),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[23]~144_combout ),
	.datad(\Add1~46_combout ),
	.cin(gnd),
	.combout(\myif.out[23]~145_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~145 .lut_mask = 16'h6C20;
defparam \myif.out[23]~145 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N10
cycloneive_lcell_comb \myif.out[23]~146 (
// Equation(s):
// \myif.out[23]~146_combout  = (\ShiftRight0~90_combout  & (\myif.out[23]~143_combout )) # (!\ShiftRight0~90_combout  & ((\myif.out[23]~145_combout )))

	.dataa(gnd),
	.datab(\myif.out[23]~143_combout ),
	.datac(\ShiftRight0~90_combout ),
	.datad(\myif.out[23]~145_combout ),
	.cin(gnd),
	.combout(\myif.out[23]~146_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~146 .lut_mask = 16'hCFC0;
defparam \myif.out[23]~146 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N16
cycloneive_lcell_comb \myif.out[23]~148 (
// Equation(s):
// \myif.out[23]~148_combout  = (idex_ifaluop_o_2 & (\myif.out[23]~147_combout )) # (!idex_ifaluop_o_2 & ((\myif.out[23]~146_combout )))

	.dataa(idex_ifaluop_o_2),
	.datab(gnd),
	.datac(\myif.out[23]~147_combout ),
	.datad(\myif.out[23]~146_combout ),
	.cin(gnd),
	.combout(\myif.out[23]~148_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~148 .lut_mask = 16'hF5A0;
defparam \myif.out[23]~148 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N2
cycloneive_lcell_comb \myif.out[23]~149 (
// Equation(s):
// \myif.out[23]~149_combout  = (\myif.out[13]~23_combout  & (((\myif.out[23]~148_combout )))) # (!\myif.out[13]~23_combout  & (\myif.out[23]~139_combout  & (\myif.out[23]~141_combout )))

	.dataa(\myif.out[13]~23_combout ),
	.datab(\myif.out[23]~139_combout ),
	.datac(\myif.out[23]~141_combout ),
	.datad(\myif.out[23]~148_combout ),
	.cin(gnd),
	.combout(\myif.out[23]~149_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[23]~149 .lut_mask = 16'hEA40;
defparam \myif.out[23]~149 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N16
cycloneive_lcell_comb \out~54 (
// Equation(s):
// \out~54_combout  = \rdat1[16]~19_combout  $ (((\port_b~21_combout ) # ((\port_b~0_combout  & fuifrtReplace_16))))

	.dataa(port_b),
	.datab(port_b11),
	.datac(rdat1_16),
	.datad(fuifrtReplace_16),
	.cin(gnd),
	.combout(\out~54_combout ),
	.cout());
// synopsys translate_off
defparam \out~54 .lut_mask = 16'h1E3C;
defparam \out~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N26
cycloneive_lcell_comb \out~53 (
// Equation(s):
// \out~53_combout  = (\rdat1[16]~19_combout  & ((\port_b~21_combout ) # ((\port_b~0_combout  & fuifrtReplace_16))))

	.dataa(port_b),
	.datab(fuifrtReplace_16),
	.datac(port_b11),
	.datad(rdat1_16),
	.cin(gnd),
	.combout(\out~53_combout ),
	.cout());
// synopsys translate_off
defparam \out~53 .lut_mask = 16'hF800;
defparam \out~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N24
cycloneive_lcell_comb \myif.out[16]~155 (
// Equation(s):
// \myif.out[16]~155_combout  = (\myif.out[13]~84_combout  & (((\out~53_combout ) # (!\myif.out[13]~83_combout )))) # (!\myif.out[13]~84_combout  & (\ShiftLeft0~102_combout  & ((\myif.out[13]~83_combout ))))

	.dataa(\ShiftLeft0~102_combout ),
	.datab(\myif.out[13]~84_combout ),
	.datac(\out~53_combout ),
	.datad(\myif.out[13]~83_combout ),
	.cin(gnd),
	.combout(\myif.out[16]~155_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[16]~155 .lut_mask = 16'hE2CC;
defparam \myif.out[16]~155 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N14
cycloneive_lcell_comb \myif.out[16]~156 (
// Equation(s):
// \myif.out[16]~156_combout  = (\myif.out[13]~82_combout  & (((\myif.out[16]~155_combout )))) # (!\myif.out[13]~82_combout  & ((\myif.out[16]~155_combout  & (\ShiftLeft0~39_combout )) # (!\myif.out[16]~155_combout  & ((\ShiftLeft0~30_combout )))))

	.dataa(\ShiftLeft0~39_combout ),
	.datab(\myif.out[13]~82_combout ),
	.datac(\ShiftLeft0~30_combout ),
	.datad(\myif.out[16]~155_combout ),
	.cin(gnd),
	.combout(\myif.out[16]~156_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[16]~156 .lut_mask = 16'hEE30;
defparam \myif.out[16]~156 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N28
cycloneive_lcell_comb \out~52 (
// Equation(s):
// \out~52_combout  = (\port_b~21_combout ) # ((\rdat1[16]~19_combout ) # ((\port_b~0_combout  & fuifrtReplace_16)))

	.dataa(port_b),
	.datab(fuifrtReplace_16),
	.datac(port_b11),
	.datad(rdat1_16),
	.cin(gnd),
	.combout(\out~52_combout ),
	.cout());
// synopsys translate_off
defparam \out~52 .lut_mask = 16'hFFF8;
defparam \out~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N6
cycloneive_lcell_comb \ShiftRight0~101 (
// Equation(s):
// \ShiftRight0~101_combout  = (\port_b~14_combout  & ((\port_b~10_combout  & ((\ShiftRight0~67_combout ))) # (!\port_b~10_combout  & (\ShiftRight0~62_combout ))))

	.dataa(port_b7),
	.datab(\ShiftRight0~62_combout ),
	.datac(port_b6),
	.datad(\ShiftRight0~67_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~101_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~101 .lut_mask = 16'hA808;
defparam \ShiftRight0~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N28
cycloneive_lcell_comb \ShiftRight0~102 (
// Equation(s):
// \ShiftRight0~102_combout  = (\ShiftRight0~101_combout ) # ((!\port_b~14_combout  & \ShiftRight0~93_combout ))

	.dataa(gnd),
	.datab(port_b7),
	.datac(\ShiftRight0~93_combout ),
	.datad(\ShiftRight0~101_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~102_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~102 .lut_mask = 16'hFF30;
defparam \ShiftRight0~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N18
cycloneive_lcell_comb \myif.out[16]~153 (
// Equation(s):
// \myif.out[16]~153_combout  = (idex_ifaluop_o_2 & ((\out~52_combout ) # ((!\myif.out[13]~23_combout )))) # (!idex_ifaluop_o_2 & (((\myif.out[13]~23_combout  & \ShiftRight0~102_combout ))))

	.dataa(\out~52_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\myif.out[13]~23_combout ),
	.datad(\ShiftRight0~102_combout ),
	.cin(gnd),
	.combout(\myif.out[16]~153_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[16]~153 .lut_mask = 16'hBC8C;
defparam \myif.out[16]~153 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N20
cycloneive_lcell_comb \myif.out[16]~154 (
// Equation(s):
// \myif.out[16]~154_combout  = (idex_ifaluop_o_1 & ((\myif.out[16]~153_combout  & ((!\out~52_combout ))) # (!\myif.out[16]~153_combout  & (\Add1~32_combout )))) # (!idex_ifaluop_o_1 & (((\myif.out[16]~153_combout ))))

	.dataa(\Add1~32_combout ),
	.datab(idex_ifaluop_o_1),
	.datac(\out~52_combout ),
	.datad(\myif.out[16]~153_combout ),
	.cin(gnd),
	.combout(\myif.out[16]~154_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[16]~154 .lut_mask = 16'h3F88;
defparam \myif.out[16]~154 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N0
cycloneive_lcell_comb \myif.out[16]~157 (
// Equation(s):
// \myif.out[16]~157_combout  = (\myif.out[23]~150_combout  & ((\myif.out[23]~135_combout ) # ((\myif.out[16]~154_combout )))) # (!\myif.out[23]~150_combout  & (!\myif.out[23]~135_combout  & (\myif.out[16]~156_combout )))

	.dataa(\myif.out[23]~150_combout ),
	.datab(\myif.out[23]~135_combout ),
	.datac(\myif.out[16]~156_combout ),
	.datad(\myif.out[16]~154_combout ),
	.cin(gnd),
	.combout(\myif.out[16]~157_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[16]~157 .lut_mask = 16'hBA98;
defparam \myif.out[16]~157 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N0
cycloneive_lcell_comb \out~55 (
// Equation(s):
// \out~55_combout  = (\rdat1[17]~63_combout  & ((\port_b~23_combout ) # ((\port_b~0_combout  & fuifrtReplace_17))))

	.dataa(port_b),
	.datab(port_b13),
	.datac(fuifrtReplace_17),
	.datad(rdat1_17),
	.cin(gnd),
	.combout(\out~55_combout ),
	.cout());
// synopsys translate_off
defparam \out~55 .lut_mask = 16'hEC00;
defparam \out~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N2
cycloneive_lcell_comb \myif.out[17]~159 (
// Equation(s):
// \myif.out[17]~159_combout  = (\myif.out[13]~84_combout  & (((\out~55_combout ) # (!\myif.out[13]~83_combout )))) # (!\myif.out[13]~84_combout  & (\ShiftLeft0~14_combout  & ((\myif.out[13]~83_combout ))))

	.dataa(\ShiftLeft0~14_combout ),
	.datab(\out~55_combout ),
	.datac(\myif.out[13]~84_combout ),
	.datad(\myif.out[13]~83_combout ),
	.cin(gnd),
	.combout(\myif.out[17]~159_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[17]~159 .lut_mask = 16'hCAF0;
defparam \myif.out[17]~159 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N12
cycloneive_lcell_comb \myif.out[17]~160 (
// Equation(s):
// \myif.out[17]~160_combout  = (\myif.out[13]~82_combout  & (((\myif.out[17]~159_combout )))) # (!\myif.out[13]~82_combout  & ((\myif.out[17]~159_combout  & ((\ShiftLeft0~72_combout ))) # (!\myif.out[17]~159_combout  & (\ShiftLeft0~61_combout ))))

	.dataa(\myif.out[13]~82_combout ),
	.datab(\ShiftLeft0~61_combout ),
	.datac(\ShiftLeft0~72_combout ),
	.datad(\myif.out[17]~159_combout ),
	.cin(gnd),
	.combout(\myif.out[17]~160_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[17]~160 .lut_mask = 16'hFA44;
defparam \myif.out[17]~160 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N16
cycloneive_lcell_comb \myif.out[17]~163 (
// Equation(s):
// \myif.out[17]~163_combout  = (idex_ifaluop_o_1 & (((\Add1~34_combout )))) # (!idex_ifaluop_o_1 & ((\myif.out[17]~161_combout ) # ((\rdat1[17]~63_combout ))))

	.dataa(\myif.out[17]~161_combout ),
	.datab(rdat1_17),
	.datac(idex_ifaluop_o_1),
	.datad(\Add1~34_combout ),
	.cin(gnd),
	.combout(\myif.out[17]~163_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[17]~163 .lut_mask = 16'hFE0E;
defparam \myif.out[17]~163 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N18
cycloneive_lcell_comb \myif.out[17]~164 (
// Equation(s):
// \myif.out[17]~164_combout  = (\myif.out[23]~135_combout  & (((\Add0~34_combout )))) # (!\myif.out[23]~135_combout  & ((idex_ifaluop_o_2) # ((\myif.out[17]~163_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\myif.out[23]~135_combout ),
	.datac(\Add0~34_combout ),
	.datad(\myif.out[17]~163_combout ),
	.cin(gnd),
	.combout(\myif.out[17]~164_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[17]~164 .lut_mask = 16'hF3E2;
defparam \myif.out[17]~164 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N4
cycloneive_lcell_comb \myif.out[17]~161 (
// Equation(s):
// \myif.out[17]~161_combout  = \rdat1[17]~63_combout  $ (((\port_b~23_combout ) # ((\port_b~0_combout  & fuifrtReplace_17))))

	.dataa(rdat1_17),
	.datab(port_b),
	.datac(port_b13),
	.datad(fuifrtReplace_17),
	.cin(gnd),
	.combout(\myif.out[17]~161_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[17]~161 .lut_mask = 16'h565A;
defparam \myif.out[17]~161 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N26
cycloneive_lcell_comb \myif.out[17]~162 (
// Equation(s):
// \myif.out[17]~162_combout  = (idex_ifaluop_o_1 & (((!\rdat1[17]~63_combout  & !\myif.out[17]~161_combout )) # (!idex_ifaluop_o_2))) # (!idex_ifaluop_o_1 & (((idex_ifaluop_o_2))))

	.dataa(rdat1_17),
	.datab(idex_ifaluop_o_1),
	.datac(idex_ifaluop_o_2),
	.datad(\myif.out[17]~161_combout ),
	.cin(gnd),
	.combout(\myif.out[17]~162_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[17]~162 .lut_mask = 16'h3C7C;
defparam \myif.out[17]~162 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N8
cycloneive_lcell_comb \myif.out[17]~165 (
// Equation(s):
// \myif.out[17]~165_combout  = (\port_b~23_combout ) # ((\port_b~0_combout  & fuifrtReplace_17))

	.dataa(port_b),
	.datab(gnd),
	.datac(fuifrtReplace_17),
	.datad(port_b13),
	.cin(gnd),
	.combout(\myif.out[17]~165_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[17]~165 .lut_mask = 16'hFFA0;
defparam \myif.out[17]~165 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N14
cycloneive_lcell_comb \myif.out[17]~170 (
// Equation(s):
// \myif.out[17]~170_combout  = (\rdat1[17]~63_combout  & (!idex_ifaluop_o_1)) # (!\rdat1[17]~63_combout  & ((idex_ifaluop_o_1 & (!\myif.out[17]~165_combout  & \Add1~34_combout )) # (!idex_ifaluop_o_1 & (\myif.out[17]~165_combout ))))

	.dataa(rdat1_17),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[17]~165_combout ),
	.datad(\Add1~34_combout ),
	.cin(gnd),
	.combout(\myif.out[17]~170_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[17]~170 .lut_mask = 16'h3632;
defparam \myif.out[17]~170 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N4
cycloneive_lcell_comb \myif.out[17]~167 (
// Equation(s):
// \myif.out[17]~167_combout  = (\port_b~23_combout ) # ((\rdat1[17]~63_combout ) # ((\port_b~0_combout  & fuifrtReplace_17)))

	.dataa(port_b),
	.datab(port_b13),
	.datac(fuifrtReplace_17),
	.datad(rdat1_17),
	.cin(gnd),
	.combout(\myif.out[17]~167_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[17]~167 .lut_mask = 16'hFFEC;
defparam \myif.out[17]~167 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N6
cycloneive_lcell_comb \myif.out[17]~168 (
// Equation(s):
// \myif.out[17]~168_combout  = (idex_ifaluop_o_1 & (\Add1~34_combout  & ((!\myif.out[17]~167_combout ) # (!idex_ifaluop_o_2)))) # (!idex_ifaluop_o_1 & (idex_ifaluop_o_2 & (\myif.out[17]~167_combout )))

	.dataa(idex_ifaluop_o_2),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[17]~167_combout ),
	.datad(\Add1~34_combout ),
	.cin(gnd),
	.combout(\myif.out[17]~168_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[17]~168 .lut_mask = 16'h6C20;
defparam \myif.out[17]~168 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N28
cycloneive_lcell_comb \myif.out[17]~169 (
// Equation(s):
// \myif.out[17]~169_combout  = (\ShiftRight0~30_combout  & (\myif.out[17]~166_combout )) # (!\ShiftRight0~30_combout  & ((\myif.out[17]~168_combout )))

	.dataa(\myif.out[17]~166_combout ),
	.datab(gnd),
	.datac(\ShiftRight0~30_combout ),
	.datad(\myif.out[17]~168_combout ),
	.cin(gnd),
	.combout(\myif.out[17]~169_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[17]~169 .lut_mask = 16'hAFA0;
defparam \myif.out[17]~169 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N24
cycloneive_lcell_comb \myif.out[17]~171 (
// Equation(s):
// \myif.out[17]~171_combout  = (idex_ifaluop_o_2 & (\myif.out[17]~170_combout )) # (!idex_ifaluop_o_2 & ((\myif.out[17]~169_combout )))

	.dataa(gnd),
	.datab(idex_ifaluop_o_2),
	.datac(\myif.out[17]~170_combout ),
	.datad(\myif.out[17]~169_combout ),
	.cin(gnd),
	.combout(\myif.out[17]~171_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[17]~171 .lut_mask = 16'hF3C0;
defparam \myif.out[17]~171 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N30
cycloneive_lcell_comb \myif.out[17]~172 (
// Equation(s):
// \myif.out[17]~172_combout  = (\myif.out[13]~23_combout  & (((\myif.out[17]~171_combout )))) # (!\myif.out[13]~23_combout  & (\myif.out[17]~164_combout  & (\myif.out[17]~162_combout )))

	.dataa(\myif.out[13]~23_combout ),
	.datab(\myif.out[17]~164_combout ),
	.datac(\myif.out[17]~162_combout ),
	.datad(\myif.out[17]~171_combout ),
	.cin(gnd),
	.combout(\myif.out[17]~172_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[17]~172 .lut_mask = 16'hEA40;
defparam \myif.out[17]~172 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N20
cycloneive_lcell_comb \myif.out[17]~173 (
// Equation(s):
// \myif.out[17]~173_combout  = (\myif.out[23]~150_combout  & ((\myif.out[17]~161_combout ) # ((!\myif.out[23]~135_combout )))) # (!\myif.out[23]~150_combout  & (((\myif.out[23]~135_combout  & \myif.out[17]~164_combout ))))

	.dataa(\myif.out[17]~161_combout ),
	.datab(\myif.out[23]~150_combout ),
	.datac(\myif.out[23]~135_combout ),
	.datad(\myif.out[17]~164_combout ),
	.cin(gnd),
	.combout(\myif.out[17]~173_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[17]~173 .lut_mask = 16'hBC8C;
defparam \myif.out[17]~173 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N2
cycloneive_lcell_comb \out~58 (
// Equation(s):
// \out~58_combout  = \rdat1[18]~59_combout  $ (((\port_b~25_combout ) # ((\port_b~0_combout  & fuifrtReplace_18))))

	.dataa(rdat1_18),
	.datab(port_b),
	.datac(fuifrtReplace_18),
	.datad(port_b15),
	.cin(gnd),
	.combout(\out~58_combout ),
	.cout());
// synopsys translate_off
defparam \out~58 .lut_mask = 16'h556A;
defparam \out~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N18
cycloneive_lcell_comb \out~56 (
// Equation(s):
// \out~56_combout  = (\port_b~25_combout ) # ((\rdat1[18]~59_combout ) # ((fuifrtReplace_18 & \port_b~0_combout )))

	.dataa(port_b15),
	.datab(fuifrtReplace_18),
	.datac(rdat1_18),
	.datad(port_b),
	.cin(gnd),
	.combout(\out~56_combout ),
	.cout());
// synopsys translate_off
defparam \out~56 .lut_mask = 16'hFEFA;
defparam \out~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N24
cycloneive_lcell_comb \ShiftRight0~103 (
// Equation(s):
// \ShiftRight0~103_combout  = (\port_b~14_combout  & (\ShiftRight0~70_combout )) # (!\port_b~14_combout  & ((\ShiftRight0~98_combout )))

	.dataa(gnd),
	.datab(port_b7),
	.datac(\ShiftRight0~70_combout ),
	.datad(\ShiftRight0~98_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~103_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~103 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N22
cycloneive_lcell_comb \myif.out[18]~175 (
// Equation(s):
// \myif.out[18]~175_combout  = (idex_ifaluop_o_2 & ((\out~56_combout ) # ((!\myif.out[13]~23_combout )))) # (!idex_ifaluop_o_2 & (((\myif.out[13]~23_combout  & \ShiftRight0~103_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\out~56_combout ),
	.datac(\myif.out[13]~23_combout ),
	.datad(\ShiftRight0~103_combout ),
	.cin(gnd),
	.combout(\myif.out[18]~175_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[18]~175 .lut_mask = 16'hDA8A;
defparam \myif.out[18]~175 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N8
cycloneive_lcell_comb \myif.out[18]~176 (
// Equation(s):
// \myif.out[18]~176_combout  = (idex_ifaluop_o_1 & ((\myif.out[18]~175_combout  & (!\out~56_combout )) # (!\myif.out[18]~175_combout  & ((\Add1~36_combout ))))) # (!idex_ifaluop_o_1 & (((\myif.out[18]~175_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(\out~56_combout ),
	.datac(\myif.out[18]~175_combout ),
	.datad(\Add1~36_combout ),
	.cin(gnd),
	.combout(\myif.out[18]~176_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[18]~176 .lut_mask = 16'h7A70;
defparam \myif.out[18]~176 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N4
cycloneive_lcell_comb \ShiftLeft0~103 (
// Equation(s):
// \ShiftLeft0~103_combout  = (!\port_b~14_combout  & (!\port_b~10_combout  & \ShiftLeft0~16_combout ))

	.dataa(port_b7),
	.datab(gnd),
	.datac(port_b6),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~103_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~103 .lut_mask = 16'h0500;
defparam \ShiftLeft0~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N16
cycloneive_lcell_comb \myif.out[18]~177 (
// Equation(s):
// \myif.out[18]~177_combout  = (\myif.out[13]~84_combout  & ((\out~57_combout ) # ((!\myif.out[13]~83_combout )))) # (!\myif.out[13]~84_combout  & (((\ShiftLeft0~103_combout  & \myif.out[13]~83_combout ))))

	.dataa(\out~57_combout ),
	.datab(\ShiftLeft0~103_combout ),
	.datac(\myif.out[13]~84_combout ),
	.datad(\myif.out[13]~83_combout ),
	.cin(gnd),
	.combout(\myif.out[18]~177_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[18]~177 .lut_mask = 16'hACF0;
defparam \myif.out[18]~177 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N10
cycloneive_lcell_comb \myif.out[18]~178 (
// Equation(s):
// \myif.out[18]~178_combout  = (\myif.out[13]~82_combout  & (((\myif.out[18]~177_combout )))) # (!\myif.out[13]~82_combout  & ((\myif.out[18]~177_combout  & (\ShiftLeft0~53_combout )) # (!\myif.out[18]~177_combout  & ((\ShiftLeft0~48_combout )))))

	.dataa(\ShiftLeft0~53_combout ),
	.datab(\ShiftLeft0~48_combout ),
	.datac(\myif.out[13]~82_combout ),
	.datad(\myif.out[18]~177_combout ),
	.cin(gnd),
	.combout(\myif.out[18]~178_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[18]~178 .lut_mask = 16'hFA0C;
defparam \myif.out[18]~178 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N0
cycloneive_lcell_comb \myif.out[18]~179 (
// Equation(s):
// \myif.out[18]~179_combout  = (\myif.out[23]~135_combout  & (\myif.out[23]~150_combout )) # (!\myif.out[23]~135_combout  & ((\myif.out[23]~150_combout  & (\myif.out[18]~176_combout )) # (!\myif.out[23]~150_combout  & ((\myif.out[18]~178_combout )))))

	.dataa(\myif.out[23]~135_combout ),
	.datab(\myif.out[23]~150_combout ),
	.datac(\myif.out[18]~176_combout ),
	.datad(\myif.out[18]~178_combout ),
	.cin(gnd),
	.combout(\myif.out[18]~179_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[18]~179 .lut_mask = 16'hD9C8;
defparam \myif.out[18]~179 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N30
cycloneive_lcell_comb \myif.out[19]~183 (
// Equation(s):
// \myif.out[19]~183_combout  = \rdat1[19]~61_combout  $ (((\port_b~27_combout ) # ((\port_b~0_combout  & fuifrtReplace_19))))

	.dataa(port_b17),
	.datab(rdat1_19),
	.datac(port_b),
	.datad(fuifrtReplace_19),
	.cin(gnd),
	.combout(\myif.out[19]~183_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[19]~183 .lut_mask = 16'h3666;
defparam \myif.out[19]~183 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N6
cycloneive_lcell_comb \myif.out[19]~185 (
// Equation(s):
// \myif.out[19]~185_combout  = (idex_ifaluop_o_1 & (((\Add1~38_combout )))) # (!idex_ifaluop_o_1 & ((\rdat1[19]~61_combout ) # ((\myif.out[19]~183_combout ))))

	.dataa(rdat1_19),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[19]~183_combout ),
	.datad(\Add1~38_combout ),
	.cin(gnd),
	.combout(\myif.out[19]~185_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[19]~185 .lut_mask = 16'hFE32;
defparam \myif.out[19]~185 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N0
cycloneive_lcell_comb \myif.out[19]~186 (
// Equation(s):
// \myif.out[19]~186_combout  = (\myif.out[23]~135_combout  & (((\Add0~38_combout )))) # (!\myif.out[23]~135_combout  & ((idex_ifaluop_o_2) # ((\myif.out[19]~185_combout ))))

	.dataa(\myif.out[23]~135_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\Add0~38_combout ),
	.datad(\myif.out[19]~185_combout ),
	.cin(gnd),
	.combout(\myif.out[19]~186_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[19]~186 .lut_mask = 16'hF5E4;
defparam \myif.out[19]~186 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N24
cycloneive_lcell_comb \myif.out[19]~195 (
// Equation(s):
// \myif.out[19]~195_combout  = (\myif.out[23]~135_combout  & ((\myif.out[23]~150_combout  & (\myif.out[19]~183_combout )) # (!\myif.out[23]~150_combout  & ((\myif.out[19]~186_combout ))))) # (!\myif.out[23]~135_combout  & (!\myif.out[23]~150_combout ))

	.dataa(\myif.out[23]~135_combout ),
	.datab(\myif.out[23]~150_combout ),
	.datac(\myif.out[19]~183_combout ),
	.datad(\myif.out[19]~186_combout ),
	.cin(gnd),
	.combout(\myif.out[19]~195_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[19]~195 .lut_mask = 16'hB391;
defparam \myif.out[19]~195 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N14
cycloneive_lcell_comb \out~59 (
// Equation(s):
// \out~59_combout  = (\rdat1[19]~61_combout  & ((\port_b~27_combout ) # ((\port_b~0_combout  & fuifrtReplace_19))))

	.dataa(port_b),
	.datab(port_b17),
	.datac(fuifrtReplace_19),
	.datad(rdat1_19),
	.cin(gnd),
	.combout(\out~59_combout ),
	.cout());
// synopsys translate_off
defparam \out~59 .lut_mask = 16'hEC00;
defparam \out~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N0
cycloneive_lcell_comb \myif.out[19]~181 (
// Equation(s):
// \myif.out[19]~181_combout  = (\myif.out[13]~84_combout  & (((\out~59_combout ) # (!\myif.out[13]~83_combout )))) # (!\myif.out[13]~84_combout  & (\ShiftLeft0~109_combout  & ((\myif.out[13]~83_combout ))))

	.dataa(\ShiftLeft0~109_combout ),
	.datab(\myif.out[13]~84_combout ),
	.datac(\out~59_combout ),
	.datad(\myif.out[13]~83_combout ),
	.cin(gnd),
	.combout(\myif.out[19]~181_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[19]~181 .lut_mask = 16'hE2CC;
defparam \myif.out[19]~181 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N26
cycloneive_lcell_comb \myif.out[19]~182 (
// Equation(s):
// \myif.out[19]~182_combout  = (\myif.out[13]~82_combout  & (((\myif.out[19]~181_combout )))) # (!\myif.out[13]~82_combout  & ((\myif.out[19]~181_combout  & (\ShiftLeft0~84_combout )) # (!\myif.out[19]~181_combout  & ((\ShiftLeft0~78_combout )))))

	.dataa(\ShiftLeft0~84_combout ),
	.datab(\myif.out[13]~82_combout ),
	.datac(\ShiftLeft0~78_combout ),
	.datad(\myif.out[19]~181_combout ),
	.cin(gnd),
	.combout(\myif.out[19]~182_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[19]~182 .lut_mask = 16'hEE30;
defparam \myif.out[19]~182 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N16
cycloneive_lcell_comb \myif.out[19]~184 (
// Equation(s):
// \myif.out[19]~184_combout  = (idex_ifaluop_o_2 & (((!\myif.out[19]~183_combout  & !\rdat1[19]~61_combout )) # (!idex_ifaluop_o_1))) # (!idex_ifaluop_o_2 & (idex_ifaluop_o_1))

	.dataa(idex_ifaluop_o_2),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[19]~183_combout ),
	.datad(rdat1_19),
	.cin(gnd),
	.combout(\myif.out[19]~184_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[19]~184 .lut_mask = 16'h666E;
defparam \myif.out[19]~184 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N4
cycloneive_lcell_comb \myif.out[19]~187 (
// Equation(s):
// \myif.out[19]~187_combout  = (\port_b~27_combout ) # ((\port_b~0_combout  & fuifrtReplace_19))

	.dataa(port_b17),
	.datab(port_b),
	.datac(gnd),
	.datad(fuifrtReplace_19),
	.cin(gnd),
	.combout(\myif.out[19]~187_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[19]~187 .lut_mask = 16'hEEAA;
defparam \myif.out[19]~187 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N14
cycloneive_lcell_comb \myif.out[19]~192 (
// Equation(s):
// \myif.out[19]~192_combout  = (\rdat1[19]~61_combout  & (!idex_ifaluop_o_1)) # (!\rdat1[19]~61_combout  & ((idex_ifaluop_o_1 & (!\myif.out[19]~187_combout  & \Add1~38_combout )) # (!idex_ifaluop_o_1 & (\myif.out[19]~187_combout ))))

	.dataa(rdat1_19),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[19]~187_combout ),
	.datad(\Add1~38_combout ),
	.cin(gnd),
	.combout(\myif.out[19]~192_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[19]~192 .lut_mask = 16'h3632;
defparam \myif.out[19]~192 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N28
cycloneive_lcell_comb \ShiftRight0~104 (
// Equation(s):
// \ShiftRight0~104_combout  = (\port_b~10_combout  & (\ShiftRight0~73_combout )) # (!\port_b~10_combout  & ((\ShiftRight0~75_combout )))

	.dataa(\ShiftRight0~73_combout ),
	.datab(port_b6),
	.datac(gnd),
	.datad(\ShiftRight0~75_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~104_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~104 .lut_mask = 16'hBB88;
defparam \ShiftRight0~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N6
cycloneive_lcell_comb \ShiftRight0~105 (
// Equation(s):
// \ShiftRight0~105_combout  = (\port_b~14_combout  & (\ShiftRight0~104_combout )) # (!\port_b~14_combout  & ((\ShiftRight0~100_combout )))

	.dataa(port_b7),
	.datab(\ShiftRight0~104_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~100_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~105_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~105 .lut_mask = 16'hDD88;
defparam \ShiftRight0~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N24
cycloneive_lcell_comb \myif.out[19]~189 (
// Equation(s):
// \myif.out[19]~189_combout  = (\port_b~27_combout ) # ((\rdat1[19]~61_combout ) # ((\port_b~0_combout  & fuifrtReplace_19)))

	.dataa(port_b17),
	.datab(rdat1_19),
	.datac(port_b),
	.datad(fuifrtReplace_19),
	.cin(gnd),
	.combout(\myif.out[19]~189_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[19]~189 .lut_mask = 16'hFEEE;
defparam \myif.out[19]~189 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N12
cycloneive_lcell_comb \myif.out[19]~190 (
// Equation(s):
// \myif.out[19]~190_combout  = (idex_ifaluop_o_1 & (\Add1~38_combout  & ((!\myif.out[19]~189_combout ) # (!idex_ifaluop_o_2)))) # (!idex_ifaluop_o_1 & (idex_ifaluop_o_2 & (\myif.out[19]~189_combout )))

	.dataa(idex_ifaluop_o_2),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[19]~189_combout ),
	.datad(\Add1~38_combout ),
	.cin(gnd),
	.combout(\myif.out[19]~190_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[19]~190 .lut_mask = 16'h6C20;
defparam \myif.out[19]~190 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N20
cycloneive_lcell_comb \myif.out[19]~191 (
// Equation(s):
// \myif.out[19]~191_combout  = (\ShiftRight0~105_combout  & (\myif.out[19]~188_combout )) # (!\ShiftRight0~105_combout  & ((\myif.out[19]~190_combout )))

	.dataa(\myif.out[19]~188_combout ),
	.datab(\ShiftRight0~105_combout ),
	.datac(gnd),
	.datad(\myif.out[19]~190_combout ),
	.cin(gnd),
	.combout(\myif.out[19]~191_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[19]~191 .lut_mask = 16'hBB88;
defparam \myif.out[19]~191 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N4
cycloneive_lcell_comb \myif.out[19]~193 (
// Equation(s):
// \myif.out[19]~193_combout  = (idex_ifaluop_o_2 & (\myif.out[19]~192_combout )) # (!idex_ifaluop_o_2 & ((\myif.out[19]~191_combout )))

	.dataa(idex_ifaluop_o_2),
	.datab(gnd),
	.datac(\myif.out[19]~192_combout ),
	.datad(\myif.out[19]~191_combout ),
	.cin(gnd),
	.combout(\myif.out[19]~193_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[19]~193 .lut_mask = 16'hF5A0;
defparam \myif.out[19]~193 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N18
cycloneive_lcell_comb \myif.out[19]~194 (
// Equation(s):
// \myif.out[19]~194_combout  = (\myif.out[13]~23_combout  & (((\myif.out[19]~193_combout )))) # (!\myif.out[13]~23_combout  & (\myif.out[19]~184_combout  & ((\myif.out[19]~186_combout ))))

	.dataa(\myif.out[19]~184_combout ),
	.datab(\myif.out[13]~23_combout ),
	.datac(\myif.out[19]~193_combout ),
	.datad(\myif.out[19]~186_combout ),
	.cin(gnd),
	.combout(\myif.out[19]~194_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[19]~194 .lut_mask = 16'hE2C0;
defparam \myif.out[19]~194 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N12
cycloneive_lcell_comb \out~62 (
// Equation(s):
// \out~62_combout  = \rdat1[30]~39_combout  $ (((\port_b~57_combout ) # ((fuifrtReplace_30 & \port_b~0_combout ))))

	.dataa(fuifrtReplace_30),
	.datab(port_b),
	.datac(port_b47),
	.datad(rdat1_30),
	.cin(gnd),
	.combout(\out~62_combout ),
	.cout());
// synopsys translate_off
defparam \out~62 .lut_mask = 16'h07F8;
defparam \out~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N24
cycloneive_lcell_comb \Add0~56 (
// Equation(s):
// \Add0~56_combout  = ((\rdat1[28]~41_combout  $ (\port_b~54_combout  $ (!\Add0~55 )))) # (GND)
// \Add0~57  = CARRY((\rdat1[28]~41_combout  & ((\port_b~54_combout ) # (!\Add0~55 ))) # (!\rdat1[28]~41_combout  & (\port_b~54_combout  & !\Add0~55 )))

	.dataa(rdat1_28),
	.datab(port_b44),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~55 ),
	.combout(\Add0~56_combout ),
	.cout(\Add0~57 ));
// synopsys translate_off
defparam \Add0~56 .lut_mask = 16'h698E;
defparam \Add0~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N26
cycloneive_lcell_comb \Add0~58 (
// Equation(s):
// \Add0~58_combout  = (\port_b~56_combout  & ((\rdat1[29]~37_combout  & (\Add0~57  & VCC)) # (!\rdat1[29]~37_combout  & (!\Add0~57 )))) # (!\port_b~56_combout  & ((\rdat1[29]~37_combout  & (!\Add0~57 )) # (!\rdat1[29]~37_combout  & ((\Add0~57 ) # (GND)))))
// \Add0~59  = CARRY((\port_b~56_combout  & (!\rdat1[29]~37_combout  & !\Add0~57 )) # (!\port_b~56_combout  & ((!\Add0~57 ) # (!\rdat1[29]~37_combout ))))

	.dataa(port_b46),
	.datab(rdat1_29),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~57 ),
	.combout(\Add0~58_combout ),
	.cout(\Add0~59 ));
// synopsys translate_off
defparam \Add0~58 .lut_mask = 16'h9617;
defparam \Add0~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N28
cycloneive_lcell_comb \Add0~60 (
// Equation(s):
// \Add0~60_combout  = ((\rdat1[30]~39_combout  $ (\port_b~58_combout  $ (!\Add0~59 )))) # (GND)
// \Add0~61  = CARRY((\rdat1[30]~39_combout  & ((\port_b~58_combout ) # (!\Add0~59 ))) # (!\rdat1[30]~39_combout  & (\port_b~58_combout  & !\Add0~59 )))

	.dataa(rdat1_30),
	.datab(port_b48),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~59 ),
	.combout(\Add0~60_combout ),
	.cout(\Add0~61 ));
// synopsys translate_off
defparam \Add0~60 .lut_mask = 16'h698E;
defparam \Add0~60 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N10
cycloneive_lcell_comb \ShiftLeft0~41 (
// Equation(s):
// \ShiftLeft0~41_combout  = (\port_b~4_combout  & ((\rdat1[19]~61_combout ))) # (!\port_b~4_combout  & (\rdat1[21]~55_combout ))

	.dataa(gnd),
	.datab(rdat1_21),
	.datac(port_b2),
	.datad(rdat1_19),
	.cin(gnd),
	.combout(\ShiftLeft0~41_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~41 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N24
cycloneive_lcell_comb \ShiftLeft0~43 (
// Equation(s):
// \ShiftLeft0~43_combout  = (\port_b~7_combout  & (\ShiftLeft0~41_combout )) # (!\port_b~7_combout  & ((\ShiftLeft0~42_combout )))

	.dataa(gnd),
	.datab(port_b4),
	.datac(\ShiftLeft0~41_combout ),
	.datad(\ShiftLeft0~42_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~43_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~43 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N26
cycloneive_lcell_comb \ShiftLeft0~105 (
// Equation(s):
// \ShiftLeft0~105_combout  = (\port_b~10_combout  & ((\ShiftLeft0~46_combout ) # ((\ShiftLeft0~47_combout )))) # (!\port_b~10_combout  & (((\ShiftLeft0~43_combout ))))

	.dataa(\ShiftLeft0~46_combout ),
	.datab(\ShiftLeft0~47_combout ),
	.datac(port_b6),
	.datad(\ShiftLeft0~43_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~105_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~105 .lut_mask = 16'hEFE0;
defparam \ShiftLeft0~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N0
cycloneive_lcell_comb \myif.negative~0 (
// Equation(s):
// \myif.negative~0_combout  = (\port_b~10_combout ) # ((!\port_b~4_combout  & \port_b~7_combout ))

	.dataa(port_b2),
	.datab(port_b4),
	.datac(gnd),
	.datad(port_b6),
	.cin(gnd),
	.combout(\myif.negative~0_combout ),
	.cout());
// synopsys translate_off
defparam \myif.negative~0 .lut_mask = 16'hFF44;
defparam \myif.negative~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N4
cycloneive_lcell_comb \ShiftLeft0~50 (
// Equation(s):
// \ShiftLeft0~50_combout  = (\port_b~7_combout  & (\rdat1[25]~47_combout )) # (!\port_b~7_combout  & ((\rdat1[26]~43_combout )))

	.dataa(gnd),
	.datab(port_b4),
	.datac(rdat1_25),
	.datad(rdat1_26),
	.cin(gnd),
	.combout(\ShiftLeft0~50_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~50 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N14
cycloneive_lcell_comb \ShiftLeft0~49 (
// Equation(s):
// \ShiftLeft0~49_combout  = (\port_b~4_combout  & ((\port_b~7_combout  & ((\rdat1[23]~53_combout ))) # (!\port_b~7_combout  & (\rdat1[24]~49_combout ))))

	.dataa(rdat1_24),
	.datab(port_b4),
	.datac(rdat1_23),
	.datad(port_b2),
	.cin(gnd),
	.combout(\ShiftLeft0~49_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~49 .lut_mask = 16'hE200;
defparam \ShiftLeft0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N30
cycloneive_lcell_comb \ShiftLeft0~51 (
// Equation(s):
// \ShiftLeft0~51_combout  = (\ShiftLeft0~49_combout ) # ((!\port_b~4_combout  & \ShiftLeft0~50_combout ))

	.dataa(gnd),
	.datab(port_b2),
	.datac(\ShiftLeft0~50_combout ),
	.datad(\ShiftLeft0~49_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~51_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~51 .lut_mask = 16'hFF30;
defparam \ShiftLeft0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N18
cycloneive_lcell_comb \ShiftLeft0~104 (
// Equation(s):
// \ShiftLeft0~104_combout  = (\port_b~7_combout  & ((\rdat1[27]~45_combout ))) # (!\port_b~7_combout  & (\rdat1[28]~41_combout ))

	.dataa(rdat1_28),
	.datab(port_b4),
	.datac(gnd),
	.datad(rdat1_27),
	.cin(gnd),
	.combout(\ShiftLeft0~104_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~104 .lut_mask = 16'hEE22;
defparam \ShiftLeft0~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N4
cycloneive_lcell_comb \myif.out[30]~199 (
// Equation(s):
// \myif.out[30]~199_combout  = (\ShiftLeft0~13_combout  & (((\ShiftLeft0~104_combout ) # (\myif.negative~0_combout )))) # (!\ShiftLeft0~13_combout  & (\rdat1[30]~39_combout  & ((!\myif.negative~0_combout ))))

	.dataa(\ShiftLeft0~13_combout ),
	.datab(rdat1_30),
	.datac(\ShiftLeft0~104_combout ),
	.datad(\myif.negative~0_combout ),
	.cin(gnd),
	.combout(\myif.out[30]~199_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[30]~199 .lut_mask = 16'hAAE4;
defparam \myif.out[30]~199 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N18
cycloneive_lcell_comb \myif.out[30]~200 (
// Equation(s):
// \myif.out[30]~200_combout  = (\myif.negative~0_combout  & ((\myif.out[30]~199_combout  & ((\ShiftLeft0~51_combout ))) # (!\myif.out[30]~199_combout  & (\rdat1[29]~37_combout )))) # (!\myif.negative~0_combout  & (((\myif.out[30]~199_combout ))))

	.dataa(rdat1_29),
	.datab(\myif.negative~0_combout ),
	.datac(\ShiftLeft0~51_combout ),
	.datad(\myif.out[30]~199_combout ),
	.cin(gnd),
	.combout(\myif.out[30]~200_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[30]~200 .lut_mask = 16'hF388;
defparam \myif.out[30]~200 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N20
cycloneive_lcell_comb \myif.out[30]~201 (
// Equation(s):
// \myif.out[30]~201_combout  = (\myif.out[13]~84_combout  & ((\out~61_combout ) # ((!\myif.out[13]~83_combout )))) # (!\myif.out[13]~84_combout  & (((\myif.out[13]~83_combout  & \ShiftLeft0~94_combout ))))

	.dataa(\out~61_combout ),
	.datab(\myif.out[13]~84_combout ),
	.datac(\myif.out[13]~83_combout ),
	.datad(\ShiftLeft0~94_combout ),
	.cin(gnd),
	.combout(\myif.out[30]~201_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[30]~201 .lut_mask = 16'hBC8C;
defparam \myif.out[30]~201 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N22
cycloneive_lcell_comb \myif.out[30]~202 (
// Equation(s):
// \myif.out[30]~202_combout  = (\myif.out[13]~82_combout  & (((\myif.out[30]~201_combout )))) # (!\myif.out[13]~82_combout  & ((\myif.out[30]~201_combout  & (\ShiftLeft0~105_combout )) # (!\myif.out[30]~201_combout  & ((\myif.out[30]~200_combout )))))

	.dataa(\myif.out[13]~82_combout ),
	.datab(\ShiftLeft0~105_combout ),
	.datac(\myif.out[30]~200_combout ),
	.datad(\myif.out[30]~201_combout ),
	.cin(gnd),
	.combout(\myif.out[30]~202_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[30]~202 .lut_mask = 16'hEE50;
defparam \myif.out[30]~202 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N24
cycloneive_lcell_comb \Add1~56 (
// Equation(s):
// \Add1~56_combout  = ((\port_b~54_combout  $ (\rdat1[28]~41_combout  $ (\Add1~55 )))) # (GND)
// \Add1~57  = CARRY((\port_b~54_combout  & (\rdat1[28]~41_combout  & !\Add1~55 )) # (!\port_b~54_combout  & ((\rdat1[28]~41_combout ) # (!\Add1~55 ))))

	.dataa(port_b44),
	.datab(rdat1_28),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~55 ),
	.combout(\Add1~56_combout ),
	.cout(\Add1~57 ));
// synopsys translate_off
defparam \Add1~56 .lut_mask = 16'h964D;
defparam \Add1~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N26
cycloneive_lcell_comb \Add1~58 (
// Equation(s):
// \Add1~58_combout  = (\port_b~56_combout  & ((\rdat1[29]~37_combout  & (!\Add1~57 )) # (!\rdat1[29]~37_combout  & ((\Add1~57 ) # (GND))))) # (!\port_b~56_combout  & ((\rdat1[29]~37_combout  & (\Add1~57  & VCC)) # (!\rdat1[29]~37_combout  & (!\Add1~57 ))))
// \Add1~59  = CARRY((\port_b~56_combout  & ((!\Add1~57 ) # (!\rdat1[29]~37_combout ))) # (!\port_b~56_combout  & (!\rdat1[29]~37_combout  & !\Add1~57 )))

	.dataa(port_b46),
	.datab(rdat1_29),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~57 ),
	.combout(\Add1~58_combout ),
	.cout(\Add1~59 ));
// synopsys translate_off
defparam \Add1~58 .lut_mask = 16'h692B;
defparam \Add1~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N28
cycloneive_lcell_comb \Add1~60 (
// Equation(s):
// \Add1~60_combout  = ((\port_b~58_combout  $ (\rdat1[30]~39_combout  $ (\Add1~59 )))) # (GND)
// \Add1~61  = CARRY((\port_b~58_combout  & (\rdat1[30]~39_combout  & !\Add1~59 )) # (!\port_b~58_combout  & ((\rdat1[30]~39_combout ) # (!\Add1~59 ))))

	.dataa(port_b48),
	.datab(rdat1_30),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~59 ),
	.combout(\Add1~60_combout ),
	.cout(\Add1~61 ));
// synopsys translate_off
defparam \Add1~60 .lut_mask = 16'h964D;
defparam \Add1~60 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N20
cycloneive_lcell_comb \out~60 (
// Equation(s):
// \out~60_combout  = (\rdat1[30]~39_combout ) # ((\port_b~57_combout ) # ((\port_b~0_combout  & fuifrtReplace_30)))

	.dataa(port_b),
	.datab(rdat1_30),
	.datac(port_b47),
	.datad(fuifrtReplace_30),
	.cin(gnd),
	.combout(\out~60_combout ),
	.cout());
// synopsys translate_off
defparam \out~60 .lut_mask = 16'hFEFC;
defparam \out~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N18
cycloneive_lcell_comb \myif.out[30]~198 (
// Equation(s):
// \myif.out[30]~198_combout  = (\myif.out[30]~197_combout  & (((!\out~60_combout )) # (!idex_ifaluop_o_1))) # (!\myif.out[30]~197_combout  & (idex_ifaluop_o_1 & (\Add1~60_combout )))

	.dataa(\myif.out[30]~197_combout ),
	.datab(idex_ifaluop_o_1),
	.datac(\Add1~60_combout ),
	.datad(\out~60_combout ),
	.cin(gnd),
	.combout(\myif.out[30]~198_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[30]~198 .lut_mask = 16'h62EA;
defparam \myif.out[30]~198 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N0
cycloneive_lcell_comb \myif.out[30]~203 (
// Equation(s):
// \myif.out[30]~203_combout  = (\myif.out[23]~150_combout  & ((\myif.out[23]~135_combout ) # ((\myif.out[30]~198_combout )))) # (!\myif.out[23]~150_combout  & (!\myif.out[23]~135_combout  & (\myif.out[30]~202_combout )))

	.dataa(\myif.out[23]~150_combout ),
	.datab(\myif.out[23]~135_combout ),
	.datac(\myif.out[30]~202_combout ),
	.datad(\myif.out[30]~198_combout ),
	.cin(gnd),
	.combout(\myif.out[30]~203_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[30]~203 .lut_mask = 16'hBA98;
defparam \myif.out[30]~203 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N2
cycloneive_lcell_comb \myif.out[21]~207 (
// Equation(s):
// \myif.out[21]~207_combout  = \rdat1[21]~55_combout  $ (((\port_b~31_combout ) # ((fuifrtReplace_21 & \port_b~0_combout ))))

	.dataa(fuifrtReplace_21),
	.datab(port_b21),
	.datac(rdat1_21),
	.datad(port_b),
	.cin(gnd),
	.combout(\myif.out[21]~207_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[21]~207 .lut_mask = 16'h1E3C;
defparam \myif.out[21]~207 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N22
cycloneive_lcell_comb \myif.out[21]~209 (
// Equation(s):
// \myif.out[21]~209_combout  = (idex_ifaluop_o_1 & (((\Add1~42_combout )))) # (!idex_ifaluop_o_1 & ((\rdat1[21]~55_combout ) # ((\myif.out[21]~207_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(rdat1_21),
	.datac(\Add1~42_combout ),
	.datad(\myif.out[21]~207_combout ),
	.cin(gnd),
	.combout(\myif.out[21]~209_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[21]~209 .lut_mask = 16'hF5E4;
defparam \myif.out[21]~209 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N4
cycloneive_lcell_comb \myif.out[21]~210 (
// Equation(s):
// \myif.out[21]~210_combout  = (\myif.out[23]~135_combout  & (((\Add0~42_combout )))) # (!\myif.out[23]~135_combout  & ((idex_ifaluop_o_2) # ((\myif.out[21]~209_combout ))))

	.dataa(\myif.out[23]~135_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\myif.out[21]~209_combout ),
	.datad(\Add0~42_combout ),
	.cin(gnd),
	.combout(\myif.out[21]~210_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[21]~210 .lut_mask = 16'hFE54;
defparam \myif.out[21]~210 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N0
cycloneive_lcell_comb \myif.out[21]~219 (
// Equation(s):
// \myif.out[21]~219_combout  = (\myif.out[23]~135_combout  & ((\myif.out[23]~150_combout  & ((\myif.out[21]~207_combout ))) # (!\myif.out[23]~150_combout  & (\myif.out[21]~210_combout )))) # (!\myif.out[23]~135_combout  & (\myif.out[23]~150_combout ))

	.dataa(\myif.out[23]~135_combout ),
	.datab(\myif.out[23]~150_combout ),
	.datac(\myif.out[21]~210_combout ),
	.datad(\myif.out[21]~207_combout ),
	.cin(gnd),
	.combout(\myif.out[21]~219_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[21]~219 .lut_mask = 16'hEC64;
defparam \myif.out[21]~219 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N14
cycloneive_lcell_comb \ShiftLeft0~106 (
// Equation(s):
// \ShiftLeft0~106_combout  = (\port_b~10_combout  & ((\ShiftLeft0~60_combout ))) # (!\port_b~10_combout  & (\ShiftLeft0~63_combout ))

	.dataa(\ShiftLeft0~63_combout ),
	.datab(gnd),
	.datac(port_b6),
	.datad(\ShiftLeft0~60_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~106_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~106 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N24
cycloneive_lcell_comb \out~63 (
// Equation(s):
// \out~63_combout  = (\rdat1[21]~55_combout  & ((\port_b~31_combout ) # ((fuifrtReplace_21 & \port_b~0_combout ))))

	.dataa(fuifrtReplace_21),
	.datab(port_b21),
	.datac(rdat1_21),
	.datad(port_b),
	.cin(gnd),
	.combout(\out~63_combout ),
	.cout());
// synopsys translate_off
defparam \out~63 .lut_mask = 16'hE0C0;
defparam \out~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N26
cycloneive_lcell_comb \myif.out[21]~205 (
// Equation(s):
// \myif.out[21]~205_combout  = (\myif.out[13]~83_combout  & ((\myif.out[13]~84_combout  & (\out~63_combout )) # (!\myif.out[13]~84_combout  & ((\ShiftLeft0~88_combout ))))) # (!\myif.out[13]~83_combout  & (((\myif.out[13]~84_combout ))))

	.dataa(\myif.out[13]~83_combout ),
	.datab(\out~63_combout ),
	.datac(\ShiftLeft0~88_combout ),
	.datad(\myif.out[13]~84_combout ),
	.cin(gnd),
	.combout(\myif.out[21]~205_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[21]~205 .lut_mask = 16'hDDA0;
defparam \myif.out[21]~205 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N8
cycloneive_lcell_comb \myif.out[21]~206 (
// Equation(s):
// \myif.out[21]~206_combout  = (\myif.out[13]~82_combout  & (((\myif.out[21]~205_combout )))) # (!\myif.out[13]~82_combout  & ((\myif.out[21]~205_combout  & ((\ShiftLeft0~90_combout ))) # (!\myif.out[21]~205_combout  & (\ShiftLeft0~106_combout ))))

	.dataa(\ShiftLeft0~106_combout ),
	.datab(\myif.out[13]~82_combout ),
	.datac(\myif.out[21]~205_combout ),
	.datad(\ShiftLeft0~90_combout ),
	.cin(gnd),
	.combout(\myif.out[21]~206_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[21]~206 .lut_mask = 16'hF2C2;
defparam \myif.out[21]~206 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N28
cycloneive_lcell_comb \myif.out[21]~208 (
// Equation(s):
// \myif.out[21]~208_combout  = (idex_ifaluop_o_1 & (((!\myif.out[21]~207_combout  & !\rdat1[21]~55_combout )) # (!idex_ifaluop_o_2))) # (!idex_ifaluop_o_1 & (((idex_ifaluop_o_2))))

	.dataa(idex_ifaluop_o_1),
	.datab(\myif.out[21]~207_combout ),
	.datac(rdat1_21),
	.datad(idex_ifaluop_o_2),
	.cin(gnd),
	.combout(\myif.out[21]~208_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[21]~208 .lut_mask = 16'h57AA;
defparam \myif.out[21]~208 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N30
cycloneive_lcell_comb \myif.out[21]~211 (
// Equation(s):
// \myif.out[21]~211_combout  = (\port_b~31_combout ) # ((\port_b~0_combout  & fuifrtReplace_21))

	.dataa(port_b),
	.datab(gnd),
	.datac(port_b21),
	.datad(fuifrtReplace_21),
	.cin(gnd),
	.combout(\myif.out[21]~211_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[21]~211 .lut_mask = 16'hFAF0;
defparam \myif.out[21]~211 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N30
cycloneive_lcell_comb \myif.out[21]~216 (
// Equation(s):
// \myif.out[21]~216_combout  = (idex_ifaluop_o_1 & (!\rdat1[21]~55_combout  & (\Add1~42_combout  & !\myif.out[21]~211_combout ))) # (!idex_ifaluop_o_1 & ((\rdat1[21]~55_combout ) # ((\myif.out[21]~211_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(rdat1_21),
	.datac(\Add1~42_combout ),
	.datad(\myif.out[21]~211_combout ),
	.cin(gnd),
	.combout(\myif.out[21]~216_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[21]~216 .lut_mask = 16'h5564;
defparam \myif.out[21]~216 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N20
cycloneive_lcell_comb \myif.out[21]~213 (
// Equation(s):
// \myif.out[21]~213_combout  = (\port_b~31_combout ) # ((\rdat1[21]~55_combout ) # ((fuifrtReplace_21 & \port_b~0_combout )))

	.dataa(fuifrtReplace_21),
	.datab(port_b21),
	.datac(rdat1_21),
	.datad(port_b),
	.cin(gnd),
	.combout(\myif.out[21]~213_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[21]~213 .lut_mask = 16'hFEFC;
defparam \myif.out[21]~213 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N14
cycloneive_lcell_comb \myif.out[21]~214 (
// Equation(s):
// \myif.out[21]~214_combout  = (idex_ifaluop_o_1 & (\Add1~42_combout  & ((!\myif.out[21]~213_combout ) # (!idex_ifaluop_o_2)))) # (!idex_ifaluop_o_1 & (idex_ifaluop_o_2 & ((\myif.out[21]~213_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(idex_ifaluop_o_2),
	.datac(\Add1~42_combout ),
	.datad(\myif.out[21]~213_combout ),
	.cin(gnd),
	.combout(\myif.out[21]~214_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[21]~214 .lut_mask = 16'h64A0;
defparam \myif.out[21]~214 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N16
cycloneive_lcell_comb \myif.out[21]~215 (
// Equation(s):
// \myif.out[21]~215_combout  = (\ShiftRight0~79_combout  & (\myif.out[21]~212_combout )) # (!\ShiftRight0~79_combout  & ((\myif.out[21]~214_combout )))

	.dataa(\myif.out[21]~212_combout ),
	.datab(gnd),
	.datac(\myif.out[21]~214_combout ),
	.datad(\ShiftRight0~79_combout ),
	.cin(gnd),
	.combout(\myif.out[21]~215_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[21]~215 .lut_mask = 16'hAAF0;
defparam \myif.out[21]~215 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N12
cycloneive_lcell_comb \myif.out[21]~217 (
// Equation(s):
// \myif.out[21]~217_combout  = (idex_ifaluop_o_2 & (\myif.out[21]~216_combout )) # (!idex_ifaluop_o_2 & ((\myif.out[21]~215_combout )))

	.dataa(gnd),
	.datab(idex_ifaluop_o_2),
	.datac(\myif.out[21]~216_combout ),
	.datad(\myif.out[21]~215_combout ),
	.cin(gnd),
	.combout(\myif.out[21]~217_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[21]~217 .lut_mask = 16'hF3C0;
defparam \myif.out[21]~217 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N18
cycloneive_lcell_comb \myif.out[21]~218 (
// Equation(s):
// \myif.out[21]~218_combout  = (\myif.out[13]~23_combout  & (((\myif.out[21]~217_combout )))) # (!\myif.out[13]~23_combout  & (\myif.out[21]~208_combout  & (\myif.out[21]~210_combout )))

	.dataa(\myif.out[13]~23_combout ),
	.datab(\myif.out[21]~208_combout ),
	.datac(\myif.out[21]~210_combout ),
	.datad(\myif.out[21]~217_combout ),
	.cin(gnd),
	.combout(\myif.out[21]~218_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[21]~218 .lut_mask = 16'hEA40;
defparam \myif.out[21]~218 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N14
cycloneive_lcell_comb \out~66 (
// Equation(s):
// \out~66_combout  = \rdat1[31]~35_combout  $ (((\port_b~19_combout ) # ((\port_b~0_combout  & fuifrtReplace_31))))

	.dataa(port_b),
	.datab(port_b9),
	.datac(rdat1_311),
	.datad(fuifrtReplace_31),
	.cin(gnd),
	.combout(\out~66_combout ),
	.cout());
// synopsys translate_off
defparam \out~66 .lut_mask = 16'h1E3C;
defparam \out~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N26
cycloneive_lcell_comb \out~64 (
// Equation(s):
// \out~64_combout  = (\port_b~19_combout ) # ((\rdat1[31]~35_combout ) # ((\port_b~0_combout  & fuifrtReplace_31)))

	.dataa(port_b),
	.datab(port_b9),
	.datac(rdat1_311),
	.datad(fuifrtReplace_31),
	.cin(gnd),
	.combout(\out~64_combout ),
	.cout());
// synopsys translate_off
defparam \out~64 .lut_mask = 16'hFEFC;
defparam \out~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N14
cycloneive_lcell_comb \myif.negative~1 (
// Equation(s):
// \myif.negative~1_combout  = (idex_ifaluop_o_2 & ((\out~64_combout ) # ((!\myif.out[13]~23_combout )))) # (!idex_ifaluop_o_2 & (((\ShiftRight0~96_combout  & \myif.out[13]~23_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\out~64_combout ),
	.datac(\ShiftRight0~96_combout ),
	.datad(\myif.out[13]~23_combout ),
	.cin(gnd),
	.combout(\myif.negative~1_combout ),
	.cout());
// synopsys translate_off
defparam \myif.negative~1 .lut_mask = 16'hD8AA;
defparam \myif.negative~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N30
cycloneive_lcell_comb \Add1~62 (
// Equation(s):
// \Add1~62_combout  = \rdat1[31]~35_combout  $ (\Add1~61  $ (!\port_b~20_combout ))

	.dataa(gnd),
	.datab(rdat1_311),
	.datac(gnd),
	.datad(port_b10),
	.cin(\Add1~61 ),
	.combout(\Add1~62_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~62 .lut_mask = 16'h3CC3;
defparam \Add1~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N4
cycloneive_lcell_comb \myif.negative~2 (
// Equation(s):
// \myif.negative~2_combout  = (idex_ifaluop_o_1 & ((\myif.negative~1_combout  & ((!\out~64_combout ))) # (!\myif.negative~1_combout  & (\Add1~62_combout )))) # (!idex_ifaluop_o_1 & (\myif.negative~1_combout ))

	.dataa(idex_ifaluop_o_1),
	.datab(\myif.negative~1_combout ),
	.datac(\Add1~62_combout ),
	.datad(\out~64_combout ),
	.cin(gnd),
	.combout(\myif.negative~2_combout ),
	.cout());
// synopsys translate_off
defparam \myif.negative~2 .lut_mask = 16'h64EC;
defparam \myif.negative~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N26
cycloneive_lcell_comb \myif.negative~5 (
// Equation(s):
// \myif.negative~5_combout  = (\myif.out[13]~84_combout  & ((\out~65_combout ) # ((!\myif.out[13]~83_combout )))) # (!\myif.out[13]~84_combout  & (((\myif.out[13]~83_combout  & \ShiftLeft0~100_combout ))))

	.dataa(\out~65_combout ),
	.datab(\myif.out[13]~84_combout ),
	.datac(\myif.out[13]~83_combout ),
	.datad(\ShiftLeft0~100_combout ),
	.cin(gnd),
	.combout(\myif.negative~5_combout ),
	.cout());
// synopsys translate_off
defparam \myif.negative~5 .lut_mask = 16'hBC8C;
defparam \myif.negative~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N8
cycloneive_lcell_comb \myif.negative~6 (
// Equation(s):
// \myif.negative~6_combout  = (\myif.out[13]~82_combout  & (((\myif.negative~5_combout )))) # (!\myif.out[13]~82_combout  & ((\myif.negative~5_combout  & ((\ShiftLeft0~101_combout ))) # (!\myif.negative~5_combout  & (\myif.negative~4_combout ))))

	.dataa(\myif.negative~4_combout ),
	.datab(\myif.out[13]~82_combout ),
	.datac(\myif.negative~5_combout ),
	.datad(\ShiftLeft0~101_combout ),
	.cin(gnd),
	.combout(\myif.negative~6_combout ),
	.cout());
// synopsys translate_off
defparam \myif.negative~6 .lut_mask = 16'hF2C2;
defparam \myif.negative~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N30
cycloneive_lcell_comb \Add0~62 (
// Equation(s):
// \Add0~62_combout  = \port_b~20_combout  $ (\Add0~61  $ (\rdat1[31]~35_combout ))

	.dataa(port_b10),
	.datab(gnd),
	.datac(gnd),
	.datad(rdat1_311),
	.cin(\Add0~61 ),
	.combout(\Add0~62_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~62 .lut_mask = 16'hA55A;
defparam \Add0~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N18
cycloneive_lcell_comb \myif.negative~7 (
// Equation(s):
// \myif.negative~7_combout  = (\myif.out[23]~150_combout  & (\myif.out[23]~135_combout )) # (!\myif.out[23]~150_combout  & ((\myif.out[23]~135_combout  & ((\Add0~62_combout ))) # (!\myif.out[23]~135_combout  & (\myif.negative~6_combout ))))

	.dataa(\myif.out[23]~150_combout ),
	.datab(\myif.out[23]~135_combout ),
	.datac(\myif.negative~6_combout ),
	.datad(\Add0~62_combout ),
	.cin(gnd),
	.combout(\myif.negative~7_combout ),
	.cout());
// synopsys translate_off
defparam \myif.negative~7 .lut_mask = 16'hDC98;
defparam \myif.negative~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N24
cycloneive_lcell_comb \out~69 (
// Equation(s):
// \out~69_combout  = \rdat1[22]~51_combout  $ (((\port_b~33_combout ) # ((fuifrtReplace_22 & \port_b~0_combout ))))

	.dataa(port_b23),
	.datab(rdat1_22),
	.datac(fuifrtReplace_22),
	.datad(port_b),
	.cin(gnd),
	.combout(\out~69_combout ),
	.cout());
// synopsys translate_off
defparam \out~69 .lut_mask = 16'h3666;
defparam \out~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N2
cycloneive_lcell_comb \out~68 (
// Equation(s):
// \out~68_combout  = (\rdat1[22]~51_combout  & ((\port_b~33_combout ) # ((fuifrtReplace_22 & \port_b~0_combout ))))

	.dataa(port_b23),
	.datab(fuifrtReplace_22),
	.datac(rdat1_22),
	.datad(port_b),
	.cin(gnd),
	.combout(\out~68_combout ),
	.cout());
// synopsys translate_off
defparam \out~68 .lut_mask = 16'hE0A0;
defparam \out~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N18
cycloneive_lcell_comb \myif.out[22]~223 (
// Equation(s):
// \myif.out[22]~223_combout  = (\myif.out[13]~84_combout  & (((\out~68_combout ) # (!\myif.out[13]~83_combout )))) # (!\myif.out[13]~84_combout  & (\ShiftLeft0~20_combout  & ((\myif.out[13]~83_combout ))))

	.dataa(\myif.out[13]~84_combout ),
	.datab(\ShiftLeft0~20_combout ),
	.datac(\out~68_combout ),
	.datad(\myif.out[13]~83_combout ),
	.cin(gnd),
	.combout(\myif.out[22]~223_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[22]~223 .lut_mask = 16'hE4AA;
defparam \myif.out[22]~223 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N8
cycloneive_lcell_comb \myif.out[22]~224 (
// Equation(s):
// \myif.out[22]~224_combout  = (\myif.out[22]~223_combout  & ((\ShiftLeft0~93_combout ) # ((\myif.out[13]~82_combout )))) # (!\myif.out[22]~223_combout  & (((\ShiftLeft0~105_combout  & !\myif.out[13]~82_combout ))))

	.dataa(\ShiftLeft0~93_combout ),
	.datab(\myif.out[22]~223_combout ),
	.datac(\ShiftLeft0~105_combout ),
	.datad(\myif.out[13]~82_combout ),
	.cin(gnd),
	.combout(\myif.out[22]~224_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[22]~224 .lut_mask = 16'hCCB8;
defparam \myif.out[22]~224 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N20
cycloneive_lcell_comb \out~67 (
// Equation(s):
// \out~67_combout  = (\port_b~33_combout ) # ((\rdat1[22]~51_combout ) # ((fuifrtReplace_22 & \port_b~0_combout )))

	.dataa(port_b23),
	.datab(fuifrtReplace_22),
	.datac(rdat1_22),
	.datad(port_b),
	.cin(gnd),
	.combout(\out~67_combout ),
	.cout());
// synopsys translate_off
defparam \out~67 .lut_mask = 16'hFEFA;
defparam \out~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N26
cycloneive_lcell_comb \myif.out[22]~221 (
// Equation(s):
// \myif.out[22]~221_combout  = (idex_ifaluop_o_2 & ((\out~67_combout ) # ((!\myif.out[13]~23_combout )))) # (!idex_ifaluop_o_2 & (((\myif.out[13]~23_combout  & \ShiftRight0~53_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\out~67_combout ),
	.datac(\myif.out[13]~23_combout ),
	.datad(\ShiftRight0~53_combout ),
	.cin(gnd),
	.combout(\myif.out[22]~221_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[22]~221 .lut_mask = 16'hDA8A;
defparam \myif.out[22]~221 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N16
cycloneive_lcell_comb \myif.out[22]~222 (
// Equation(s):
// \myif.out[22]~222_combout  = (idex_ifaluop_o_1 & ((\myif.out[22]~221_combout  & (!\out~67_combout )) # (!\myif.out[22]~221_combout  & ((\Add1~44_combout ))))) # (!idex_ifaluop_o_1 & (((\myif.out[22]~221_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(\out~67_combout ),
	.datac(\myif.out[22]~221_combout ),
	.datad(\Add1~44_combout ),
	.cin(gnd),
	.combout(\myif.out[22]~222_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[22]~222 .lut_mask = 16'h7A70;
defparam \myif.out[22]~222 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N22
cycloneive_lcell_comb \myif.out[22]~225 (
// Equation(s):
// \myif.out[22]~225_combout  = (\myif.out[23]~150_combout  & ((\myif.out[23]~135_combout ) # ((\myif.out[22]~222_combout )))) # (!\myif.out[23]~150_combout  & (!\myif.out[23]~135_combout  & (\myif.out[22]~224_combout )))

	.dataa(\myif.out[23]~150_combout ),
	.datab(\myif.out[23]~135_combout ),
	.datac(\myif.out[22]~224_combout ),
	.datad(\myif.out[22]~222_combout ),
	.cin(gnd),
	.combout(\myif.out[22]~225_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[22]~225 .lut_mask = 16'hBA98;
defparam \myif.out[22]~225 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N10
cycloneive_lcell_comb \out~72 (
// Equation(s):
// \out~72_combout  = \rdat1[20]~57_combout  $ (((\port_b~29_combout ) # ((\port_b~0_combout  & fuifrtReplace_20))))

	.dataa(rdat1_20),
	.datab(port_b),
	.datac(port_b19),
	.datad(fuifrtReplace_20),
	.cin(gnd),
	.combout(\out~72_combout ),
	.cout());
// synopsys translate_off
defparam \out~72 .lut_mask = 16'h565A;
defparam \out~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N4
cycloneive_lcell_comb \ShiftLeft0~29 (
// Equation(s):
// \ShiftLeft0~29_combout  = (!\port_b~7_combout  & ((\port_b~4_combout  & (\rdat1[14]~23_combout )) # (!\port_b~4_combout  & ((\rdat1[16]~19_combout )))))

	.dataa(rdat1_14),
	.datab(port_b4),
	.datac(port_b2),
	.datad(rdat1_16),
	.cin(gnd),
	.combout(\ShiftLeft0~29_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~29 .lut_mask = 16'h2320;
defparam \ShiftLeft0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N6
cycloneive_lcell_comb \ShiftLeft0~33 (
// Equation(s):
// \ShiftLeft0~33_combout  = (\ShiftLeft0~31_combout ) # ((\port_b~7_combout  & \ShiftLeft0~32_combout ))

	.dataa(\ShiftLeft0~31_combout ),
	.datab(port_b4),
	.datac(gnd),
	.datad(\ShiftLeft0~32_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~33_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~33 .lut_mask = 16'hEEAA;
defparam \ShiftLeft0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N30
cycloneive_lcell_comb \ShiftLeft0~108 (
// Equation(s):
// \ShiftLeft0~108_combout  = (\port_b~10_combout  & ((\ShiftLeft0~28_combout ) # ((\ShiftLeft0~29_combout )))) # (!\port_b~10_combout  & (((\ShiftLeft0~33_combout ))))

	.dataa(port_b6),
	.datab(\ShiftLeft0~28_combout ),
	.datac(\ShiftLeft0~29_combout ),
	.datad(\ShiftLeft0~33_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~108_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~108 .lut_mask = 16'hFDA8;
defparam \ShiftLeft0~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N28
cycloneive_lcell_comb \myif.out[20]~229 (
// Equation(s):
// \myif.out[20]~229_combout  = (\myif.out[13]~84_combout  & ((\out~71_combout ) # ((!\myif.out[13]~83_combout )))) # (!\myif.out[13]~84_combout  & (((\ShiftLeft0~24_combout  & \myif.out[13]~83_combout ))))

	.dataa(\out~71_combout ),
	.datab(\myif.out[13]~84_combout ),
	.datac(\ShiftLeft0~24_combout ),
	.datad(\myif.out[13]~83_combout ),
	.cin(gnd),
	.combout(\myif.out[20]~229_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[20]~229 .lut_mask = 16'hB8CC;
defparam \myif.out[20]~229 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N26
cycloneive_lcell_comb \myif.out[20]~230 (
// Equation(s):
// \myif.out[20]~230_combout  = (\myif.out[13]~82_combout  & (((\myif.out[20]~229_combout )))) # (!\myif.out[13]~82_combout  & ((\myif.out[20]~229_combout  & (\ShiftLeft0~96_combout )) # (!\myif.out[20]~229_combout  & ((\ShiftLeft0~108_combout )))))

	.dataa(\myif.out[13]~82_combout ),
	.datab(\ShiftLeft0~96_combout ),
	.datac(\ShiftLeft0~108_combout ),
	.datad(\myif.out[20]~229_combout ),
	.cin(gnd),
	.combout(\myif.out[20]~230_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[20]~230 .lut_mask = 16'hEE50;
defparam \myif.out[20]~230 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N14
cycloneive_lcell_comb \out~70 (
// Equation(s):
// \out~70_combout  = (\port_b~29_combout ) # ((\rdat1[20]~57_combout ) # ((\port_b~0_combout  & fuifrtReplace_20)))

	.dataa(port_b19),
	.datab(port_b),
	.datac(rdat1_20),
	.datad(fuifrtReplace_20),
	.cin(gnd),
	.combout(\out~70_combout ),
	.cout());
// synopsys translate_off
defparam \out~70 .lut_mask = 16'hFEFA;
defparam \out~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N8
cycloneive_lcell_comb \myif.out[20]~227 (
// Equation(s):
// \myif.out[20]~227_combout  = (idex_ifaluop_o_2 & (((\out~70_combout )) # (!\myif.out[13]~23_combout ))) # (!idex_ifaluop_o_2 & (\myif.out[13]~23_combout  & ((\ShiftRight0~68_combout ))))

	.dataa(idex_ifaluop_o_2),
	.datab(\myif.out[13]~23_combout ),
	.datac(\out~70_combout ),
	.datad(\ShiftRight0~68_combout ),
	.cin(gnd),
	.combout(\myif.out[20]~227_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[20]~227 .lut_mask = 16'hE6A2;
defparam \myif.out[20]~227 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N18
cycloneive_lcell_comb \myif.out[20]~228 (
// Equation(s):
// \myif.out[20]~228_combout  = (idex_ifaluop_o_1 & ((\myif.out[20]~227_combout  & (!\out~70_combout )) # (!\myif.out[20]~227_combout  & ((\Add1~40_combout ))))) # (!idex_ifaluop_o_1 & (((\myif.out[20]~227_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(\out~70_combout ),
	.datac(\myif.out[20]~227_combout ),
	.datad(\Add1~40_combout ),
	.cin(gnd),
	.combout(\myif.out[20]~228_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[20]~228 .lut_mask = 16'h7A70;
defparam \myif.out[20]~228 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N20
cycloneive_lcell_comb \myif.out[20]~231 (
// Equation(s):
// \myif.out[20]~231_combout  = (\myif.out[23]~135_combout  & (\myif.out[23]~150_combout )) # (!\myif.out[23]~135_combout  & ((\myif.out[23]~150_combout  & ((\myif.out[20]~228_combout ))) # (!\myif.out[23]~150_combout  & (\myif.out[20]~230_combout ))))

	.dataa(\myif.out[23]~135_combout ),
	.datab(\myif.out[23]~150_combout ),
	.datac(\myif.out[20]~230_combout ),
	.datad(\myif.out[20]~228_combout ),
	.cin(gnd),
	.combout(\myif.out[20]~231_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[20]~231 .lut_mask = 16'hDC98;
defparam \myif.out[20]~231 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N4
cycloneive_lcell_comb \myif.out[0]~237 (
// Equation(s):
// \myif.out[0]~237_combout  = (idex_ifaluop_o_0 & (!idex_ifaluop_o_2)) # (!idex_ifaluop_o_0 & ((\Add0~0_combout )))

	.dataa(gnd),
	.datab(idex_ifaluop_o_2),
	.datac(idex_ifaluop_o_0),
	.datad(\Add0~0_combout ),
	.cin(gnd),
	.combout(\myif.out[0]~237_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[0]~237 .lut_mask = 16'h3F30;
defparam \myif.out[0]~237 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N10
cycloneive_lcell_comb \out~73 (
// Equation(s):
// \out~73_combout  = (\port_b~6_combout ) # ((\rdat1[0]~3_combout ) # ((fuifrtReplace_0 & \port_b~0_combout )))

	.dataa(fuifrtReplace_0),
	.datab(port_b),
	.datac(port_b3),
	.datad(rdat1_0),
	.cin(gnd),
	.combout(\out~73_combout ),
	.cout());
// synopsys translate_off
defparam \out~73 .lut_mask = 16'hFFF8;
defparam \out~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N22
cycloneive_lcell_comb \myif.out[0]~238 (
// Equation(s):
// \myif.out[0]~238_combout  = (\myif.out[0]~237_combout  & ((\Add1~0_combout ) # ((!idex_ifaluop_o_0)))) # (!\myif.out[0]~237_combout  & (((idex_ifaluop_o_0 & !\out~73_combout ))))

	.dataa(\Add1~0_combout ),
	.datab(\myif.out[0]~237_combout ),
	.datac(idex_ifaluop_o_0),
	.datad(\out~73_combout ),
	.cin(gnd),
	.combout(\myif.out[0]~238_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[0]~238 .lut_mask = 16'h8CBC;
defparam \myif.out[0]~238 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N30
cycloneive_lcell_comb \ShiftLeft0~102 (
// Equation(s):
// \ShiftLeft0~102_combout  = (!\port_b~14_combout  & (!\port_b~10_combout  & \ShiftLeft0~21_combout ))

	.dataa(gnd),
	.datab(port_b7),
	.datac(port_b6),
	.datad(\ShiftLeft0~21_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~102_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~102 .lut_mask = 16'h0300;
defparam \ShiftLeft0~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N26
cycloneive_lcell_comb \myif.out[0]~235 (
// Equation(s):
// \myif.out[0]~235_combout  = (\myif.out[0]~234_combout  & ((idex_ifaluop_o_2) # ((\ShiftLeft0~102_combout  & !\ShiftLeft0~11_combout ))))

	.dataa(\myif.out[0]~234_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\ShiftLeft0~102_combout ),
	.datad(\ShiftLeft0~11_combout ),
	.cin(gnd),
	.combout(\myif.out[0]~235_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[0]~235 .lut_mask = 16'h88A8;
defparam \myif.out[0]~235 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N12
cycloneive_lcell_comb \ShiftRight0~111 (
// Equation(s):
// \ShiftRight0~111_combout  = (!\ShiftLeft0~11_combout  & ((\port_b~17_combout  & ((\ShiftRight0~102_combout ))) # (!\port_b~17_combout  & (\ShiftRight0~110_combout ))))

	.dataa(\ShiftRight0~110_combout ),
	.datab(\ShiftLeft0~11_combout ),
	.datac(port_b8),
	.datad(\ShiftRight0~102_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~111_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~111 .lut_mask = 16'h3202;
defparam \ShiftRight0~111 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N8
cycloneive_lcell_comb \myif.out[0]~236 (
// Equation(s):
// \myif.out[0]~236_combout  = (idex_ifaluop_o_0 & ((\myif.out[0]~235_combout  & (\out~73_combout )) # (!\myif.out[0]~235_combout  & ((\ShiftRight0~111_combout ))))) # (!idex_ifaluop_o_0 & (((\myif.out[0]~235_combout ))))

	.dataa(\out~73_combout ),
	.datab(idex_ifaluop_o_0),
	.datac(\myif.out[0]~235_combout ),
	.datad(\ShiftRight0~111_combout ),
	.cin(gnd),
	.combout(\myif.out[0]~236_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[0]~236 .lut_mask = 16'hBCB0;
defparam \myif.out[0]~236 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N0
cycloneive_lcell_comb \LessThan1~1 (
// Equation(s):
// \LessThan1~1_cout  = CARRY((\port_b~7_combout  & !\rdat1[0]~3_combout ))

	.dataa(port_b4),
	.datab(rdat1_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan1~1_cout ));
// synopsys translate_off
defparam \LessThan1~1 .lut_mask = 16'h0022;
defparam \LessThan1~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N2
cycloneive_lcell_comb \LessThan1~3 (
// Equation(s):
// \LessThan1~3_cout  = CARRY((\rdat1[1]~1_combout  & ((!\LessThan1~1_cout ) # (!\port_b~4_combout ))) # (!\rdat1[1]~1_combout  & (!\port_b~4_combout  & !\LessThan1~1_cout )))

	.dataa(rdat1_1),
	.datab(port_b2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~1_cout ),
	.combout(),
	.cout(\LessThan1~3_cout ));
// synopsys translate_off
defparam \LessThan1~3 .lut_mask = 16'h002B;
defparam \LessThan1~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N4
cycloneive_lcell_comb \LessThan1~5 (
// Equation(s):
// \LessThan1~5_cout  = CARRY((\port_b~10_combout  & ((!\LessThan1~3_cout ) # (!\rdat1[2]~5_combout ))) # (!\port_b~10_combout  & (!\rdat1[2]~5_combout  & !\LessThan1~3_cout )))

	.dataa(port_b6),
	.datab(rdat1_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~3_cout ),
	.combout(),
	.cout(\LessThan1~5_cout ));
// synopsys translate_off
defparam \LessThan1~5 .lut_mask = 16'h002B;
defparam \LessThan1~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N6
cycloneive_lcell_comb \LessThan1~7 (
// Equation(s):
// \LessThan1~7_cout  = CARRY((\port_b~14_combout  & (\rdat1[3]~9_combout  & !\LessThan1~5_cout )) # (!\port_b~14_combout  & ((\rdat1[3]~9_combout ) # (!\LessThan1~5_cout ))))

	.dataa(port_b7),
	.datab(rdat1_31),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~5_cout ),
	.combout(),
	.cout(\LessThan1~7_cout ));
// synopsys translate_off
defparam \LessThan1~7 .lut_mask = 16'h004D;
defparam \LessThan1~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N8
cycloneive_lcell_comb \LessThan1~9 (
// Equation(s):
// \LessThan1~9_cout  = CARRY((\rdat1[4]~7_combout  & (\port_b~17_combout  & !\LessThan1~7_cout )) # (!\rdat1[4]~7_combout  & ((\port_b~17_combout ) # (!\LessThan1~7_cout ))))

	.dataa(rdat1_41),
	.datab(port_b8),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~7_cout ),
	.combout(),
	.cout(\LessThan1~9_cout ));
// synopsys translate_off
defparam \LessThan1~9 .lut_mask = 16'h004D;
defparam \LessThan1~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N10
cycloneive_lcell_comb \LessThan1~11 (
// Equation(s):
// \LessThan1~11_cout  = CARRY((\port_b~44_combout  & (\rdat1[5]~17_combout  & !\LessThan1~9_cout )) # (!\port_b~44_combout  & ((\rdat1[5]~17_combout ) # (!\LessThan1~9_cout ))))

	.dataa(port_b34),
	.datab(rdat1_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~9_cout ),
	.combout(),
	.cout(\LessThan1~11_cout ));
// synopsys translate_off
defparam \LessThan1~11 .lut_mask = 16'h004D;
defparam \LessThan1~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N12
cycloneive_lcell_comb \LessThan1~13 (
// Equation(s):
// \LessThan1~13_cout  = CARRY((\port_b~46_combout  & ((!\LessThan1~11_cout ) # (!\rdat1[6]~15_combout ))) # (!\port_b~46_combout  & (!\rdat1[6]~15_combout  & !\LessThan1~11_cout )))

	.dataa(port_b36),
	.datab(rdat1_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~11_cout ),
	.combout(),
	.cout(\LessThan1~13_cout ));
// synopsys translate_off
defparam \LessThan1~13 .lut_mask = 16'h002B;
defparam \LessThan1~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N14
cycloneive_lcell_comb \LessThan1~15 (
// Equation(s):
// \LessThan1~15_cout  = CARRY((\rdat1[7]~13_combout  & ((!\LessThan1~13_cout ) # (!\port_b~48_combout ))) # (!\rdat1[7]~13_combout  & (!\port_b~48_combout  & !\LessThan1~13_cout )))

	.dataa(rdat1_7),
	.datab(port_b38),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~13_cout ),
	.combout(),
	.cout(\LessThan1~15_cout ));
// synopsys translate_off
defparam \LessThan1~15 .lut_mask = 16'h002B;
defparam \LessThan1~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N16
cycloneive_lcell_comb \LessThan1~17 (
// Equation(s):
// \LessThan1~17_cout  = CARRY((\rdat1[8]~11_combout  & (\port_b~50_combout  & !\LessThan1~15_cout )) # (!\rdat1[8]~11_combout  & ((\port_b~50_combout ) # (!\LessThan1~15_cout ))))

	.dataa(rdat1_8),
	.datab(port_b40),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~15_cout ),
	.combout(),
	.cout(\LessThan1~17_cout ));
// synopsys translate_off
defparam \LessThan1~17 .lut_mask = 16'h004D;
defparam \LessThan1~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N18
cycloneive_lcell_comb \LessThan1~19 (
// Equation(s):
// \LessThan1~19_cout  = CARRY((\port_b~60_combout  & (\rdat1[9]~33_combout  & !\LessThan1~17_cout )) # (!\port_b~60_combout  & ((\rdat1[9]~33_combout ) # (!\LessThan1~17_cout ))))

	.dataa(port_b50),
	.datab(rdat1_9),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~17_cout ),
	.combout(),
	.cout(\LessThan1~19_cout ));
// synopsys translate_off
defparam \LessThan1~19 .lut_mask = 16'h004D;
defparam \LessThan1~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N20
cycloneive_lcell_comb \LessThan1~21 (
// Equation(s):
// \LessThan1~21_cout  = CARRY((\port_b~65_combout  & ((!\LessThan1~19_cout ) # (!\rdat1[10]~31_combout ))) # (!\port_b~65_combout  & (!\rdat1[10]~31_combout  & !\LessThan1~19_cout )))

	.dataa(port_b55),
	.datab(rdat1_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~19_cout ),
	.combout(),
	.cout(\LessThan1~21_cout ));
// synopsys translate_off
defparam \LessThan1~21 .lut_mask = 16'h002B;
defparam \LessThan1~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N22
cycloneive_lcell_comb \LessThan1~23 (
// Equation(s):
// \LessThan1~23_cout  = CARRY((\port_b~67_combout  & (\rdat1[11]~29_combout  & !\LessThan1~21_cout )) # (!\port_b~67_combout  & ((\rdat1[11]~29_combout ) # (!\LessThan1~21_cout ))))

	.dataa(port_b57),
	.datab(rdat1_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~21_cout ),
	.combout(),
	.cout(\LessThan1~23_cout ));
// synopsys translate_off
defparam \LessThan1~23 .lut_mask = 16'h004D;
defparam \LessThan1~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N24
cycloneive_lcell_comb \LessThan1~25 (
// Equation(s):
// \LessThan1~25_cout  = CARRY((\rdat1[12]~27_combout  & (\port_b~72_combout  & !\LessThan1~23_cout )) # (!\rdat1[12]~27_combout  & ((\port_b~72_combout ) # (!\LessThan1~23_cout ))))

	.dataa(rdat1_12),
	.datab(port_b62),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~23_cout ),
	.combout(),
	.cout(\LessThan1~25_cout ));
// synopsys translate_off
defparam \LessThan1~25 .lut_mask = 16'h004D;
defparam \LessThan1~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N26
cycloneive_lcell_comb \LessThan1~27 (
// Equation(s):
// \LessThan1~27_cout  = CARRY((\rdat1[13]~25_combout  & ((!\LessThan1~25_cout ) # (!\port_b~70_combout ))) # (!\rdat1[13]~25_combout  & (!\port_b~70_combout  & !\LessThan1~25_cout )))

	.dataa(rdat1_13),
	.datab(port_b60),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~25_cout ),
	.combout(),
	.cout(\LessThan1~27_cout ));
// synopsys translate_off
defparam \LessThan1~27 .lut_mask = 16'h002B;
defparam \LessThan1~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N28
cycloneive_lcell_comb \LessThan1~29 (
// Equation(s):
// \LessThan1~29_cout  = CARRY((\rdat1[14]~23_combout  & (\port_b~71_combout  & !\LessThan1~27_cout )) # (!\rdat1[14]~23_combout  & ((\port_b~71_combout ) # (!\LessThan1~27_cout ))))

	.dataa(rdat1_14),
	.datab(port_b61),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~27_cout ),
	.combout(),
	.cout(\LessThan1~29_cout ));
// synopsys translate_off
defparam \LessThan1~29 .lut_mask = 16'h004D;
defparam \LessThan1~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N30
cycloneive_lcell_comb \LessThan1~31 (
// Equation(s):
// \LessThan1~31_cout  = CARRY((\port_b~63_combout  & (\rdat1[15]~21_combout  & !\LessThan1~29_cout )) # (!\port_b~63_combout  & ((\rdat1[15]~21_combout ) # (!\LessThan1~29_cout ))))

	.dataa(port_b53),
	.datab(rdat1_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~29_cout ),
	.combout(),
	.cout(\LessThan1~31_cout ));
// synopsys translate_off
defparam \LessThan1~31 .lut_mask = 16'h004D;
defparam \LessThan1~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N0
cycloneive_lcell_comb \LessThan1~33 (
// Equation(s):
// \LessThan1~33_cout  = CARRY((\port_b~22_combout  & ((!\LessThan1~31_cout ) # (!\rdat1[16]~19_combout ))) # (!\port_b~22_combout  & (!\rdat1[16]~19_combout  & !\LessThan1~31_cout )))

	.dataa(port_b12),
	.datab(rdat1_16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~31_cout ),
	.combout(),
	.cout(\LessThan1~33_cout ));
// synopsys translate_off
defparam \LessThan1~33 .lut_mask = 16'h002B;
defparam \LessThan1~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N2
cycloneive_lcell_comb \LessThan1~35 (
// Equation(s):
// \LessThan1~35_cout  = CARRY((\rdat1[17]~63_combout  & ((!\LessThan1~33_cout ) # (!\port_b~24_combout ))) # (!\rdat1[17]~63_combout  & (!\port_b~24_combout  & !\LessThan1~33_cout )))

	.dataa(rdat1_17),
	.datab(port_b14),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~33_cout ),
	.combout(),
	.cout(\LessThan1~35_cout ));
// synopsys translate_off
defparam \LessThan1~35 .lut_mask = 16'h002B;
defparam \LessThan1~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N4
cycloneive_lcell_comb \LessThan1~37 (
// Equation(s):
// \LessThan1~37_cout  = CARRY((\port_b~26_combout  & ((!\LessThan1~35_cout ) # (!\rdat1[18]~59_combout ))) # (!\port_b~26_combout  & (!\rdat1[18]~59_combout  & !\LessThan1~35_cout )))

	.dataa(port_b16),
	.datab(rdat1_18),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~35_cout ),
	.combout(),
	.cout(\LessThan1~37_cout ));
// synopsys translate_off
defparam \LessThan1~37 .lut_mask = 16'h002B;
defparam \LessThan1~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N6
cycloneive_lcell_comb \LessThan1~39 (
// Equation(s):
// \LessThan1~39_cout  = CARRY((\rdat1[19]~61_combout  & ((!\LessThan1~37_cout ) # (!\port_b~28_combout ))) # (!\rdat1[19]~61_combout  & (!\port_b~28_combout  & !\LessThan1~37_cout )))

	.dataa(rdat1_19),
	.datab(port_b18),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~37_cout ),
	.combout(),
	.cout(\LessThan1~39_cout ));
// synopsys translate_off
defparam \LessThan1~39 .lut_mask = 16'h002B;
defparam \LessThan1~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N8
cycloneive_lcell_comb \LessThan1~41 (
// Equation(s):
// \LessThan1~41_cout  = CARRY((\port_b~30_combout  & ((!\LessThan1~39_cout ) # (!\rdat1[20]~57_combout ))) # (!\port_b~30_combout  & (!\rdat1[20]~57_combout  & !\LessThan1~39_cout )))

	.dataa(port_b20),
	.datab(rdat1_20),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~39_cout ),
	.combout(),
	.cout(\LessThan1~41_cout ));
// synopsys translate_off
defparam \LessThan1~41 .lut_mask = 16'h002B;
defparam \LessThan1~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N10
cycloneive_lcell_comb \LessThan1~43 (
// Equation(s):
// \LessThan1~43_cout  = CARRY((\port_b~32_combout  & (\rdat1[21]~55_combout  & !\LessThan1~41_cout )) # (!\port_b~32_combout  & ((\rdat1[21]~55_combout ) # (!\LessThan1~41_cout ))))

	.dataa(port_b22),
	.datab(rdat1_21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~41_cout ),
	.combout(),
	.cout(\LessThan1~43_cout ));
// synopsys translate_off
defparam \LessThan1~43 .lut_mask = 16'h004D;
defparam \LessThan1~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N12
cycloneive_lcell_comb \LessThan1~45 (
// Equation(s):
// \LessThan1~45_cout  = CARRY((\port_b~34_combout  & ((!\LessThan1~43_cout ) # (!\rdat1[22]~51_combout ))) # (!\port_b~34_combout  & (!\rdat1[22]~51_combout  & !\LessThan1~43_cout )))

	.dataa(port_b24),
	.datab(rdat1_22),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~43_cout ),
	.combout(),
	.cout(\LessThan1~45_cout ));
// synopsys translate_off
defparam \LessThan1~45 .lut_mask = 16'h002B;
defparam \LessThan1~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N14
cycloneive_lcell_comb \LessThan1~47 (
// Equation(s):
// \LessThan1~47_cout  = CARRY((\port_b~36_combout  & (\rdat1[23]~53_combout  & !\LessThan1~45_cout )) # (!\port_b~36_combout  & ((\rdat1[23]~53_combout ) # (!\LessThan1~45_cout ))))

	.dataa(port_b26),
	.datab(rdat1_23),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~45_cout ),
	.combout(),
	.cout(\LessThan1~47_cout ));
// synopsys translate_off
defparam \LessThan1~47 .lut_mask = 16'h004D;
defparam \LessThan1~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N16
cycloneive_lcell_comb \LessThan1~49 (
// Equation(s):
// \LessThan1~49_cout  = CARRY((\rdat1[24]~49_combout  & (\port_b~38_combout  & !\LessThan1~47_cout )) # (!\rdat1[24]~49_combout  & ((\port_b~38_combout ) # (!\LessThan1~47_cout ))))

	.dataa(rdat1_24),
	.datab(port_b28),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~47_cout ),
	.combout(),
	.cout(\LessThan1~49_cout ));
// synopsys translate_off
defparam \LessThan1~49 .lut_mask = 16'h004D;
defparam \LessThan1~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N18
cycloneive_lcell_comb \LessThan1~51 (
// Equation(s):
// \LessThan1~51_cout  = CARRY((\rdat1[25]~47_combout  & ((!\LessThan1~49_cout ) # (!\port_b~40_combout ))) # (!\rdat1[25]~47_combout  & (!\port_b~40_combout  & !\LessThan1~49_cout )))

	.dataa(rdat1_25),
	.datab(port_b30),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~49_cout ),
	.combout(),
	.cout(\LessThan1~51_cout ));
// synopsys translate_off
defparam \LessThan1~51 .lut_mask = 16'h002B;
defparam \LessThan1~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N20
cycloneive_lcell_comb \LessThan1~53 (
// Equation(s):
// \LessThan1~53_cout  = CARRY((\port_b~42_combout  & ((!\LessThan1~51_cout ) # (!\rdat1[26]~43_combout ))) # (!\port_b~42_combout  & (!\rdat1[26]~43_combout  & !\LessThan1~51_cout )))

	.dataa(port_b32),
	.datab(rdat1_26),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~51_cout ),
	.combout(),
	.cout(\LessThan1~53_cout ));
// synopsys translate_off
defparam \LessThan1~53 .lut_mask = 16'h002B;
defparam \LessThan1~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N22
cycloneive_lcell_comb \LessThan1~55 (
// Equation(s):
// \LessThan1~55_cout  = CARRY((\rdat1[27]~45_combout  & ((!\LessThan1~53_cout ) # (!\port_b~52_combout ))) # (!\rdat1[27]~45_combout  & (!\port_b~52_combout  & !\LessThan1~53_cout )))

	.dataa(rdat1_27),
	.datab(port_b42),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~53_cout ),
	.combout(),
	.cout(\LessThan1~55_cout ));
// synopsys translate_off
defparam \LessThan1~55 .lut_mask = 16'h002B;
defparam \LessThan1~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N24
cycloneive_lcell_comb \LessThan1~57 (
// Equation(s):
// \LessThan1~57_cout  = CARRY((\port_b~54_combout  & ((!\LessThan1~55_cout ) # (!\rdat1[28]~41_combout ))) # (!\port_b~54_combout  & (!\rdat1[28]~41_combout  & !\LessThan1~55_cout )))

	.dataa(port_b44),
	.datab(rdat1_28),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~55_cout ),
	.combout(),
	.cout(\LessThan1~57_cout ));
// synopsys translate_off
defparam \LessThan1~57 .lut_mask = 16'h002B;
defparam \LessThan1~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N26
cycloneive_lcell_comb \LessThan1~59 (
// Equation(s):
// \LessThan1~59_cout  = CARRY((\port_b~56_combout  & (\rdat1[29]~37_combout  & !\LessThan1~57_cout )) # (!\port_b~56_combout  & ((\rdat1[29]~37_combout ) # (!\LessThan1~57_cout ))))

	.dataa(port_b46),
	.datab(rdat1_29),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~57_cout ),
	.combout(),
	.cout(\LessThan1~59_cout ));
// synopsys translate_off
defparam \LessThan1~59 .lut_mask = 16'h004D;
defparam \LessThan1~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N28
cycloneive_lcell_comb \LessThan1~61 (
// Equation(s):
// \LessThan1~61_cout  = CARRY((\port_b~58_combout  & ((!\LessThan1~59_cout ) # (!\rdat1[30]~39_combout ))) # (!\port_b~58_combout  & (!\rdat1[30]~39_combout  & !\LessThan1~59_cout )))

	.dataa(port_b48),
	.datab(rdat1_30),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~59_cout ),
	.combout(),
	.cout(\LessThan1~61_cout ));
// synopsys translate_off
defparam \LessThan1~61 .lut_mask = 16'h002B;
defparam \LessThan1~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N30
cycloneive_lcell_comb \LessThan1~62 (
// Equation(s):
// \LessThan1~62_combout  = (\rdat1[31]~35_combout  & (\LessThan1~61_cout  & \port_b~20_combout )) # (!\rdat1[31]~35_combout  & ((\LessThan1~61_cout ) # (\port_b~20_combout )))

	.dataa(rdat1_311),
	.datab(gnd),
	.datac(gnd),
	.datad(port_b10),
	.cin(\LessThan1~61_cout ),
	.combout(\LessThan1~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan1~62 .lut_mask = 16'hF550;
defparam \LessThan1~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N16
cycloneive_lcell_comb \myif.out[0]~294 (
// Equation(s):
// \myif.out[0]~294_combout  = (!idex_ifaluop_o_2 & ((idex_ifaluop_o_0 & ((\LessThan1~62_combout ))) # (!idex_ifaluop_o_0 & (\LessThan0~62_combout ))))

	.dataa(\LessThan0~62_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(idex_ifaluop_o_0),
	.datad(\LessThan1~62_combout ),
	.cin(gnd),
	.combout(\myif.out[0]~294_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[0]~294 .lut_mask = 16'h3202;
defparam \myif.out[0]~294 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N6
cycloneive_lcell_comb \myif.out[0]~295 (
// Equation(s):
// \myif.out[0]~295_combout  = (idex_ifaluop_o_3 & (idex_ifaluop_o_1 & ((\myif.out[0]~294_combout )))) # (!idex_ifaluop_o_3 & (!idex_ifaluop_o_1 & (\myif.out[0]~236_combout )))

	.dataa(idex_ifaluop_o_3),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[0]~236_combout ),
	.datad(\myif.out[0]~294_combout ),
	.cin(gnd),
	.combout(\myif.out[0]~295_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[0]~295 .lut_mask = 16'h9810;
defparam \myif.out[0]~295 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N12
cycloneive_lcell_comb \Equal10~8 (
// Equation(s):
// \Equal10~8_combout  = (myifout_22) # ((myifout_20) # ((myifnegative) # (myifout_21)))

	.dataa(myifout_22),
	.datab(myifout_20),
	.datac(myifnegative),
	.datad(myifout_21),
	.cin(gnd),
	.combout(\Equal10~8_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~8 .lut_mask = 16'hFFFE;
defparam \Equal10~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N6
cycloneive_lcell_comb \Equal10~9 (
// Equation(s):
// \Equal10~9_combout  = (idex_ifaluop_o_3) # ((!myifout_30 & (!myifout_19 & !\Equal10~8_combout )))

	.dataa(myifout_30),
	.datab(idex_ifaluop_o_3),
	.datac(myifout_19),
	.datad(\Equal10~8_combout ),
	.cin(gnd),
	.combout(\Equal10~9_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~9 .lut_mask = 16'hCCCD;
defparam \Equal10~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N8
cycloneive_lcell_comb \Equal10~4 (
// Equation(s):
// \Equal10~4_combout  = (idex_ifaluop_o_3) # ((!myifout_15 & (!myifout_12 & !myifout_14)))

	.dataa(myifout_15),
	.datab(idex_ifaluop_o_3),
	.datac(myifout_12),
	.datad(myifout_14),
	.cin(gnd),
	.combout(\Equal10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~4 .lut_mask = 16'hCCCD;
defparam \Equal10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N6
cycloneive_lcell_comb \Equal10~3 (
// Equation(s):
// \Equal10~3_combout  = (idex_ifaluop_o_3) # ((!myifout_8 & (!myifout_13 & !myifout_9)))

	.dataa(myifout_8),
	.datab(idex_ifaluop_o_3),
	.datac(myifout_13),
	.datad(myifout_9),
	.cin(gnd),
	.combout(\Equal10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~3 .lut_mask = 16'hCCCD;
defparam \Equal10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N8
cycloneive_lcell_comb \Equal10~6 (
// Equation(s):
// \Equal10~6_combout  = (idex_ifaluop_o_3) # ((!myifout_18 & (!myifout_16 & !myifout_17)))

	.dataa(idex_ifaluop_o_3),
	.datab(myifout_18),
	.datac(myifout_16),
	.datad(myifout_17),
	.cin(gnd),
	.combout(\Equal10~6_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~6 .lut_mask = 16'hAAAB;
defparam \Equal10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N18
cycloneive_lcell_comb \Equal10~5 (
// Equation(s):
// \Equal10~5_combout  = (idex_ifaluop_o_3) # ((!myifout_11 & (!myifout_10 & !myifout_23)))

	.dataa(idex_ifaluop_o_3),
	.datab(myifout_11),
	.datac(myifout_10),
	.datad(myifout_23),
	.cin(gnd),
	.combout(\Equal10~5_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~5 .lut_mask = 16'hAAAB;
defparam \Equal10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N26
cycloneive_lcell_comb \Equal10~7 (
// Equation(s):
// \Equal10~7_combout  = (\Equal10~4_combout  & (\Equal10~3_combout  & (\Equal10~6_combout  & \Equal10~5_combout )))

	.dataa(\Equal10~4_combout ),
	.datab(\Equal10~3_combout ),
	.datac(\Equal10~6_combout ),
	.datad(\Equal10~5_combout ),
	.cin(gnd),
	.combout(\Equal10~7_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~7 .lut_mask = 16'h8000;
defparam \Equal10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N10
cycloneive_lcell_comb \Equal10~1 (
// Equation(s):
// \Equal10~1_combout  = (!myifout_24 & (!myifout_27 & (!myifout_26 & !myifout_25)))

	.dataa(myifout_24),
	.datab(myifout_27),
	.datac(myifout_26),
	.datad(myifout_25),
	.cin(gnd),
	.combout(\Equal10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~1 .lut_mask = 16'h0001;
defparam \Equal10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N14
cycloneive_lcell_comb \Equal10~0 (
// Equation(s):
// \Equal10~0_combout  = (!myifout_6 & !myifout_4)

	.dataa(gnd),
	.datab(gnd),
	.datac(myifout_6),
	.datad(myifout_4),
	.cin(gnd),
	.combout(\Equal10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~0 .lut_mask = 16'h000F;
defparam \Equal10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N18
cycloneive_lcell_comb \Equal10~2 (
// Equation(s):
// \Equal10~2_combout  = (!myifout_7 & (!myifout_5 & (\Equal10~1_combout  & \Equal10~0_combout )))

	.dataa(myifout_7),
	.datab(myifout_5),
	.datac(\Equal10~1_combout ),
	.datad(\Equal10~0_combout ),
	.cin(gnd),
	.combout(\Equal10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~2 .lut_mask = 16'h1000;
defparam \Equal10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N22
cycloneive_lcell_comb \myif.out[3]~246 (
// Equation(s):
// \myif.out[3]~246_combout  = (idex_ifaluop_o_2 & idex_ifaluop_o_1)

	.dataa(gnd),
	.datab(gnd),
	.datac(idex_ifaluop_o_2),
	.datad(idex_ifaluop_o_1),
	.cin(gnd),
	.combout(\myif.out[3]~246_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[3]~246 .lut_mask = 16'hF000;
defparam \myif.out[3]~246 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N24
cycloneive_lcell_comb \myif.out[28]~247 (
// Equation(s):
// \myif.out[28]~247_combout  = (\myif.out[5]~245_combout  & (\myif.out[3]~246_combout  & (\rdat1[28]~41_combout  $ (\port_b~54_combout ))))

	.dataa(\myif.out[5]~245_combout ),
	.datab(\myif.out[3]~246_combout ),
	.datac(rdat1_28),
	.datad(port_b44),
	.cin(gnd),
	.combout(\myif.out[28]~247_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[28]~247 .lut_mask = 16'h0880;
defparam \myif.out[28]~247 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N22
cycloneive_lcell_comb \out~75 (
// Equation(s):
// \out~75_combout  = (\port_b~53_combout ) # ((\rdat1[28]~41_combout ) # ((\port_b~0_combout  & fuifrtReplace_28)))

	.dataa(port_b),
	.datab(port_b43),
	.datac(rdat1_28),
	.datad(fuifrtReplace_28),
	.cin(gnd),
	.combout(\out~75_combout ),
	.cout());
// synopsys translate_off
defparam \out~75 .lut_mask = 16'hFEFC;
defparam \out~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N28
cycloneive_lcell_comb \myif.out[28]~249 (
// Equation(s):
// \myif.out[28]~249_combout  = (\myif.out[13]~23_combout  & ((idex_ifaluop_o_2 & ((\out~75_combout ))) # (!idex_ifaluop_o_2 & (\ShiftRight0~95_combout )))) # (!\myif.out[13]~23_combout  & (((idex_ifaluop_o_2))))

	.dataa(\ShiftRight0~95_combout ),
	.datab(\myif.out[13]~23_combout ),
	.datac(idex_ifaluop_o_2),
	.datad(\out~75_combout ),
	.cin(gnd),
	.combout(\myif.out[28]~249_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[28]~249 .lut_mask = 16'hF838;
defparam \myif.out[28]~249 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N16
cycloneive_lcell_comb \myif.out[28]~292 (
// Equation(s):
// \myif.out[28]~292_combout  = (idex_ifaluop_o_1 & ((\myif.out[28]~249_combout  & ((!\out~75_combout ))) # (!\myif.out[28]~249_combout  & (\Add1~56_combout )))) # (!idex_ifaluop_o_1 & (((\myif.out[28]~249_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(\Add1~56_combout ),
	.datac(\out~75_combout ),
	.datad(\myif.out[28]~249_combout ),
	.cin(gnd),
	.combout(\myif.out[28]~292_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[28]~292 .lut_mask = 16'h5F88;
defparam \myif.out[28]~292 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N30
cycloneive_lcell_comb \myif.out[28]~293 (
// Equation(s):
// \myif.out[28]~293_combout  = (\myif.out[28]~247_combout ) # ((!idex_ifaluop_o_3 & (idex_ifaluop_o_0 & \myif.out[28]~292_combout )))

	.dataa(\myif.out[28]~247_combout ),
	.datab(idex_ifaluop_o_3),
	.datac(idex_ifaluop_o_0),
	.datad(\myif.out[28]~292_combout ),
	.cin(gnd),
	.combout(\myif.out[28]~293_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[28]~293 .lut_mask = 16'hBAAA;
defparam \myif.out[28]~293 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N8
cycloneive_lcell_comb \out~74 (
// Equation(s):
// \out~74_combout  = (\rdat1[28]~41_combout  & ((\port_b~53_combout ) # ((fuifrtReplace_28 & \port_b~0_combout ))))

	.dataa(fuifrtReplace_28),
	.datab(port_b),
	.datac(rdat1_28),
	.datad(port_b43),
	.cin(gnd),
	.combout(\out~74_combout ),
	.cout());
// synopsys translate_off
defparam \out~74 .lut_mask = 16'hF080;
defparam \out~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N2
cycloneive_lcell_comb \myif.out[3]~240 (
// Equation(s):
// \myif.out[3]~240_combout  = (idex_ifaluop_o_1) # ((\port_b~17_combout  & !idex_ifaluop_o_2))

	.dataa(idex_ifaluop_o_1),
	.datab(port_b8),
	.datac(idex_ifaluop_o_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\myif.out[3]~240_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[3]~240 .lut_mask = 16'hAEAE;
defparam \myif.out[3]~240 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N30
cycloneive_lcell_comb \myif.out[3]~241 (
// Equation(s):
// \myif.out[3]~241_combout  = (\port_b~14_combout ) # ((\port_b~4_combout  & !\port_b~10_combout ))

	.dataa(port_b2),
	.datab(port_b6),
	.datac(port_b7),
	.datad(gnd),
	.cin(gnd),
	.combout(\myif.out[3]~241_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[3]~241 .lut_mask = 16'hF2F2;
defparam \myif.out[3]~241 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N12
cycloneive_lcell_comb \myif.out[28]~242 (
// Equation(s):
// \myif.out[28]~242_combout  = (\ShiftRight0~112_combout  & (((!\myif.out[3]~241_combout  & \ShiftLeft0~104_combout )))) # (!\ShiftRight0~112_combout  & ((\ShiftLeft0~36_combout ) # ((\myif.out[3]~241_combout ))))

	.dataa(\ShiftRight0~112_combout ),
	.datab(\ShiftLeft0~36_combout ),
	.datac(\myif.out[3]~241_combout ),
	.datad(\ShiftLeft0~104_combout ),
	.cin(gnd),
	.combout(\myif.out[28]~242_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[28]~242 .lut_mask = 16'h5E54;
defparam \myif.out[28]~242 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N2
cycloneive_lcell_comb \myif.out[28]~243 (
// Equation(s):
// \myif.out[28]~243_combout  = (\myif.out[3]~241_combout  & ((\myif.out[28]~242_combout  & (\ShiftLeft0~108_combout )) # (!\myif.out[28]~242_combout  & ((\ShiftLeft0~50_combout ))))) # (!\myif.out[3]~241_combout  & (((\myif.out[28]~242_combout ))))

	.dataa(\ShiftLeft0~108_combout ),
	.datab(\ShiftLeft0~50_combout ),
	.datac(\myif.out[3]~241_combout ),
	.datad(\myif.out[28]~242_combout ),
	.cin(gnd),
	.combout(\myif.out[28]~243_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[28]~243 .lut_mask = 16'hAFC0;
defparam \myif.out[28]~243 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N0
cycloneive_lcell_comb \myif.out[28]~244 (
// Equation(s):
// \myif.out[28]~244_combout  = (\myif.out[1]~8_combout  & (((!\myif.out[3]~240_combout  & \myif.out[28]~243_combout )))) # (!\myif.out[1]~8_combout  & ((\out~74_combout ) # ((\myif.out[3]~240_combout ))))

	.dataa(\myif.out[1]~8_combout ),
	.datab(\out~74_combout ),
	.datac(\myif.out[3]~240_combout ),
	.datad(\myif.out[28]~243_combout ),
	.cin(gnd),
	.combout(\myif.out[28]~244_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[28]~244 .lut_mask = 16'h5E54;
defparam \myif.out[28]~244 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N14
cycloneive_lcell_comb \myif.out[28]~248 (
// Equation(s):
// \myif.out[28]~248_combout  = (\myif.out[28]~247_combout ) # ((\myif.out[3]~240_combout  & \ShiftLeft0~97_combout ))

	.dataa(gnd),
	.datab(\myif.out[3]~240_combout ),
	.datac(\ShiftLeft0~97_combout ),
	.datad(\myif.out[28]~247_combout ),
	.cin(gnd),
	.combout(\myif.out[28]~248_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[28]~248 .lut_mask = 16'hFFC0;
defparam \myif.out[28]~248 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N22
cycloneive_lcell_comb \myif.out[28]~251 (
// Equation(s):
// \myif.out[28]~251_combout  = (\myif.out[3]~240_combout  & (!\myif.out[28]~247_combout  & !\Add0~56_combout ))

	.dataa(gnd),
	.datab(\myif.out[3]~240_combout ),
	.datac(\myif.out[28]~247_combout ),
	.datad(\Add0~56_combout ),
	.cin(gnd),
	.combout(\myif.out[28]~251_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[28]~251 .lut_mask = 16'h000C;
defparam \myif.out[28]~251 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N8
cycloneive_lcell_comb \myif.out[5]~245 (
// Equation(s):
// \myif.out[5]~245_combout  = (!idex_ifaluop_o_3 & !idex_ifaluop_o_0)

	.dataa(gnd),
	.datab(gnd),
	.datac(idex_ifaluop_o_3),
	.datad(idex_ifaluop_o_0),
	.cin(gnd),
	.combout(\myif.out[5]~245_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[5]~245 .lut_mask = 16'h000F;
defparam \myif.out[5]~245 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N28
cycloneive_lcell_comb \myif.out[28]~250 (
// Equation(s):
// \myif.out[28]~250_combout  = (!\myif.out[3]~246_combout  & (\myif.out[5]~245_combout  & ((!\ShiftLeft0~11_combout ) # (!\myif.out[1]~8_combout ))))

	.dataa(\myif.out[3]~246_combout ),
	.datab(\myif.out[1]~8_combout ),
	.datac(\myif.out[5]~245_combout ),
	.datad(\ShiftLeft0~11_combout ),
	.cin(gnd),
	.combout(\myif.out[28]~250_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[28]~250 .lut_mask = 16'h1050;
defparam \myif.out[28]~250 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N18
cycloneive_lcell_comb \myif.out[28]~290 (
// Equation(s):
// \myif.out[28]~290_combout  = (\myif.out[28]~250_combout  & (((!idex_ifaluop_o_1 & !idex_ifaluop_o_2)) # (!\myif.out[28]~251_combout )))

	.dataa(idex_ifaluop_o_1),
	.datab(idex_ifaluop_o_2),
	.datac(\myif.out[28]~251_combout ),
	.datad(\myif.out[28]~250_combout ),
	.cin(gnd),
	.combout(\myif.out[28]~290_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[28]~290 .lut_mask = 16'h1F00;
defparam \myif.out[28]~290 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N28
cycloneive_lcell_comb \myif.out[29]~260 (
// Equation(s):
// \myif.out[29]~260_combout  = (\port_b~55_combout ) # ((\rdat1[29]~37_combout ) # ((fuifrtReplace_29 & \port_b~0_combout )))

	.dataa(fuifrtReplace_29),
	.datab(port_b),
	.datac(port_b45),
	.datad(rdat1_29),
	.cin(gnd),
	.combout(\myif.out[29]~260_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[29]~260 .lut_mask = 16'hFFF8;
defparam \myif.out[29]~260 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N30
cycloneive_lcell_comb \myif.out[29]~261 (
// Equation(s):
// \myif.out[29]~261_combout  = (idex_ifaluop_o_2 & (((\myif.out[29]~260_combout ) # (!\myif.out[13]~23_combout )))) # (!idex_ifaluop_o_2 & (\ShiftRight0~91_combout  & ((\myif.out[13]~23_combout ))))

	.dataa(\ShiftRight0~91_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\myif.out[29]~260_combout ),
	.datad(\myif.out[13]~23_combout ),
	.cin(gnd),
	.combout(\myif.out[29]~261_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[29]~261 .lut_mask = 16'hE2CC;
defparam \myif.out[29]~261 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N30
cycloneive_lcell_comb \myif.out[29]~253 (
// Equation(s):
// \myif.out[29]~253_combout  = (\myif.out[5]~245_combout  & (\myif.out[3]~246_combout  & (\port_b~56_combout  $ (\rdat1[29]~37_combout ))))

	.dataa(\myif.out[5]~245_combout ),
	.datab(\myif.out[3]~246_combout ),
	.datac(port_b46),
	.datad(rdat1_29),
	.cin(gnd),
	.combout(\myif.out[29]~253_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[29]~253 .lut_mask = 16'h0880;
defparam \myif.out[29]~253 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N0
cycloneive_lcell_comb \myif.out[29]~262 (
// Equation(s):
// \myif.out[29]~262_combout  = (\myif.out[29]~253_combout  & ((!\myif.out[29]~261_combout ))) # (!\myif.out[29]~253_combout  & (\myif.out[29]~260_combout  & \myif.out[29]~261_combout ))

	.dataa(\myif.out[29]~260_combout ),
	.datab(\myif.out[29]~253_combout ),
	.datac(\myif.out[29]~261_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\myif.out[29]~262_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[29]~262 .lut_mask = 16'h2C2C;
defparam \myif.out[29]~262 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N6
cycloneive_lcell_comb \myif.out[29]~263 (
// Equation(s):
// \myif.out[29]~263_combout  = (\myif.out[29]~261_combout  & (((!\myif.out[29]~262_combout )) # (!idex_ifaluop_o_1))) # (!\myif.out[29]~261_combout  & ((\myif.out[29]~262_combout ) # ((idex_ifaluop_o_1 & \Add1~58_combout ))))

	.dataa(\myif.out[29]~261_combout ),
	.datab(idex_ifaluop_o_1),
	.datac(\Add1~58_combout ),
	.datad(\myif.out[29]~262_combout ),
	.cin(gnd),
	.combout(\myif.out[29]~263_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[29]~263 .lut_mask = 16'h77EA;
defparam \myif.out[29]~263 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N8
cycloneive_lcell_comb \myif.out[29]~259 (
// Equation(s):
// \myif.out[29]~259_combout  = (\myif.out[29]~253_combout ) # ((!idex_ifaluop_o_3 & idex_ifaluop_o_0))

	.dataa(gnd),
	.datab(idex_ifaluop_o_3),
	.datac(\myif.out[29]~253_combout ),
	.datad(idex_ifaluop_o_0),
	.cin(gnd),
	.combout(\myif.out[29]~259_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[29]~259 .lut_mask = 16'hF3F0;
defparam \myif.out[29]~259 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N26
cycloneive_lcell_comb \myif.out[29]~254 (
// Equation(s):
// \myif.out[29]~254_combout  = (\myif.out[3]~240_combout  & (((\Add0~58_combout )))) # (!\myif.out[3]~240_combout  & (\port_b~56_combout  & (\rdat1[29]~37_combout )))

	.dataa(port_b46),
	.datab(\myif.out[3]~240_combout ),
	.datac(rdat1_29),
	.datad(\Add0~58_combout ),
	.cin(gnd),
	.combout(\myif.out[29]~254_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[29]~254 .lut_mask = 16'hEC20;
defparam \myif.out[29]~254 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N12
cycloneive_lcell_comb \ShiftLeft0~107 (
// Equation(s):
// \ShiftLeft0~107_combout  = (\port_b~7_combout  & (\rdat1[28]~41_combout )) # (!\port_b~7_combout  & ((\rdat1[29]~37_combout )))

	.dataa(gnd),
	.datab(port_b4),
	.datac(rdat1_28),
	.datad(rdat1_29),
	.cin(gnd),
	.combout(\ShiftLeft0~107_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~107 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N24
cycloneive_lcell_comb \myif.out[29]~255 (
// Equation(s):
// \myif.out[29]~255_combout  = (\ShiftRight0~112_combout  & (!\myif.out[3]~241_combout  & (\ShiftLeft0~107_combout ))) # (!\ShiftRight0~112_combout  & ((\myif.out[3]~241_combout ) # ((\ShiftLeft0~65_combout ))))

	.dataa(\ShiftRight0~112_combout ),
	.datab(\myif.out[3]~241_combout ),
	.datac(\ShiftLeft0~107_combout ),
	.datad(\ShiftLeft0~65_combout ),
	.cin(gnd),
	.combout(\myif.out[29]~255_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[29]~255 .lut_mask = 16'h7564;
defparam \myif.out[29]~255 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N10
cycloneive_lcell_comb \myif.out[29]~256 (
// Equation(s):
// \myif.out[29]~256_combout  = (\myif.out[3]~241_combout  & ((\myif.out[29]~255_combout  & ((\ShiftLeft0~106_combout ))) # (!\myif.out[29]~255_combout  & (\ShiftLeft0~80_combout )))) # (!\myif.out[3]~241_combout  & (((\myif.out[29]~255_combout ))))

	.dataa(\ShiftLeft0~80_combout ),
	.datab(\myif.out[3]~241_combout ),
	.datac(\ShiftLeft0~106_combout ),
	.datad(\myif.out[29]~255_combout ),
	.cin(gnd),
	.combout(\myif.out[29]~256_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[29]~256 .lut_mask = 16'hF388;
defparam \myif.out[29]~256 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N12
cycloneive_lcell_comb \myif.out[29]~257 (
// Equation(s):
// \myif.out[29]~257_combout  = (\myif.out[3]~240_combout  & (\ShiftLeft0~91_combout )) # (!\myif.out[3]~240_combout  & ((\myif.out[29]~256_combout )))

	.dataa(gnd),
	.datab(\myif.out[3]~240_combout ),
	.datac(\ShiftLeft0~91_combout ),
	.datad(\myif.out[29]~256_combout ),
	.cin(gnd),
	.combout(\myif.out[29]~257_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[29]~257 .lut_mask = 16'hF3C0;
defparam \myif.out[29]~257 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N18
cycloneive_lcell_comb \myif.out[29]~258 (
// Equation(s):
// \myif.out[29]~258_combout  = (\myif.out[29]~253_combout ) # ((\myif.out[1]~8_combout  & ((\myif.out[29]~257_combout ))) # (!\myif.out[1]~8_combout  & (\myif.out[29]~254_combout )))

	.dataa(\myif.out[29]~254_combout ),
	.datab(\myif.out[1]~8_combout ),
	.datac(\myif.out[29]~253_combout ),
	.datad(\myif.out[29]~257_combout ),
	.cin(gnd),
	.combout(\myif.out[29]~258_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[29]~258 .lut_mask = 16'hFEF2;
defparam \myif.out[29]~258 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N2
cycloneive_lcell_comb \myif.out[3]~273 (
// Equation(s):
// \myif.out[3]~273_combout  = (idex_ifaluop_o_1 & (idex_ifaluop_o_2 & (!idex_ifaluop_o_3 & idex_ifaluop_o_0)))

	.dataa(idex_ifaluop_o_1),
	.datab(idex_ifaluop_o_2),
	.datac(idex_ifaluop_o_3),
	.datad(idex_ifaluop_o_0),
	.cin(gnd),
	.combout(\myif.out[3]~273_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[3]~273 .lut_mask = 16'h0800;
defparam \myif.out[3]~273 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N26
cycloneive_lcell_comb \out~76 (
// Equation(s):
// \out~76_combout  = (\port_b~9_combout ) # ((\rdat1[2]~5_combout ) # ((\port_b~0_combout  & fuifrtReplace_2)))

	.dataa(port_b5),
	.datab(port_b),
	.datac(fuifrtReplace_2),
	.datad(rdat1_2),
	.cin(gnd),
	.combout(\out~76_combout ),
	.cout());
// synopsys translate_off
defparam \out~76 .lut_mask = 16'hFFEA;
defparam \out~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N12
cycloneive_lcell_comb \myif.out[2]~265 (
// Equation(s):
// \myif.out[2]~265_combout  = (!\port_b~0_combout ) # (!fuifrtReplace_2)

	.dataa(gnd),
	.datab(gnd),
	.datac(fuifrtReplace_2),
	.datad(port_b),
	.cin(gnd),
	.combout(\myif.out[2]~265_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[2]~265 .lut_mask = 16'h0FFF;
defparam \myif.out[2]~265 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N22
cycloneive_lcell_comb \myif.out[2]~266 (
// Equation(s):
// \myif.out[2]~266_combout  = (\rdat1[2]~5_combout  $ (((\port_b~9_combout ) # (!\myif.out[2]~265_combout )))) # (!idex_ifaluop_o_1)

	.dataa(port_b5),
	.datab(idex_ifaluop_o_1),
	.datac(rdat1_2),
	.datad(\myif.out[2]~265_combout ),
	.cin(gnd),
	.combout(\myif.out[2]~266_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[2]~266 .lut_mask = 16'h7B3F;
defparam \myif.out[2]~266 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N22
cycloneive_lcell_comb \myif.out[2]~267 (
// Equation(s):
// \myif.out[2]~267_combout  = (idex_ifaluop_o_2 & ((\port_b~9_combout ) # ((\port_b~0_combout  & fuifrtReplace_2))))

	.dataa(port_b),
	.datab(fuifrtReplace_2),
	.datac(port_b5),
	.datad(idex_ifaluop_o_2),
	.cin(gnd),
	.combout(\myif.out[2]~267_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[2]~267 .lut_mask = 16'hF800;
defparam \myif.out[2]~267 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N0
cycloneive_lcell_comb \myif.out[2]~268 (
// Equation(s):
// \myif.out[2]~268_combout  = (idex_ifaluop_o_1 & (\Add0~4_combout  & ((!\myif.out[2]~267_combout ) # (!\rdat1[2]~5_combout )))) # (!idex_ifaluop_o_1 & (\rdat1[2]~5_combout  & ((\myif.out[2]~267_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(rdat1_2),
	.datac(\Add0~4_combout ),
	.datad(\myif.out[2]~267_combout ),
	.cin(gnd),
	.combout(\myif.out[2]~268_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[2]~268 .lut_mask = 16'h64A0;
defparam \myif.out[2]~268 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N22
cycloneive_lcell_comb \myif.out[2]~269 (
// Equation(s):
// \myif.out[2]~269_combout  = (\ShiftLeft0~103_combout  & ((idex_ifaluop_o_2 & ((\myif.out[2]~268_combout ))) # (!idex_ifaluop_o_2 & (\myif.out[2]~266_combout )))) # (!\ShiftLeft0~103_combout  & (((\myif.out[2]~268_combout ))))

	.dataa(\ShiftLeft0~103_combout ),
	.datab(idex_ifaluop_o_2),
	.datac(\myif.out[2]~266_combout ),
	.datad(\myif.out[2]~268_combout ),
	.cin(gnd),
	.combout(\myif.out[2]~269_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[2]~269 .lut_mask = 16'hFD20;
defparam \myif.out[2]~269 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N4
cycloneive_lcell_comb \myif.out[2]~270 (
// Equation(s):
// \myif.out[2]~270_combout  = \rdat1[2]~5_combout  $ (((\port_b~9_combout ) # ((\port_b~0_combout  & fuifrtReplace_2))))

	.dataa(port_b5),
	.datab(port_b),
	.datac(fuifrtReplace_2),
	.datad(rdat1_2),
	.cin(gnd),
	.combout(\myif.out[2]~270_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[2]~270 .lut_mask = 16'h15EA;
defparam \myif.out[2]~270 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N14
cycloneive_lcell_comb \myif.out[2]~271 (
// Equation(s):
// \myif.out[2]~271_combout  = (idex_ifaluop_o_2 & (((\myif.out[2]~270_combout )) # (!idex_ifaluop_o_1))) # (!idex_ifaluop_o_2 & (((\myif.out[2]~268_combout ))))

	.dataa(idex_ifaluop_o_1),
	.datab(idex_ifaluop_o_2),
	.datac(\myif.out[2]~270_combout ),
	.datad(\myif.out[2]~268_combout ),
	.cin(gnd),
	.combout(\myif.out[2]~271_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[2]~271 .lut_mask = 16'hF7C4;
defparam \myif.out[2]~271 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N24
cycloneive_lcell_comb \myif.out[2]~272 (
// Equation(s):
// \myif.out[2]~272_combout  = (\myif.out[13]~23_combout  & (\myif.out[2]~269_combout )) # (!\myif.out[13]~23_combout  & ((\myif.out[2]~271_combout )))

	.dataa(\myif.out[2]~269_combout ),
	.datab(gnd),
	.datac(\myif.out[2]~271_combout ),
	.datad(\myif.out[13]~23_combout ),
	.cin(gnd),
	.combout(\myif.out[2]~272_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[2]~272 .lut_mask = 16'hAAF0;
defparam \myif.out[2]~272 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N22
cycloneive_lcell_comb \out~80 (
// Equation(s):
// \out~80_combout  = (\rdat1[3]~8_combout ) # ((\port_b~14_combout ) # ((\mem_data~12_combout  & always03)))

	.dataa(mem_data1),
	.datab(always0),
	.datac(rdat1_3),
	.datad(port_b7),
	.cin(gnd),
	.combout(\out~80_combout ),
	.cout());
// synopsys translate_off
defparam \out~80 .lut_mask = 16'hFFF8;
defparam \out~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N28
cycloneive_lcell_comb \ShiftRight0~99 (
// Equation(s):
// \ShiftRight0~99_combout  = (\port_b~10_combout  & ((\ShiftRight0~84_combout ) # ((\ShiftRight0~83_combout )))) # (!\port_b~10_combout  & (((\ShiftRight0~80_combout ))))

	.dataa(\ShiftRight0~84_combout ),
	.datab(port_b6),
	.datac(\ShiftRight0~83_combout ),
	.datad(\ShiftRight0~80_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~99_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~99 .lut_mask = 16'hFBC8;
defparam \ShiftRight0~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N10
cycloneive_lcell_comb \ShiftRight0~112 (
// Equation(s):
// \ShiftRight0~112_combout  = (!\port_b~9_combout  & (!\port_b~14_combout  & ((!fuifrtReplace_2) # (!\port_b~0_combout ))))

	.dataa(port_b),
	.datab(port_b5),
	.datac(fuifrtReplace_2),
	.datad(port_b7),
	.cin(gnd),
	.combout(\ShiftRight0~112_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~112 .lut_mask = 16'h0013;
defparam \ShiftRight0~112 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N12
cycloneive_lcell_comb \myif.out[3]~280 (
// Equation(s):
// \myif.out[3]~280_combout  = (\ShiftRight0~112_combout  & (\ShiftRight0~3_combout  & (!\myif.out[3]~241_combout ))) # (!\ShiftRight0~112_combout  & (((\myif.out[3]~241_combout ) # (\ShiftRight0~86_combout ))))

	.dataa(\ShiftRight0~3_combout ),
	.datab(\ShiftRight0~112_combout ),
	.datac(\myif.out[3]~241_combout ),
	.datad(\ShiftRight0~86_combout ),
	.cin(gnd),
	.combout(\myif.out[3]~280_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[3]~280 .lut_mask = 16'h3B38;
defparam \myif.out[3]~280 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N18
cycloneive_lcell_comb \myif.out[3]~281 (
// Equation(s):
// \myif.out[3]~281_combout  = (\myif.out[3]~241_combout  & ((\myif.out[3]~280_combout  & ((\ShiftRight0~99_combout ))) # (!\myif.out[3]~280_combout  & (\ShiftRight0~6_combout )))) # (!\myif.out[3]~241_combout  & (((\myif.out[3]~280_combout ))))

	.dataa(\myif.out[3]~241_combout ),
	.datab(\ShiftRight0~6_combout ),
	.datac(\ShiftRight0~99_combout ),
	.datad(\myif.out[3]~280_combout ),
	.cin(gnd),
	.combout(\myif.out[3]~281_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[3]~281 .lut_mask = 16'hF588;
defparam \myif.out[3]~281 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N8
cycloneive_lcell_comb \myif.out[3]~282 (
// Equation(s):
// \myif.out[3]~282_combout  = (\myif.out[3]~240_combout  & (((!\myif.out[1]~8_combout )))) # (!\myif.out[3]~240_combout  & ((\myif.out[1]~8_combout  & ((\myif.out[3]~281_combout ))) # (!\myif.out[1]~8_combout  & (\out~80_combout ))))

	.dataa(\out~80_combout ),
	.datab(\myif.out[3]~240_combout ),
	.datac(\myif.out[1]~8_combout ),
	.datad(\myif.out[3]~281_combout ),
	.cin(gnd),
	.combout(\myif.out[3]~282_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[3]~282 .lut_mask = 16'h3E0E;
defparam \myif.out[3]~282 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N10
cycloneive_lcell_comb \myif.out[5]~284 (
// Equation(s):
// \myif.out[5]~284_combout  = (!idex_ifaluop_o_3 & idex_ifaluop_o_0)

	.dataa(gnd),
	.datab(gnd),
	.datac(idex_ifaluop_o_3),
	.datad(idex_ifaluop_o_0),
	.cin(gnd),
	.combout(\myif.out[5]~284_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[5]~284 .lut_mask = 16'h0F00;
defparam \myif.out[5]~284 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N6
cycloneive_lcell_comb \ShiftRight0~59 (
// Equation(s):
// \ShiftRight0~59_combout  = (\port_b~7_combout  & ((\rdat1[5]~17_combout ))) # (!\port_b~7_combout  & (\rdat1[4]~7_combout ))

	.dataa(port_b4),
	.datab(gnd),
	.datac(rdat1_41),
	.datad(rdat1_5),
	.cin(gnd),
	.combout(\ShiftRight0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~59 .lut_mask = 16'hFA50;
defparam \ShiftRight0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N12
cycloneive_lcell_comb \ShiftRight0~107 (
// Equation(s):
// \ShiftRight0~107_combout  = (\port_b~7_combout  & (\rdat1[3]~9_combout )) # (!\port_b~7_combout  & ((\rdat1[2]~5_combout )))

	.dataa(rdat1_31),
	.datab(gnd),
	.datac(port_b4),
	.datad(rdat1_2),
	.cin(gnd),
	.combout(\ShiftRight0~107_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~107 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N28
cycloneive_lcell_comb \ShiftRight0~44 (
// Equation(s):
// \ShiftRight0~44_combout  = (\port_b~4_combout  & ((\ShiftRight0~42_combout ))) # (!\port_b~4_combout  & (\ShiftRight0~43_combout ))

	.dataa(gnd),
	.datab(port_b2),
	.datac(\ShiftRight0~43_combout ),
	.datad(\ShiftRight0~42_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~44_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~44 .lut_mask = 16'hFC30;
defparam \ShiftRight0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N4
cycloneive_lcell_comb \myif.out[2]~286 (
// Equation(s):
// \myif.out[2]~286_combout  = (\myif.out[3]~241_combout  & (((!\ShiftRight0~112_combout )))) # (!\myif.out[3]~241_combout  & ((\ShiftRight0~112_combout  & (\ShiftRight0~107_combout )) # (!\ShiftRight0~112_combout  & ((\ShiftRight0~44_combout )))))

	.dataa(\myif.out[3]~241_combout ),
	.datab(\ShiftRight0~107_combout ),
	.datac(\ShiftRight0~112_combout ),
	.datad(\ShiftRight0~44_combout ),
	.cin(gnd),
	.combout(\myif.out[2]~286_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[2]~286 .lut_mask = 16'h4F4A;
defparam \myif.out[2]~286 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N2
cycloneive_lcell_comb \myif.out[2]~287 (
// Equation(s):
// \myif.out[2]~287_combout  = (\myif.out[3]~241_combout  & ((\myif.out[2]~286_combout  & ((\ShiftRight0~97_combout ))) # (!\myif.out[2]~286_combout  & (\ShiftRight0~59_combout )))) # (!\myif.out[3]~241_combout  & (((\myif.out[2]~286_combout ))))

	.dataa(\myif.out[3]~241_combout ),
	.datab(\ShiftRight0~59_combout ),
	.datac(\myif.out[2]~286_combout ),
	.datad(\ShiftRight0~97_combout ),
	.cin(gnd),
	.combout(\myif.out[2]~287_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[2]~287 .lut_mask = 16'hF858;
defparam \myif.out[2]~287 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N28
cycloneive_lcell_comb \myif.out[2]~288 (
// Equation(s):
// \myif.out[2]~288_combout  = (\myif.out[3]~240_combout  & ((\ShiftRight0~103_combout ) # ((!\myif.out[1]~8_combout )))) # (!\myif.out[3]~240_combout  & (((\myif.out[1]~8_combout  & \myif.out[2]~287_combout ))))

	.dataa(\ShiftRight0~103_combout ),
	.datab(\myif.out[3]~240_combout ),
	.datac(\myif.out[1]~8_combout ),
	.datad(\myif.out[2]~287_combout ),
	.cin(gnd),
	.combout(\myif.out[2]~288_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[2]~288 .lut_mask = 16'hBC8C;
defparam \myif.out[2]~288 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N14
cycloneive_lcell_comb \Equal10~11 (
// Equation(s):
// \Equal10~11_combout  = (!myifout_32 & (((!myifout_210 & !myifout_3)) # (!myifout_31)))

	.dataa(myifout_32),
	.datab(myifout_210),
	.datac(myifout_31),
	.datad(myifout_3),
	.cin(gnd),
	.combout(\Equal10~11_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~11 .lut_mask = 16'h0515;
defparam \Equal10~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N8
cycloneive_lcell_comb \ShiftLeft0~109 (
// Equation(s):
// \ShiftLeft0~109_combout  = (\ShiftRight0~112_combout  & ((\port_b~4_combout  & (\ShiftLeft0~12_combout )) # (!\port_b~4_combout  & ((\ShiftLeft0~66_combout )))))

	.dataa(\ShiftRight0~112_combout ),
	.datab(port_b2),
	.datac(\ShiftLeft0~12_combout ),
	.datad(\ShiftLeft0~66_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~109_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~109 .lut_mask = 16'hA280;
defparam \ShiftLeft0~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N16
cycloneive_lcell_comb \myif.out[3]~276 (
// Equation(s):
// \myif.out[3]~276_combout  = (\myif.out[13]~23_combout  & ((idex_ifaluop_o_2) # (\ShiftLeft0~109_combout )))

	.dataa(gnd),
	.datab(idex_ifaluop_o_2),
	.datac(\ShiftLeft0~109_combout ),
	.datad(\myif.out[13]~23_combout ),
	.cin(gnd),
	.combout(\myif.out[3]~276_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[3]~276 .lut_mask = 16'hFC00;
defparam \myif.out[3]~276 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N26
cycloneive_lcell_comb \myif.out[3]~277 (
// Equation(s):
// \myif.out[3]~277_combout  = (\rdat1[3]~9_combout  & (\port_b~14_combout  & ((idex_ifaluop_o_2) # (\myif.out[3]~276_combout )))) # (!\rdat1[3]~9_combout  & (!\port_b~14_combout  & (idex_ifaluop_o_2 $ (\myif.out[3]~276_combout ))))

	.dataa(rdat1_31),
	.datab(idex_ifaluop_o_2),
	.datac(port_b7),
	.datad(\myif.out[3]~276_combout ),
	.cin(gnd),
	.combout(\myif.out[3]~277_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[3]~277 .lut_mask = 16'hA184;
defparam \myif.out[3]~277 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N0
cycloneive_lcell_comb \myif.out[3]~278 (
// Equation(s):
// \myif.out[3]~278_combout  = (\rdat1[3]~9_combout  & (!\port_b~14_combout  & (idex_ifaluop_o_2 $ (\myif.out[3]~276_combout )))) # (!\rdat1[3]~9_combout  & (\port_b~14_combout  & (idex_ifaluop_o_2 $ (\myif.out[3]~276_combout ))))

	.dataa(rdat1_31),
	.datab(idex_ifaluop_o_2),
	.datac(port_b7),
	.datad(\myif.out[3]~276_combout ),
	.cin(gnd),
	.combout(\myif.out[3]~278_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[3]~278 .lut_mask = 16'h1248;
defparam \myif.out[3]~278 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N14
cycloneive_lcell_comb \myif.out[3]~279 (
// Equation(s):
// \myif.out[3]~279_combout  = (idex_ifaluop_o_1 & ((\Add0~6_combout  & ((\myif.out[3]~278_combout ) # (!\myif.out[3]~277_combout ))) # (!\Add0~6_combout  & (!\myif.out[3]~277_combout  & \myif.out[3]~278_combout )))) # (!idex_ifaluop_o_1 & 
// ((\myif.out[3]~277_combout  $ (\myif.out[3]~278_combout ))))

	.dataa(\Add0~6_combout ),
	.datab(idex_ifaluop_o_1),
	.datac(\myif.out[3]~277_combout ),
	.datad(\myif.out[3]~278_combout ),
	.cin(gnd),
	.combout(\myif.out[3]~279_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[3]~279 .lut_mask = 16'h8F38;
defparam \myif.out[3]~279 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N20
cycloneive_lcell_comb \myif.out[3]~275 (
// Equation(s):
// \myif.out[3]~275_combout  = (\myif.out[3]~273_combout  & !\out~80_combout )

	.dataa(\myif.out[3]~273_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\out~80_combout ),
	.cin(gnd),
	.combout(\myif.out[3]~275_combout ),
	.cout());
// synopsys translate_off
defparam \myif.out[3]~275 .lut_mask = 16'h00AA;
defparam \myif.out[3]~275 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module control_unit (
	ifid_ifinstr_o_26,
	ifid_ifinstr_o_31,
	ifid_ifinstr_o_27,
	ifid_ifinstr_o_28,
	ifid_ifinstr_o_30,
	ifid_ifinstr_o_5,
	ifid_ifinstr_o_4,
	always0,
	ifid_ifinstr_o_29,
	ifid_ifinstr_o_1,
	ifid_ifinstr_o_3,
	ifid_ifinstr_o_2,
	cuifregWEN,
	Equal0,
	ifid_ifinstr_o_0,
	Equal3,
	Equal2,
	Equal10,
	Equal14,
	Equal21,
	Equal01,
	Equal5,
	cuifregWEN1,
	Equal1,
	devpor,
	devclrn,
	devoe);
input 	ifid_ifinstr_o_26;
input 	ifid_ifinstr_o_31;
input 	ifid_ifinstr_o_27;
input 	ifid_ifinstr_o_28;
input 	ifid_ifinstr_o_30;
input 	ifid_ifinstr_o_5;
input 	ifid_ifinstr_o_4;
output 	always0;
input 	ifid_ifinstr_o_29;
input 	ifid_ifinstr_o_1;
input 	ifid_ifinstr_o_3;
input 	ifid_ifinstr_o_2;
output 	cuifregWEN;
output 	Equal0;
input 	ifid_ifinstr_o_0;
output 	Equal3;
output 	Equal2;
output 	Equal10;
output 	Equal14;
output 	Equal21;
output 	Equal01;
output 	Equal5;
output 	cuifregWEN1;
output 	Equal1;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \cuif.regWEN~3_combout ;
wire \cuif.regWEN~4_combout ;
wire \cuif.regWEN~1_combout ;
wire \cuif.regWEN~2_combout ;


// Location: LCCOMB_X61_Y26_N20
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// always0 = (ifid_ifinstr_o_5 & !ifid_ifinstr_o_4)

	.dataa(gnd),
	.datab(gnd),
	.datac(ifid_ifinstr_o_5),
	.datad(ifid_ifinstr_o_4),
	.cin(gnd),
	.combout(always0),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'h00F0;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N24
cycloneive_lcell_comb \cuif.regWEN~0 (
// Equation(s):
// cuifregWEN = (!ifid_ifinstr_o_31 & ifid_ifinstr_o_29)

	.dataa(gnd),
	.datab(ifid_ifinstr_o_31),
	.datac(gnd),
	.datad(ifid_ifinstr_o_29),
	.cin(gnd),
	.combout(cuifregWEN),
	.cout());
// synopsys translate_off
defparam \cuif.regWEN~0 .lut_mask = 16'h3300;
defparam \cuif.regWEN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N28
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// Equal0 = (!ifid_ifinstr_o_31 & !ifid_ifinstr_o_30)

	.dataa(ifid_ifinstr_o_31),
	.datab(ifid_ifinstr_o_30),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal0),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h1111;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N4
cycloneive_lcell_comb \Equal3~0 (
// Equation(s):
// Equal3 = (!ifid_ifinstr_o_2 & (!ifid_ifinstr_o_5 & (!ifid_ifinstr_o_0 & !ifid_ifinstr_o_4)))

	.dataa(ifid_ifinstr_o_2),
	.datab(ifid_ifinstr_o_5),
	.datac(ifid_ifinstr_o_0),
	.datad(ifid_ifinstr_o_4),
	.cin(gnd),
	.combout(Equal3),
	.cout());
// synopsys translate_off
defparam \Equal3~0 .lut_mask = 16'h0001;
defparam \Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N8
cycloneive_lcell_comb \Equal2~0 (
// Equation(s):
// Equal2 = (!ifid_ifinstr_o_26 & (!ifid_ifinstr_o_27 & (!ifid_ifinstr_o_28 & !ifid_ifinstr_o_29)))

	.dataa(ifid_ifinstr_o_26),
	.datab(ifid_ifinstr_o_27),
	.datac(ifid_ifinstr_o_28),
	.datad(ifid_ifinstr_o_29),
	.cin(gnd),
	.combout(Equal2),
	.cout());
// synopsys translate_off
defparam \Equal2~0 .lut_mask = 16'h0001;
defparam \Equal2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N24
cycloneive_lcell_comb \Equal10~0 (
// Equation(s):
// Equal10 = (ifid_ifinstr_o_2 & (ifid_ifinstr_o_5 & (!ifid_ifinstr_o_3 & !ifid_ifinstr_o_4)))

	.dataa(ifid_ifinstr_o_2),
	.datab(ifid_ifinstr_o_5),
	.datac(ifid_ifinstr_o_3),
	.datad(ifid_ifinstr_o_4),
	.cin(gnd),
	.combout(Equal10),
	.cout());
// synopsys translate_off
defparam \Equal10~0 .lut_mask = 16'h0008;
defparam \Equal10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N26
cycloneive_lcell_comb \Equal14~0 (
// Equation(s):
// Equal14 = (ifid_ifinstr_o_3 & (always0 & (!ifid_ifinstr_o_2 & ifid_ifinstr_o_1)))

	.dataa(ifid_ifinstr_o_3),
	.datab(always0),
	.datac(ifid_ifinstr_o_2),
	.datad(ifid_ifinstr_o_1),
	.cin(gnd),
	.combout(Equal14),
	.cout());
// synopsys translate_off
defparam \Equal14~0 .lut_mask = 16'h0800;
defparam \Equal14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y27_N24
cycloneive_lcell_comb \Equal2~1 (
// Equation(s):
// Equal21 = (!ifid_ifinstr_o_30 & (Equal2 & !ifid_ifinstr_o_31))

	.dataa(ifid_ifinstr_o_30),
	.datab(Equal2),
	.datac(gnd),
	.datad(ifid_ifinstr_o_31),
	.cin(gnd),
	.combout(Equal21),
	.cout());
// synopsys translate_off
defparam \Equal2~1 .lut_mask = 16'h0044;
defparam \Equal2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N12
cycloneive_lcell_comb \Equal0~1 (
// Equation(s):
// Equal01 = (!ifid_ifinstr_o_28 & (!ifid_ifinstr_o_31 & (!ifid_ifinstr_o_30 & ifid_ifinstr_o_27)))

	.dataa(ifid_ifinstr_o_28),
	.datab(ifid_ifinstr_o_31),
	.datac(ifid_ifinstr_o_30),
	.datad(ifid_ifinstr_o_27),
	.cin(gnd),
	.combout(Equal01),
	.cout());
// synopsys translate_off
defparam \Equal0~1 .lut_mask = 16'h0100;
defparam \Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N0
cycloneive_lcell_comb \Equal5~0 (
// Equation(s):
// Equal5 = (!ifid_ifinstr_o_1 & ifid_ifinstr_o_3)

	.dataa(ifid_ifinstr_o_1),
	.datab(ifid_ifinstr_o_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(Equal5),
	.cout());
// synopsys translate_off
defparam \Equal5~0 .lut_mask = 16'h4444;
defparam \Equal5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N14
cycloneive_lcell_comb \cuif.regWEN~5 (
// Equation(s):
// cuifregWEN1 = (\cuif.regWEN~3_combout ) # ((\cuif.regWEN~2_combout ) # ((\cuif.regWEN~4_combout  & ifid_ifinstr_o_27)))

	.dataa(\cuif.regWEN~3_combout ),
	.datab(\cuif.regWEN~4_combout ),
	.datac(ifid_ifinstr_o_27),
	.datad(\cuif.regWEN~2_combout ),
	.cin(gnd),
	.combout(cuifregWEN1),
	.cout());
// synopsys translate_off
defparam \cuif.regWEN~5 .lut_mask = 16'hFFEA;
defparam \cuif.regWEN~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N0
cycloneive_lcell_comb \Equal1~0 (
// Equation(s):
// Equal1 = (Equal01 & (ifid_ifinstr_o_26 & !ifid_ifinstr_o_29))

	.dataa(Equal01),
	.datab(gnd),
	.datac(ifid_ifinstr_o_26),
	.datad(ifid_ifinstr_o_29),
	.cin(gnd),
	.combout(Equal1),
	.cout());
// synopsys translate_off
defparam \Equal1~0 .lut_mask = 16'h00A0;
defparam \Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N26
cycloneive_lcell_comb \cuif.regWEN~3 (
// Equation(s):
// \cuif.regWEN~3_combout  = (cuifregWEN) # ((!Equal0 & ((!ifid_ifinstr_o_26) # (!ifid_ifinstr_o_27))))

	.dataa(Equal0),
	.datab(cuifregWEN),
	.datac(ifid_ifinstr_o_27),
	.datad(ifid_ifinstr_o_26),
	.cin(gnd),
	.combout(\cuif.regWEN~3_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.regWEN~3 .lut_mask = 16'hCDDD;
defparam \cuif.regWEN~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N20
cycloneive_lcell_comb \cuif.regWEN~4 (
// Equation(s):
// \cuif.regWEN~4_combout  = (ifid_ifinstr_o_28 & (((!ifid_ifinstr_o_29 & ifid_ifinstr_o_26)) # (!ifid_ifinstr_o_30))) # (!ifid_ifinstr_o_28 & (!ifid_ifinstr_o_29 & ((ifid_ifinstr_o_26))))

	.dataa(ifid_ifinstr_o_28),
	.datab(ifid_ifinstr_o_29),
	.datac(ifid_ifinstr_o_30),
	.datad(ifid_ifinstr_o_26),
	.cin(gnd),
	.combout(\cuif.regWEN~4_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.regWEN~4 .lut_mask = 16'h3B0A;
defparam \cuif.regWEN~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N6
cycloneive_lcell_comb \cuif.regWEN~1 (
// Equation(s):
// \cuif.regWEN~1_combout  = (((ifid_ifinstr_o_26) # (ifid_ifinstr_o_1)) # (!Equal3)) # (!ifid_ifinstr_o_3)

	.dataa(ifid_ifinstr_o_3),
	.datab(Equal3),
	.datac(ifid_ifinstr_o_26),
	.datad(ifid_ifinstr_o_1),
	.cin(gnd),
	.combout(\cuif.regWEN~1_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.regWEN~1 .lut_mask = 16'hFFF7;
defparam \cuif.regWEN~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N28
cycloneive_lcell_comb \cuif.regWEN~2 (
// Equation(s):
// \cuif.regWEN~2_combout  = (!ifid_ifinstr_o_28 & ((ifid_ifinstr_o_30) # ((!ifid_ifinstr_o_27 & \cuif.regWEN~1_combout ))))

	.dataa(ifid_ifinstr_o_28),
	.datab(ifid_ifinstr_o_27),
	.datac(ifid_ifinstr_o_30),
	.datad(\cuif.regWEN~1_combout ),
	.cin(gnd),
	.combout(\cuif.regWEN~2_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.regWEN~2 .lut_mask = 16'h5150;
defparam \cuif.regWEN~2 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module ex_mem (
	exmem_ifout_o_1,
	exmem_ifdWEN_o,
	exmem_ifdREN_o,
	exmem_ifout_o_0,
	exmem_ifout_o_3,
	exmem_ifout_o_2,
	exmem_ifout_o_5,
	exmem_ifout_o_4,
	exmem_ifout_o_7,
	exmem_ifout_o_6,
	exmem_ifout_o_9,
	exmem_ifout_o_8,
	exmem_ifout_o_11,
	exmem_ifout_o_10,
	exmem_ifout_o_13,
	exmem_ifout_o_12,
	exmem_ifout_o_15,
	exmem_ifout_o_14,
	exmem_ifout_o_17,
	exmem_ifout_o_16,
	exmem_ifout_o_19,
	exmem_ifout_o_18,
	exmem_ifout_o_21,
	exmem_ifout_o_20,
	exmem_ifout_o_23,
	exmem_ifout_o_22,
	exmem_ifout_o_25,
	exmem_ifout_o_24,
	exmem_ifout_o_27,
	exmem_ifout_o_26,
	exmem_ifout_o_29,
	exmem_ifout_o_28,
	exmem_ifout_o_31,
	exmem_ifout_o_30,
	always1,
	always11,
	exmem_ifhalt_o,
	exmem_ifrdat2_o_0,
	always12,
	idex_ifrt_o_0,
	idex_ifrt_o_1,
	exmem_ifRegDest_o_1,
	exmem_ifrt_o_1,
	exmem_ifrd_o_1,
	exmem_ifRegDest_o_0,
	exmem_ifrt_o_0,
	exmem_ifrd_o_0,
	idex_ifrt_o_2,
	idex_ifrt_o_3,
	exmem_ifrt_o_3,
	exmem_ifrd_o_3,
	exmem_ifrt_o_2,
	exmem_ifrd_o_2,
	exmem_ifregWEN_o,
	idex_ifrt_o_4,
	exmem_ifrt_o_4,
	exmem_ifrd_o_4,
	exmem_ifjal_o,
	exmem_iflui_o,
	exmem_ifnext_pc_o_1,
	exmem_ifmemToReg_o,
	fuifrtReplace_1,
	idex_ifimm_o_1,
	idex_ifrdat2_o_1,
	idex_ifimm_o_0,
	idex_ifrdat2_o_0,
	exmem_ifnext_pc_o_0,
	fuifrtReplace_0,
	exmem_ifnext_pc_o_2,
	exmem_ifnext_pc_o_4,
	exmem_ifnext_pc_o_3,
	idex_ifimm_o_2,
	idex_ifrdat2_o_2,
	fuifrtReplace_2,
	exmem_ifnext_pc_o_8,
	exmem_ifnext_pc_o_7,
	exmem_ifnext_pc_o_6,
	exmem_ifnext_pc_o_5,
	idex_ifrdat2_o_3,
	idex_ifimm_o_3,
	fuifrtReplace_3,
	exmem_ifimm_o_0,
	exmem_ifnext_pc_o_16,
	exmem_ifnext_pc_o_15,
	exmem_ifnext_pc_o_14,
	exmem_ifnext_pc_o_13,
	exmem_ifnext_pc_o_12,
	exmem_ifnext_pc_o_11,
	exmem_ifnext_pc_o_10,
	exmem_ifnext_pc_o_9,
	idex_ifrdat2_o_4,
	idex_ifimm_o_4,
	fuifrtReplace_4,
	exmem_ifnext_pc_o_31,
	exmem_ifimm_o_15,
	exmem_ifnext_pc_o_29,
	exmem_ifimm_o_13,
	exmem_ifimm_o_14,
	exmem_ifnext_pc_o_30,
	exmem_ifimm_o_12,
	exmem_ifnext_pc_o_28,
	exmem_ifimm_o_10,
	exmem_ifnext_pc_o_26,
	exmem_ifnext_pc_o_27,
	exmem_ifimm_o_11,
	exmem_ifnext_pc_o_25,
	exmem_ifimm_o_9,
	exmem_ifimm_o_8,
	exmem_ifnext_pc_o_24,
	exmem_ifimm_o_6,
	exmem_ifnext_pc_o_22,
	exmem_ifnext_pc_o_23,
	exmem_ifimm_o_7,
	exmem_ifnext_pc_o_21,
	exmem_ifimm_o_5,
	exmem_ifimm_o_4,
	exmem_ifnext_pc_o_20,
	exmem_ifimm_o_2,
	exmem_ifnext_pc_o_18,
	exmem_ifnext_pc_o_19,
	exmem_ifimm_o_3,
	exmem_ifnext_pc_o_17,
	exmem_ifimm_o_1,
	idex_ifimm_o_15,
	idex_ifrdat2_o_31,
	fuifrtReplace_31,
	idex_ifrdat2_o_16,
	fuifrtReplace_16,
	idex_ifrdat2_o_17,
	fuifrtReplace_17,
	idex_ifrdat2_o_18,
	fuifrtReplace_18,
	idex_ifrdat2_o_19,
	fuifrtReplace_19,
	idex_ifrdat2_o_20,
	fuifrtReplace_20,
	idex_ifrdat2_o_21,
	fuifrtReplace_21,
	idex_ifrdat2_o_22,
	fuifrtReplace_22,
	idex_ifrdat2_o_23,
	fuifrtReplace_23,
	idex_ifrdat2_o_24,
	fuifrtReplace_24,
	idex_ifrdat2_o_25,
	fuifrtReplace_25,
	idex_ifrdat2_o_26,
	fuifrtReplace_26,
	idex_ifrdat2_o_5,
	idex_ifimm_o_5,
	fuifrtReplace_5,
	idex_ifrdat2_o_6,
	idex_ifimm_o_6,
	fuifrtReplace_6,
	idex_ifrdat2_o_7,
	idex_ifimm_o_7,
	fuifrtReplace_7,
	idex_ifrdat2_o_8,
	idex_ifimm_o_8,
	fuifrtReplace_8,
	idex_ifrdat2_o_27,
	fuifrtReplace_27,
	idex_ifrdat2_o_28,
	fuifrtReplace_28,
	idex_ifrdat2_o_29,
	fuifrtReplace_29,
	idex_ifrdat2_o_30,
	fuifrtReplace_30,
	idex_ifrdat2_o_9,
	idex_ifimm_o_9,
	fuifrtReplace_9,
	idex_ifrdat2_o_14,
	idex_ifimm_o_14,
	fuifrtReplace_14,
	idex_ifrdat2_o_15,
	fuifrtReplace_15,
	idex_ifrdat2_o_10,
	idex_ifimm_o_10,
	fuifrtReplace_10,
	idex_ifrdat2_o_11,
	idex_ifimm_o_11,
	fuifrtReplace_11,
	idex_ifrdat2_o_12,
	idex_ifimm_o_12,
	fuifrtReplace_12,
	idex_ifrdat2_o_13,
	idex_ifimm_o_13,
	fuifrtReplace_13,
	idex_ifaluop_o_3,
	myifout_1,
	ramstate,
	exmem_ifimm_o_01,
	idex_ifdWEN_o,
	idex_ifdREN_o,
	idex_ifnext_pc_o_1,
	myifout_6,
	myifout_4,
	myifout_24,
	myifout_26,
	myifout_25,
	myifout_27,
	myifout_5,
	myifout_7,
	myifout_13,
	myifout_9,
	myifout_8,
	myifout_14,
	myifout_12,
	myifout_15,
	myifout_10,
	myifout_11,
	myifout_23,
	myifout_16,
	myifout_17,
	myifout_18,
	myifout_19,
	myifout_30,
	myifout_21,
	myifnegative,
	myifout_22,
	myifout_20,
	myifout_0,
	myifout_28,
	myifout_29,
	myifout_2,
	myifout_3,
	myifout_31,
	myifout_210,
	idex_ifnext_pc_o_0,
	idex_ifnext_pc_o_3,
	idex_ifnext_pc_o_2,
	idex_ifnext_pc_o_5,
	idex_ifnext_pc_o_4,
	idex_ifnext_pc_o_7,
	idex_ifnext_pc_o_6,
	idex_ifnext_pc_o_9,
	idex_ifnext_pc_o_8,
	idex_ifnext_pc_o_11,
	idex_ifnext_pc_o_10,
	idex_ifnext_pc_o_13,
	idex_ifnext_pc_o_12,
	idex_ifnext_pc_o_15,
	idex_ifnext_pc_o_14,
	idex_ifnext_pc_o_17,
	idex_ifnext_pc_o_16,
	idex_ifnext_pc_o_19,
	idex_ifnext_pc_o_18,
	idex_ifnext_pc_o_21,
	idex_ifnext_pc_o_20,
	idex_ifnext_pc_o_23,
	idex_ifnext_pc_o_22,
	idex_ifnext_pc_o_25,
	idex_ifnext_pc_o_24,
	idex_ifnext_pc_o_27,
	idex_ifnext_pc_o_26,
	idex_ifnext_pc_o_29,
	idex_ifnext_pc_o_28,
	idex_ifnext_pc_o_31,
	idex_ifnext_pc_o_30,
	exmem_ifrdat2_o_1,
	exmem_ifrdat2_o_2,
	exmem_ifrdat2_o_3,
	exmem_ifrdat2_o_4,
	exmem_ifrdat2_o_5,
	exmem_ifrdat2_o_6,
	exmem_ifrdat2_o_7,
	exmem_ifrdat2_o_8,
	exmem_ifrdat2_o_9,
	exmem_ifrdat2_o_10,
	exmem_ifrdat2_o_11,
	exmem_ifrdat2_o_12,
	exmem_ifrdat2_o_13,
	exmem_ifrdat2_o_14,
	exmem_ifrdat2_o_15,
	exmem_ifrdat2_o_16,
	exmem_ifrdat2_o_17,
	exmem_ifrdat2_o_18,
	exmem_ifrdat2_o_19,
	exmem_ifrdat2_o_20,
	exmem_ifrdat2_o_21,
	exmem_ifrdat2_o_22,
	exmem_ifrdat2_o_23,
	exmem_ifrdat2_o_24,
	exmem_ifrdat2_o_25,
	exmem_ifrdat2_o_26,
	exmem_ifrdat2_o_27,
	exmem_ifrdat2_o_28,
	exmem_ifrdat2_o_29,
	exmem_ifrdat2_o_30,
	exmem_ifrdat2_o_31,
	idex_ifhalt_o,
	fuifrdat2_ow,
	idex_ifRegDest_o_1,
	idex_ifrd_o_1,
	idex_ifRegDest_o_0,
	idex_ifrd_o_0,
	idex_ifrd_o_3,
	idex_ifrd_o_2,
	idex_ifregWEN_o,
	idex_ifrd_o_4,
	idex_ifjal_o,
	idex_iflui_o,
	idex_ifmemToReg_o,
	myifout_32,
	CPUCLK,
	nRST,
	devpor,
	devclrn,
	devoe);
output 	exmem_ifout_o_1;
output 	exmem_ifdWEN_o;
output 	exmem_ifdREN_o;
output 	exmem_ifout_o_0;
output 	exmem_ifout_o_3;
output 	exmem_ifout_o_2;
output 	exmem_ifout_o_5;
output 	exmem_ifout_o_4;
output 	exmem_ifout_o_7;
output 	exmem_ifout_o_6;
output 	exmem_ifout_o_9;
output 	exmem_ifout_o_8;
output 	exmem_ifout_o_11;
output 	exmem_ifout_o_10;
output 	exmem_ifout_o_13;
output 	exmem_ifout_o_12;
output 	exmem_ifout_o_15;
output 	exmem_ifout_o_14;
output 	exmem_ifout_o_17;
output 	exmem_ifout_o_16;
output 	exmem_ifout_o_19;
output 	exmem_ifout_o_18;
output 	exmem_ifout_o_21;
output 	exmem_ifout_o_20;
output 	exmem_ifout_o_23;
output 	exmem_ifout_o_22;
output 	exmem_ifout_o_25;
output 	exmem_ifout_o_24;
output 	exmem_ifout_o_27;
output 	exmem_ifout_o_26;
output 	exmem_ifout_o_29;
output 	exmem_ifout_o_28;
output 	exmem_ifout_o_31;
output 	exmem_ifout_o_30;
input 	always1;
input 	always11;
output 	exmem_ifhalt_o;
output 	exmem_ifrdat2_o_0;
input 	always12;
input 	idex_ifrt_o_0;
input 	idex_ifrt_o_1;
output 	exmem_ifRegDest_o_1;
output 	exmem_ifrt_o_1;
output 	exmem_ifrd_o_1;
output 	exmem_ifRegDest_o_0;
output 	exmem_ifrt_o_0;
output 	exmem_ifrd_o_0;
input 	idex_ifrt_o_2;
input 	idex_ifrt_o_3;
output 	exmem_ifrt_o_3;
output 	exmem_ifrd_o_3;
output 	exmem_ifrt_o_2;
output 	exmem_ifrd_o_2;
output 	exmem_ifregWEN_o;
input 	idex_ifrt_o_4;
output 	exmem_ifrt_o_4;
output 	exmem_ifrd_o_4;
output 	exmem_ifjal_o;
output 	exmem_iflui_o;
output 	exmem_ifnext_pc_o_1;
output 	exmem_ifmemToReg_o;
input 	fuifrtReplace_1;
input 	idex_ifimm_o_1;
input 	idex_ifrdat2_o_1;
input 	idex_ifimm_o_0;
input 	idex_ifrdat2_o_0;
output 	exmem_ifnext_pc_o_0;
input 	fuifrtReplace_0;
output 	exmem_ifnext_pc_o_2;
output 	exmem_ifnext_pc_o_4;
output 	exmem_ifnext_pc_o_3;
input 	idex_ifimm_o_2;
input 	idex_ifrdat2_o_2;
input 	fuifrtReplace_2;
output 	exmem_ifnext_pc_o_8;
output 	exmem_ifnext_pc_o_7;
output 	exmem_ifnext_pc_o_6;
output 	exmem_ifnext_pc_o_5;
input 	idex_ifrdat2_o_3;
input 	idex_ifimm_o_3;
input 	fuifrtReplace_3;
output 	exmem_ifimm_o_0;
output 	exmem_ifnext_pc_o_16;
output 	exmem_ifnext_pc_o_15;
output 	exmem_ifnext_pc_o_14;
output 	exmem_ifnext_pc_o_13;
output 	exmem_ifnext_pc_o_12;
output 	exmem_ifnext_pc_o_11;
output 	exmem_ifnext_pc_o_10;
output 	exmem_ifnext_pc_o_9;
input 	idex_ifrdat2_o_4;
input 	idex_ifimm_o_4;
input 	fuifrtReplace_4;
output 	exmem_ifnext_pc_o_31;
output 	exmem_ifimm_o_15;
output 	exmem_ifnext_pc_o_29;
output 	exmem_ifimm_o_13;
output 	exmem_ifimm_o_14;
output 	exmem_ifnext_pc_o_30;
output 	exmem_ifimm_o_12;
output 	exmem_ifnext_pc_o_28;
output 	exmem_ifimm_o_10;
output 	exmem_ifnext_pc_o_26;
output 	exmem_ifnext_pc_o_27;
output 	exmem_ifimm_o_11;
output 	exmem_ifnext_pc_o_25;
output 	exmem_ifimm_o_9;
output 	exmem_ifimm_o_8;
output 	exmem_ifnext_pc_o_24;
output 	exmem_ifimm_o_6;
output 	exmem_ifnext_pc_o_22;
output 	exmem_ifnext_pc_o_23;
output 	exmem_ifimm_o_7;
output 	exmem_ifnext_pc_o_21;
output 	exmem_ifimm_o_5;
output 	exmem_ifimm_o_4;
output 	exmem_ifnext_pc_o_20;
output 	exmem_ifimm_o_2;
output 	exmem_ifnext_pc_o_18;
output 	exmem_ifnext_pc_o_19;
output 	exmem_ifimm_o_3;
output 	exmem_ifnext_pc_o_17;
output 	exmem_ifimm_o_1;
input 	idex_ifimm_o_15;
input 	idex_ifrdat2_o_31;
input 	fuifrtReplace_31;
input 	idex_ifrdat2_o_16;
input 	fuifrtReplace_16;
input 	idex_ifrdat2_o_17;
input 	fuifrtReplace_17;
input 	idex_ifrdat2_o_18;
input 	fuifrtReplace_18;
input 	idex_ifrdat2_o_19;
input 	fuifrtReplace_19;
input 	idex_ifrdat2_o_20;
input 	fuifrtReplace_20;
input 	idex_ifrdat2_o_21;
input 	fuifrtReplace_21;
input 	idex_ifrdat2_o_22;
input 	fuifrtReplace_22;
input 	idex_ifrdat2_o_23;
input 	fuifrtReplace_23;
input 	idex_ifrdat2_o_24;
input 	fuifrtReplace_24;
input 	idex_ifrdat2_o_25;
input 	fuifrtReplace_25;
input 	idex_ifrdat2_o_26;
input 	fuifrtReplace_26;
input 	idex_ifrdat2_o_5;
input 	idex_ifimm_o_5;
input 	fuifrtReplace_5;
input 	idex_ifrdat2_o_6;
input 	idex_ifimm_o_6;
input 	fuifrtReplace_6;
input 	idex_ifrdat2_o_7;
input 	idex_ifimm_o_7;
input 	fuifrtReplace_7;
input 	idex_ifrdat2_o_8;
input 	idex_ifimm_o_8;
input 	fuifrtReplace_8;
input 	idex_ifrdat2_o_27;
input 	fuifrtReplace_27;
input 	idex_ifrdat2_o_28;
input 	fuifrtReplace_28;
input 	idex_ifrdat2_o_29;
input 	fuifrtReplace_29;
input 	idex_ifrdat2_o_30;
input 	fuifrtReplace_30;
input 	idex_ifrdat2_o_9;
input 	idex_ifimm_o_9;
input 	fuifrtReplace_9;
input 	idex_ifrdat2_o_14;
input 	idex_ifimm_o_14;
input 	fuifrtReplace_14;
input 	idex_ifrdat2_o_15;
input 	fuifrtReplace_15;
input 	idex_ifrdat2_o_10;
input 	idex_ifimm_o_10;
input 	fuifrtReplace_10;
input 	idex_ifrdat2_o_11;
input 	idex_ifimm_o_11;
input 	fuifrtReplace_11;
input 	idex_ifrdat2_o_12;
input 	idex_ifimm_o_12;
input 	fuifrtReplace_12;
input 	idex_ifrdat2_o_13;
input 	idex_ifimm_o_13;
input 	fuifrtReplace_13;
input 	idex_ifaluop_o_3;
input 	myifout_1;
input 	ramstate;
output 	exmem_ifimm_o_01;
input 	idex_ifdWEN_o;
input 	idex_ifdREN_o;
input 	idex_ifnext_pc_o_1;
input 	myifout_6;
input 	myifout_4;
input 	myifout_24;
input 	myifout_26;
input 	myifout_25;
input 	myifout_27;
input 	myifout_5;
input 	myifout_7;
input 	myifout_13;
input 	myifout_9;
input 	myifout_8;
input 	myifout_14;
input 	myifout_12;
input 	myifout_15;
input 	myifout_10;
input 	myifout_11;
input 	myifout_23;
input 	myifout_16;
input 	myifout_17;
input 	myifout_18;
input 	myifout_19;
input 	myifout_30;
input 	myifout_21;
input 	myifnegative;
input 	myifout_22;
input 	myifout_20;
input 	myifout_0;
input 	myifout_28;
input 	myifout_29;
input 	myifout_2;
input 	myifout_3;
input 	myifout_31;
input 	myifout_210;
input 	idex_ifnext_pc_o_0;
input 	idex_ifnext_pc_o_3;
input 	idex_ifnext_pc_o_2;
input 	idex_ifnext_pc_o_5;
input 	idex_ifnext_pc_o_4;
input 	idex_ifnext_pc_o_7;
input 	idex_ifnext_pc_o_6;
input 	idex_ifnext_pc_o_9;
input 	idex_ifnext_pc_o_8;
input 	idex_ifnext_pc_o_11;
input 	idex_ifnext_pc_o_10;
input 	idex_ifnext_pc_o_13;
input 	idex_ifnext_pc_o_12;
input 	idex_ifnext_pc_o_15;
input 	idex_ifnext_pc_o_14;
input 	idex_ifnext_pc_o_17;
input 	idex_ifnext_pc_o_16;
input 	idex_ifnext_pc_o_19;
input 	idex_ifnext_pc_o_18;
input 	idex_ifnext_pc_o_21;
input 	idex_ifnext_pc_o_20;
input 	idex_ifnext_pc_o_23;
input 	idex_ifnext_pc_o_22;
input 	idex_ifnext_pc_o_25;
input 	idex_ifnext_pc_o_24;
input 	idex_ifnext_pc_o_27;
input 	idex_ifnext_pc_o_26;
input 	idex_ifnext_pc_o_29;
input 	idex_ifnext_pc_o_28;
input 	idex_ifnext_pc_o_31;
input 	idex_ifnext_pc_o_30;
output 	exmem_ifrdat2_o_1;
output 	exmem_ifrdat2_o_2;
output 	exmem_ifrdat2_o_3;
output 	exmem_ifrdat2_o_4;
output 	exmem_ifrdat2_o_5;
output 	exmem_ifrdat2_o_6;
output 	exmem_ifrdat2_o_7;
output 	exmem_ifrdat2_o_8;
output 	exmem_ifrdat2_o_9;
output 	exmem_ifrdat2_o_10;
output 	exmem_ifrdat2_o_11;
output 	exmem_ifrdat2_o_12;
output 	exmem_ifrdat2_o_13;
output 	exmem_ifrdat2_o_14;
output 	exmem_ifrdat2_o_15;
output 	exmem_ifrdat2_o_16;
output 	exmem_ifrdat2_o_17;
output 	exmem_ifrdat2_o_18;
output 	exmem_ifrdat2_o_19;
output 	exmem_ifrdat2_o_20;
output 	exmem_ifrdat2_o_21;
output 	exmem_ifrdat2_o_22;
output 	exmem_ifrdat2_o_23;
output 	exmem_ifrdat2_o_24;
output 	exmem_ifrdat2_o_25;
output 	exmem_ifrdat2_o_26;
output 	exmem_ifrdat2_o_27;
output 	exmem_ifrdat2_o_28;
output 	exmem_ifrdat2_o_29;
output 	exmem_ifrdat2_o_30;
output 	exmem_ifrdat2_o_31;
input 	idex_ifhalt_o;
input 	fuifrdat2_ow;
input 	idex_ifRegDest_o_1;
input 	idex_ifrd_o_1;
input 	idex_ifRegDest_o_0;
input 	idex_ifrd_o_0;
input 	idex_ifrd_o_3;
input 	idex_ifrd_o_2;
input 	idex_ifregWEN_o;
input 	idex_ifrd_o_4;
input 	idex_ifjal_o;
input 	idex_iflui_o;
input 	idex_ifmemToReg_o;
input 	myifout_32;
input 	CPUCLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \out_o~62_combout ;
wire \dWEN_o~0_combout ;
wire \dREN_o~0_combout ;
wire \out_o~63_combout ;
wire \out_o~60_combout ;
wire \out_o~61_combout ;
wire \out_o~64_combout ;
wire \out_o~65_combout ;
wire \out_o~66_combout ;
wire \out_o~67_combout ;
wire \out_o~68_combout ;
wire \out_o~69_combout ;
wire \out_o~70_combout ;
wire \out_o~71_combout ;
wire \out_o~72_combout ;
wire \out_o~73_combout ;
wire \out_o~74_combout ;
wire \out_o~75_combout ;
wire \out_o~76_combout ;
wire \out_o~77_combout ;
wire \out_o~78_combout ;
wire \out_o~79_combout ;
wire \out_o~80_combout ;
wire \out_o~81_combout ;
wire \out_o~82_combout ;
wire \out_o~83_combout ;
wire \out_o~84_combout ;
wire \out_o~85_combout ;
wire \out_o~86_combout ;
wire \out_o~87_combout ;
wire \out_o~88_combout ;
wire \out_o~89_combout ;
wire \out_o~90_combout ;
wire \out_o~91_combout ;
wire \halt_o~0_combout ;
wire \rdat2_o~0_combout ;
wire \RegDest_o~0_combout ;
wire \rt_o~0_combout ;
wire \rd_o~0_combout ;
wire \RegDest_o~1_combout ;
wire \rt_o~1_combout ;
wire \rd_o~1_combout ;
wire \rt_o~2_combout ;
wire \rd_o~2_combout ;
wire \rt_o~3_combout ;
wire \rd_o~3_combout ;
wire \regWEN_o~0_combout ;
wire \rt_o~4_combout ;
wire \rd_o~4_combout ;
wire \jal_o~0_combout ;
wire \lui_o~0_combout ;
wire \next_pc_o~0_combout ;
wire \memToReg_o~0_combout ;
wire \next_pc_o~1_combout ;
wire \next_pc_o~2_combout ;
wire \next_pc_o~3_combout ;
wire \exmem_if.next_pc_o[4]~feeder_combout ;
wire \next_pc_o~4_combout ;
wire \next_pc_o~5_combout ;
wire \next_pc_o~6_combout ;
wire \next_pc_o~7_combout ;
wire \next_pc_o~8_combout ;
wire \imm_o~0_combout ;
wire \next_pc_o~9_combout ;
wire \next_pc_o~10_combout ;
wire \next_pc_o~11_combout ;
wire \next_pc_o~12_combout ;
wire \next_pc_o~13_combout ;
wire \next_pc_o~14_combout ;
wire \next_pc_o~15_combout ;
wire \next_pc_o~16_combout ;
wire \next_pc_o~17_combout ;
wire \imm_o~1_combout ;
wire \next_pc_o~18_combout ;
wire \imm_o~2_combout ;
wire \imm_o~3_combout ;
wire \next_pc_o~19_combout ;
wire \imm_o~4_combout ;
wire \next_pc_o~20_combout ;
wire \imm_o~5_combout ;
wire \next_pc_o~21_combout ;
wire \next_pc_o~22_combout ;
wire \imm_o~6_combout ;
wire \next_pc_o~23_combout ;
wire \imm_o~7_combout ;
wire \imm_o~8_combout ;
wire \next_pc_o~24_combout ;
wire \imm_o~9_combout ;
wire \next_pc_o~25_combout ;
wire \next_pc_o~26_combout ;
wire \imm_o~10_combout ;
wire \next_pc_o~27_combout ;
wire \exmem_if.next_pc_o[21]~feeder_combout ;
wire \imm_o~11_combout ;
wire \imm_o~12_combout ;
wire \next_pc_o~28_combout ;
wire \imm_o~13_combout ;
wire \next_pc_o~29_combout ;
wire \next_pc_o~30_combout ;
wire \imm_o~14_combout ;
wire \next_pc_o~31_combout ;
wire \imm_o~15_combout ;
wire \rdat2_o~1_combout ;
wire \rdat2_o~2_combout ;
wire \rdat2_o~3_combout ;
wire \rdat2_o~4_combout ;
wire \rdat2_o~5_combout ;
wire \rdat2_o~6_combout ;
wire \rdat2_o~7_combout ;
wire \rdat2_o~8_combout ;
wire \rdat2_o~9_combout ;
wire \rdat2_o~10_combout ;
wire \rdat2_o~11_combout ;
wire \rdat2_o~12_combout ;
wire \rdat2_o~13_combout ;
wire \rdat2_o~14_combout ;
wire \rdat2_o~15_combout ;
wire \rdat2_o~16_combout ;
wire \rdat2_o~17_combout ;
wire \rdat2_o~18_combout ;
wire \rdat2_o~19_combout ;
wire \rdat2_o~20_combout ;
wire \rdat2_o~21_combout ;
wire \rdat2_o~22_combout ;
wire \rdat2_o~23_combout ;
wire \rdat2_o~24_combout ;
wire \rdat2_o~25_combout ;
wire \rdat2_o~26_combout ;
wire \rdat2_o~27_combout ;
wire \rdat2_o~28_combout ;
wire \rdat2_o~29_combout ;
wire \rdat2_o~30_combout ;
wire \rdat2_o~31_combout ;


// Location: FF_X53_Y33_N1
dffeas \exmem_if.out_o[1] (
	.clk(CPUCLK),
	.d(\out_o~62_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[1] .is_wysiwyg = "true";
defparam \exmem_if.out_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N9
dffeas \exmem_if.dWEN_o (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\dWEN_o~0_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifdWEN_o),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.dWEN_o .is_wysiwyg = "true";
defparam \exmem_if.dWEN_o .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N25
dffeas \exmem_if.dREN_o (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\dREN_o~0_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifdREN_o),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.dREN_o .is_wysiwyg = "true";
defparam \exmem_if.dREN_o .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N25
dffeas \exmem_if.out_o[0] (
	.clk(CPUCLK),
	.d(\out_o~63_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[0] .is_wysiwyg = "true";
defparam \exmem_if.out_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N17
dffeas \exmem_if.out_o[3] (
	.clk(CPUCLK),
	.d(\out_o~60_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[3] .is_wysiwyg = "true";
defparam \exmem_if.out_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N17
dffeas \exmem_if.out_o[2] (
	.clk(CPUCLK),
	.d(\out_o~61_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[2] .is_wysiwyg = "true";
defparam \exmem_if.out_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N31
dffeas \exmem_if.out_o[5] (
	.clk(CPUCLK),
	.d(\out_o~64_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_5),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[5] .is_wysiwyg = "true";
defparam \exmem_if.out_o[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y28_N9
dffeas \exmem_if.out_o[4] (
	.clk(CPUCLK),
	.d(\out_o~65_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[4] .is_wysiwyg = "true";
defparam \exmem_if.out_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N17
dffeas \exmem_if.out_o[7] (
	.clk(CPUCLK),
	.d(\out_o~66_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_7),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[7] .is_wysiwyg = "true";
defparam \exmem_if.out_o[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N7
dffeas \exmem_if.out_o[6] (
	.clk(CPUCLK),
	.d(\out_o~67_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_6),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[6] .is_wysiwyg = "true";
defparam \exmem_if.out_o[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N27
dffeas \exmem_if.out_o[9] (
	.clk(CPUCLK),
	.d(\out_o~68_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_9),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[9] .is_wysiwyg = "true";
defparam \exmem_if.out_o[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N15
dffeas \exmem_if.out_o[8] (
	.clk(CPUCLK),
	.d(\out_o~69_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_8),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[8] .is_wysiwyg = "true";
defparam \exmem_if.out_o[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N7
dffeas \exmem_if.out_o[11] (
	.clk(CPUCLK),
	.d(\out_o~70_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_11),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[11] .is_wysiwyg = "true";
defparam \exmem_if.out_o[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N23
dffeas \exmem_if.out_o[10] (
	.clk(CPUCLK),
	.d(\out_o~71_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_10),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[10] .is_wysiwyg = "true";
defparam \exmem_if.out_o[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N9
dffeas \exmem_if.out_o[13] (
	.clk(CPUCLK),
	.d(\out_o~72_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_13),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[13] .is_wysiwyg = "true";
defparam \exmem_if.out_o[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N15
dffeas \exmem_if.out_o[12] (
	.clk(CPUCLK),
	.d(\out_o~73_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_12),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[12] .is_wysiwyg = "true";
defparam \exmem_if.out_o[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N17
dffeas \exmem_if.out_o[15] (
	.clk(CPUCLK),
	.d(\out_o~74_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_15),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[15] .is_wysiwyg = "true";
defparam \exmem_if.out_o[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N19
dffeas \exmem_if.out_o[14] (
	.clk(CPUCLK),
	.d(\out_o~75_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_14),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[14] .is_wysiwyg = "true";
defparam \exmem_if.out_o[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N21
dffeas \exmem_if.out_o[17] (
	.clk(CPUCLK),
	.d(\out_o~76_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_17),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[17] .is_wysiwyg = "true";
defparam \exmem_if.out_o[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N7
dffeas \exmem_if.out_o[16] (
	.clk(CPUCLK),
	.d(\out_o~77_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_16),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[16] .is_wysiwyg = "true";
defparam \exmem_if.out_o[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N17
dffeas \exmem_if.out_o[19] (
	.clk(CPUCLK),
	.d(\out_o~78_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_19),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[19] .is_wysiwyg = "true";
defparam \exmem_if.out_o[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N27
dffeas \exmem_if.out_o[18] (
	.clk(CPUCLK),
	.d(\out_o~79_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_18),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[18] .is_wysiwyg = "true";
defparam \exmem_if.out_o[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N23
dffeas \exmem_if.out_o[21] (
	.clk(CPUCLK),
	.d(\out_o~80_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_21),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[21] .is_wysiwyg = "true";
defparam \exmem_if.out_o[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N7
dffeas \exmem_if.out_o[20] (
	.clk(CPUCLK),
	.d(\out_o~81_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_20),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[20] .is_wysiwyg = "true";
defparam \exmem_if.out_o[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N17
dffeas \exmem_if.out_o[23] (
	.clk(CPUCLK),
	.d(\out_o~82_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_23),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[23] .is_wysiwyg = "true";
defparam \exmem_if.out_o[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N13
dffeas \exmem_if.out_o[22] (
	.clk(CPUCLK),
	.d(\out_o~83_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_22),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[22] .is_wysiwyg = "true";
defparam \exmem_if.out_o[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N15
dffeas \exmem_if.out_o[25] (
	.clk(CPUCLK),
	.d(\out_o~84_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_25),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[25] .is_wysiwyg = "true";
defparam \exmem_if.out_o[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N1
dffeas \exmem_if.out_o[24] (
	.clk(CPUCLK),
	.d(\out_o~85_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_24),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[24] .is_wysiwyg = "true";
defparam \exmem_if.out_o[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N29
dffeas \exmem_if.out_o[27] (
	.clk(CPUCLK),
	.d(\out_o~86_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_27),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[27] .is_wysiwyg = "true";
defparam \exmem_if.out_o[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N29
dffeas \exmem_if.out_o[26] (
	.clk(CPUCLK),
	.d(\out_o~87_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_26),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[26] .is_wysiwyg = "true";
defparam \exmem_if.out_o[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N9
dffeas \exmem_if.out_o[29] (
	.clk(CPUCLK),
	.d(\out_o~88_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_29),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[29] .is_wysiwyg = "true";
defparam \exmem_if.out_o[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N5
dffeas \exmem_if.out_o[28] (
	.clk(CPUCLK),
	.d(\out_o~89_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_28),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[28] .is_wysiwyg = "true";
defparam \exmem_if.out_o[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N31
dffeas \exmem_if.out_o[31] (
	.clk(CPUCLK),
	.d(\out_o~90_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_31),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[31] .is_wysiwyg = "true";
defparam \exmem_if.out_o[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N5
dffeas \exmem_if.out_o[30] (
	.clk(CPUCLK),
	.d(\out_o~91_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifout_o_30),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.out_o[30] .is_wysiwyg = "true";
defparam \exmem_if.out_o[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N29
dffeas \exmem_if.halt_o (
	.clk(CPUCLK),
	.d(\halt_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifhalt_o),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.halt_o .is_wysiwyg = "true";
defparam \exmem_if.halt_o .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N1
dffeas \exmem_if.rdat2_o[0] (
	.clk(CPUCLK),
	.d(\rdat2_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[0] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N19
dffeas \exmem_if.RegDest_o[1] (
	.clk(CPUCLK),
	.d(\RegDest_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifRegDest_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.RegDest_o[1] .is_wysiwyg = "true";
defparam \exmem_if.RegDest_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N21
dffeas \exmem_if.rt_o[1] (
	.clk(CPUCLK),
	.d(\rt_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrt_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rt_o[1] .is_wysiwyg = "true";
defparam \exmem_if.rt_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N19
dffeas \exmem_if.rd_o[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\rd_o~0_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrd_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rd_o[1] .is_wysiwyg = "true";
defparam \exmem_if.rd_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N7
dffeas \exmem_if.RegDest_o[0] (
	.clk(CPUCLK),
	.d(\RegDest_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifRegDest_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.RegDest_o[0] .is_wysiwyg = "true";
defparam \exmem_if.RegDest_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N17
dffeas \exmem_if.rt_o[0] (
	.clk(CPUCLK),
	.d(\rt_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrt_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rt_o[0] .is_wysiwyg = "true";
defparam \exmem_if.rt_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N27
dffeas \exmem_if.rd_o[0] (
	.clk(CPUCLK),
	.d(\rd_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrd_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rd_o[0] .is_wysiwyg = "true";
defparam \exmem_if.rd_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N23
dffeas \exmem_if.rt_o[3] (
	.clk(CPUCLK),
	.d(\rt_o~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrt_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rt_o[3] .is_wysiwyg = "true";
defparam \exmem_if.rt_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N13
dffeas \exmem_if.rd_o[3] (
	.clk(CPUCLK),
	.d(\rd_o~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrd_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rd_o[3] .is_wysiwyg = "true";
defparam \exmem_if.rd_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N9
dffeas \exmem_if.rt_o[2] (
	.clk(CPUCLK),
	.d(\rt_o~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrt_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rt_o[2] .is_wysiwyg = "true";
defparam \exmem_if.rt_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N11
dffeas \exmem_if.rd_o[2] (
	.clk(CPUCLK),
	.d(\rd_o~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrd_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rd_o[2] .is_wysiwyg = "true";
defparam \exmem_if.rd_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N15
dffeas \exmem_if.regWEN_o (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\regWEN_o~0_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifregWEN_o),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.regWEN_o .is_wysiwyg = "true";
defparam \exmem_if.regWEN_o .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y31_N31
dffeas \exmem_if.rt_o[4] (
	.clk(CPUCLK),
	.d(\rt_o~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrt_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rt_o[4] .is_wysiwyg = "true";
defparam \exmem_if.rt_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N5
dffeas \exmem_if.rd_o[4] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\rd_o~4_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrd_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rd_o[4] .is_wysiwyg = "true";
defparam \exmem_if.rd_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N17
dffeas \exmem_if.jal_o (
	.clk(CPUCLK),
	.d(\jal_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifjal_o),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.jal_o .is_wysiwyg = "true";
defparam \exmem_if.jal_o .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N27
dffeas \exmem_if.lui_o (
	.clk(CPUCLK),
	.d(\lui_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_iflui_o),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.lui_o .is_wysiwyg = "true";
defparam \exmem_if.lui_o .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N11
dffeas \exmem_if.next_pc_o[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\next_pc_o~0_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[1] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N9
dffeas \exmem_if.memToReg_o (
	.clk(CPUCLK),
	.d(\memToReg_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifmemToReg_o),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.memToReg_o .is_wysiwyg = "true";
defparam \exmem_if.memToReg_o .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N23
dffeas \exmem_if.next_pc_o[0] (
	.clk(CPUCLK),
	.d(\next_pc_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[0] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N13
dffeas \exmem_if.next_pc_o[2] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\next_pc_o~2_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[2] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N5
dffeas \exmem_if.next_pc_o[4] (
	.clk(CPUCLK),
	.d(\exmem_if.next_pc_o[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[4] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N13
dffeas \exmem_if.next_pc_o[3] (
	.clk(CPUCLK),
	.d(\next_pc_o~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[3] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N27
dffeas \exmem_if.next_pc_o[8] (
	.clk(CPUCLK),
	.d(\next_pc_o~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_8),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[8] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N9
dffeas \exmem_if.next_pc_o[7] (
	.clk(CPUCLK),
	.d(\next_pc_o~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_7),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[7] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N29
dffeas \exmem_if.next_pc_o[6] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\next_pc_o~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_6),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[6] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N21
dffeas \exmem_if.next_pc_o[5] (
	.clk(CPUCLK),
	.d(\next_pc_o~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_5),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[5] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N19
dffeas \exmem_if.imm_o[0] (
	.clk(CPUCLK),
	.d(\imm_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifimm_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.imm_o[0] .is_wysiwyg = "true";
defparam \exmem_if.imm_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N13
dffeas \exmem_if.next_pc_o[16] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\next_pc_o~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_16),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[16] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N21
dffeas \exmem_if.next_pc_o[15] (
	.clk(CPUCLK),
	.d(\next_pc_o~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_15),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[15] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N31
dffeas \exmem_if.next_pc_o[14] (
	.clk(CPUCLK),
	.d(\next_pc_o~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_14),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[14] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N15
dffeas \exmem_if.next_pc_o[13] (
	.clk(CPUCLK),
	.d(\next_pc_o~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_13),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[13] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N5
dffeas \exmem_if.next_pc_o[12] (
	.clk(CPUCLK),
	.d(\next_pc_o~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_12),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[12] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N17
dffeas \exmem_if.next_pc_o[11] (
	.clk(CPUCLK),
	.d(\next_pc_o~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_11),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[11] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N31
dffeas \exmem_if.next_pc_o[10] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\next_pc_o~15_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_10),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[10] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N31
dffeas \exmem_if.next_pc_o[9] (
	.clk(CPUCLK),
	.d(\next_pc_o~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_9),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[9] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N25
dffeas \exmem_if.next_pc_o[31] (
	.clk(CPUCLK),
	.d(\next_pc_o~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_31),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[31] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N15
dffeas \exmem_if.imm_o[15] (
	.clk(CPUCLK),
	.d(\imm_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifimm_o_15),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.imm_o[15] .is_wysiwyg = "true";
defparam \exmem_if.imm_o[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N23
dffeas \exmem_if.next_pc_o[29] (
	.clk(CPUCLK),
	.d(\next_pc_o~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_29),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[29] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N21
dffeas \exmem_if.imm_o[13] (
	.clk(CPUCLK),
	.d(\imm_o~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifimm_o_13),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.imm_o[13] .is_wysiwyg = "true";
defparam \exmem_if.imm_o[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y35_N9
dffeas \exmem_if.imm_o[14] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~3_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifimm_o_14),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.imm_o[14] .is_wysiwyg = "true";
defparam \exmem_if.imm_o[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y34_N25
dffeas \exmem_if.next_pc_o[30] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\next_pc_o~19_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_30),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[30] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N23
dffeas \exmem_if.imm_o[12] (
	.clk(CPUCLK),
	.d(\imm_o~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifimm_o_12),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.imm_o[12] .is_wysiwyg = "true";
defparam \exmem_if.imm_o[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N27
dffeas \exmem_if.next_pc_o[28] (
	.clk(CPUCLK),
	.d(\next_pc_o~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_28),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[28] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N9
dffeas \exmem_if.imm_o[10] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifimm_o_10),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.imm_o[10] .is_wysiwyg = "true";
defparam \exmem_if.imm_o[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N25
dffeas \exmem_if.next_pc_o[26] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\next_pc_o~21_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_26),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[26] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N5
dffeas \exmem_if.next_pc_o[27] (
	.clk(CPUCLK),
	.d(\next_pc_o~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_27),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[27] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N1
dffeas \exmem_if.imm_o[11] (
	.clk(CPUCLK),
	.d(\imm_o~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifimm_o_11),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.imm_o[11] .is_wysiwyg = "true";
defparam \exmem_if.imm_o[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N13
dffeas \exmem_if.next_pc_o[25] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\next_pc_o~23_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_25),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[25] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N13
dffeas \exmem_if.imm_o[9] (
	.clk(CPUCLK),
	.d(\imm_o~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifimm_o_9),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.imm_o[9] .is_wysiwyg = "true";
defparam \exmem_if.imm_o[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N23
dffeas \exmem_if.imm_o[8] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifimm_o_8),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.imm_o[8] .is_wysiwyg = "true";
defparam \exmem_if.imm_o[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N21
dffeas \exmem_if.next_pc_o[24] (
	.clk(CPUCLK),
	.d(\next_pc_o~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_24),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[24] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N17
dffeas \exmem_if.imm_o[6] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifimm_o_6),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.imm_o[6] .is_wysiwyg = "true";
defparam \exmem_if.imm_o[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N3
dffeas \exmem_if.next_pc_o[22] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\next_pc_o~25_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_22),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[22] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N5
dffeas \exmem_if.next_pc_o[23] (
	.clk(CPUCLK),
	.d(\next_pc_o~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_23),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[23] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N21
dffeas \exmem_if.imm_o[7] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifimm_o_7),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.imm_o[7] .is_wysiwyg = "true";
defparam \exmem_if.imm_o[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N13
dffeas \exmem_if.next_pc_o[21] (
	.clk(CPUCLK),
	.d(\exmem_if.next_pc_o[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_21),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[21] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N1
dffeas \exmem_if.imm_o[5] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~11_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifimm_o_5),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.imm_o[5] .is_wysiwyg = "true";
defparam \exmem_if.imm_o[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y37_N19
dffeas \exmem_if.imm_o[4] (
	.clk(CPUCLK),
	.d(\imm_o~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifimm_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.imm_o[4] .is_wysiwyg = "true";
defparam \exmem_if.imm_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N13
dffeas \exmem_if.next_pc_o[20] (
	.clk(CPUCLK),
	.d(\next_pc_o~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_20),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[20] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y30_N7
dffeas \exmem_if.imm_o[2] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifimm_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.imm_o[2] .is_wysiwyg = "true";
defparam \exmem_if.imm_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N19
dffeas \exmem_if.next_pc_o[18] (
	.clk(CPUCLK),
	.d(\next_pc_o~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_18),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[18] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N29
dffeas \exmem_if.next_pc_o[19] (
	.clk(CPUCLK),
	.d(\next_pc_o~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_19),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[19] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N31
dffeas \exmem_if.imm_o[3] (
	.clk(CPUCLK),
	.d(\imm_o~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifimm_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.imm_o[3] .is_wysiwyg = "true";
defparam \exmem_if.imm_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N11
dffeas \exmem_if.next_pc_o[17] (
	.clk(CPUCLK),
	.d(\next_pc_o~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifnext_pc_o_17),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.next_pc_o[17] .is_wysiwyg = "true";
defparam \exmem_if.next_pc_o[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N1
dffeas \exmem_if.imm_o[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~15_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifimm_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.imm_o[1] .is_wysiwyg = "true";
defparam \exmem_if.imm_o[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N2
cycloneive_lcell_comb \exmem_if.imm_o[0]~0 (
// Equation(s):
// exmem_ifimm_o_01 = ((!ramstate & ((always1) # (always11)))) # (!always12)

	.dataa(always1),
	.datab(ramstate),
	.datac(always12),
	.datad(always11),
	.cin(gnd),
	.combout(exmem_ifimm_o_01),
	.cout());
// synopsys translate_off
defparam \exmem_if.imm_o[0]~0 .lut_mask = 16'h3F2F;
defparam \exmem_if.imm_o[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N11
dffeas \exmem_if.rdat2_o[1] (
	.clk(CPUCLK),
	.d(\rdat2_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[1] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N7
dffeas \exmem_if.rdat2_o[2] (
	.clk(CPUCLK),
	.d(\rdat2_o~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[2] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N19
dffeas \exmem_if.rdat2_o[3] (
	.clk(CPUCLK),
	.d(\rdat2_o~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[3] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N13
dffeas \exmem_if.rdat2_o[4] (
	.clk(CPUCLK),
	.d(\rdat2_o~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[4] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N21
dffeas \exmem_if.rdat2_o[5] (
	.clk(CPUCLK),
	.d(\rdat2_o~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_5),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[5] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y28_N1
dffeas \exmem_if.rdat2_o[6] (
	.clk(CPUCLK),
	.d(\rdat2_o~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_6),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[6] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N19
dffeas \exmem_if.rdat2_o[7] (
	.clk(CPUCLK),
	.d(\rdat2_o~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_7),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[7] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N27
dffeas \exmem_if.rdat2_o[8] (
	.clk(CPUCLK),
	.d(\rdat2_o~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_8),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[8] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N29
dffeas \exmem_if.rdat2_o[9] (
	.clk(CPUCLK),
	.d(\rdat2_o~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_9),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[9] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N19
dffeas \exmem_if.rdat2_o[10] (
	.clk(CPUCLK),
	.d(\rdat2_o~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_10),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[10] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N25
dffeas \exmem_if.rdat2_o[11] (
	.clk(CPUCLK),
	.d(\rdat2_o~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_11),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[11] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N29
dffeas \exmem_if.rdat2_o[12] (
	.clk(CPUCLK),
	.d(\rdat2_o~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_12),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[12] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N3
dffeas \exmem_if.rdat2_o[13] (
	.clk(CPUCLK),
	.d(\rdat2_o~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_13),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[13] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N3
dffeas \exmem_if.rdat2_o[14] (
	.clk(CPUCLK),
	.d(\rdat2_o~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_14),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[14] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N25
dffeas \exmem_if.rdat2_o[15] (
	.clk(CPUCLK),
	.d(\rdat2_o~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_15),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[15] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N21
dffeas \exmem_if.rdat2_o[16] (
	.clk(CPUCLK),
	.d(\rdat2_o~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_16),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[16] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N5
dffeas \exmem_if.rdat2_o[17] (
	.clk(CPUCLK),
	.d(\rdat2_o~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_17),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[17] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N29
dffeas \exmem_if.rdat2_o[18] (
	.clk(CPUCLK),
	.d(\rdat2_o~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_18),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[18] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N15
dffeas \exmem_if.rdat2_o[19] (
	.clk(CPUCLK),
	.d(\rdat2_o~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_19),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[19] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N3
dffeas \exmem_if.rdat2_o[20] (
	.clk(CPUCLK),
	.d(\rdat2_o~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_20),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[20] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y34_N23
dffeas \exmem_if.rdat2_o[21] (
	.clk(CPUCLK),
	.d(\rdat2_o~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_21),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[21] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N27
dffeas \exmem_if.rdat2_o[22] (
	.clk(CPUCLK),
	.d(\rdat2_o~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_22),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[22] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N21
dffeas \exmem_if.rdat2_o[23] (
	.clk(CPUCLK),
	.d(\rdat2_o~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_23),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[23] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N1
dffeas \exmem_if.rdat2_o[24] (
	.clk(CPUCLK),
	.d(\rdat2_o~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_24),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[24] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N19
dffeas \exmem_if.rdat2_o[25] (
	.clk(CPUCLK),
	.d(\rdat2_o~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_25),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[25] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N25
dffeas \exmem_if.rdat2_o[26] (
	.clk(CPUCLK),
	.d(\rdat2_o~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_26),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[26] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N23
dffeas \exmem_if.rdat2_o[27] (
	.clk(CPUCLK),
	.d(\rdat2_o~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_27),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[27] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N15
dffeas \exmem_if.rdat2_o[28] (
	.clk(CPUCLK),
	.d(\rdat2_o~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_28),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[28] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N31
dffeas \exmem_if.rdat2_o[29] (
	.clk(CPUCLK),
	.d(\rdat2_o~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_29),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[29] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N17
dffeas \exmem_if.rdat2_o[30] (
	.clk(CPUCLK),
	.d(\rdat2_o~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_30),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[30] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N27
dffeas \exmem_if.rdat2_o[31] (
	.clk(CPUCLK),
	.d(\rdat2_o~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(exmem_ifrdat2_o_31),
	.prn(vcc));
// synopsys translate_off
defparam \exmem_if.rdat2_o[31] .is_wysiwyg = "true";
defparam \exmem_if.rdat2_o[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N0
cycloneive_lcell_comb \out_o~62 (
// Equation(s):
// \out_o~62_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & myifout_1))

	.dataa(exmem_ifdWEN_o),
	.datab(gnd),
	.datac(exmem_ifdREN_o),
	.datad(myifout_1),
	.cin(gnd),
	.combout(\out_o~62_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~62 .lut_mask = 16'h0500;
defparam \out_o~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N24
cycloneive_lcell_comb \dWEN_o~0 (
// Equation(s):
// \dWEN_o~0_combout  = (idex_ifdWEN_o & (!exmem_ifdWEN_o & !exmem_ifdREN_o))

	.dataa(idex_ifdWEN_o),
	.datab(exmem_ifdWEN_o),
	.datac(gnd),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\dWEN_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \dWEN_o~0 .lut_mask = 16'h0022;
defparam \dWEN_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N14
cycloneive_lcell_comb \dREN_o~0 (
// Equation(s):
// \dREN_o~0_combout  = (!exmem_ifdREN_o & (idex_ifdREN_o & !exmem_ifdWEN_o))

	.dataa(exmem_ifdREN_o),
	.datab(idex_ifdREN_o),
	.datac(gnd),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\dREN_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \dREN_o~0 .lut_mask = 16'h0044;
defparam \dREN_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N24
cycloneive_lcell_comb \out_o~63 (
// Equation(s):
// \out_o~63_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & myifout_0))

	.dataa(exmem_ifdWEN_o),
	.datab(gnd),
	.datac(exmem_ifdREN_o),
	.datad(myifout_0),
	.cin(gnd),
	.combout(\out_o~63_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~63 .lut_mask = 16'h0500;
defparam \out_o~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N16
cycloneive_lcell_comb \out_o~60 (
// Equation(s):
// \out_o~60_combout  = (always12 & ((myifout_32) # ((myifout_3 & myifout_31))))

	.dataa(myifout_3),
	.datab(myifout_32),
	.datac(myifout_31),
	.datad(always12),
	.cin(gnd),
	.combout(\out_o~60_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~60 .lut_mask = 16'hEC00;
defparam \out_o~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N16
cycloneive_lcell_comb \out_o~61 (
// Equation(s):
// \out_o~61_combout  = (always12 & ((myifout_2) # ((myifout_31 & myifout_210))))

	.dataa(myifout_31),
	.datab(always12),
	.datac(myifout_210),
	.datad(myifout_2),
	.cin(gnd),
	.combout(\out_o~61_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~61 .lut_mask = 16'hCC80;
defparam \out_o~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N30
cycloneive_lcell_comb \out_o~64 (
// Equation(s):
// \out_o~64_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & myifout_5))

	.dataa(exmem_ifdWEN_o),
	.datab(gnd),
	.datac(exmem_ifdREN_o),
	.datad(myifout_5),
	.cin(gnd),
	.combout(\out_o~64_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~64 .lut_mask = 16'h0500;
defparam \out_o~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N8
cycloneive_lcell_comb \out_o~65 (
// Equation(s):
// \out_o~65_combout  = (!exmem_ifdREN_o & (!exmem_ifdWEN_o & myifout_4))

	.dataa(gnd),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(myifout_4),
	.cin(gnd),
	.combout(\out_o~65_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~65 .lut_mask = 16'h0300;
defparam \out_o~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N16
cycloneive_lcell_comb \out_o~66 (
// Equation(s):
// \out_o~66_combout  = (!exmem_ifdREN_o & (myifout_7 & !exmem_ifdWEN_o))

	.dataa(exmem_ifdREN_o),
	.datab(gnd),
	.datac(myifout_7),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\out_o~66_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~66 .lut_mask = 16'h0050;
defparam \out_o~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N6
cycloneive_lcell_comb \out_o~67 (
// Equation(s):
// \out_o~67_combout  = (!exmem_ifdREN_o & (myifout_6 & !exmem_ifdWEN_o))

	.dataa(exmem_ifdREN_o),
	.datab(gnd),
	.datac(myifout_6),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\out_o~67_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~67 .lut_mask = 16'h0050;
defparam \out_o~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N26
cycloneive_lcell_comb \out_o~68 (
// Equation(s):
// \out_o~68_combout  = (!idex_ifaluop_o_3 & (!exmem_ifdREN_o & (!exmem_ifdWEN_o & myifout_9)))

	.dataa(idex_ifaluop_o_3),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(myifout_9),
	.cin(gnd),
	.combout(\out_o~68_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~68 .lut_mask = 16'h0100;
defparam \out_o~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N14
cycloneive_lcell_comb \out_o~69 (
// Equation(s):
// \out_o~69_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & (!idex_ifaluop_o_3 & myifout_8)))

	.dataa(exmem_ifdWEN_o),
	.datab(exmem_ifdREN_o),
	.datac(idex_ifaluop_o_3),
	.datad(myifout_8),
	.cin(gnd),
	.combout(\out_o~69_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~69 .lut_mask = 16'h0100;
defparam \out_o~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N6
cycloneive_lcell_comb \out_o~70 (
// Equation(s):
// \out_o~70_combout  = (!idex_ifaluop_o_3 & (!exmem_ifdWEN_o & (myifout_11 & !exmem_ifdREN_o)))

	.dataa(idex_ifaluop_o_3),
	.datab(exmem_ifdWEN_o),
	.datac(myifout_11),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\out_o~70_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~70 .lut_mask = 16'h0010;
defparam \out_o~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N22
cycloneive_lcell_comb \out_o~71 (
// Equation(s):
// \out_o~71_combout  = (!idex_ifaluop_o_3 & (!exmem_ifdREN_o & (!exmem_ifdWEN_o & myifout_10)))

	.dataa(idex_ifaluop_o_3),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(myifout_10),
	.cin(gnd),
	.combout(\out_o~71_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~71 .lut_mask = 16'h0100;
defparam \out_o~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N8
cycloneive_lcell_comb \out_o~72 (
// Equation(s):
// \out_o~72_combout  = (!idex_ifaluop_o_3 & (!exmem_ifdREN_o & (!exmem_ifdWEN_o & myifout_13)))

	.dataa(idex_ifaluop_o_3),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(myifout_13),
	.cin(gnd),
	.combout(\out_o~72_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~72 .lut_mask = 16'h0100;
defparam \out_o~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N14
cycloneive_lcell_comb \out_o~73 (
// Equation(s):
// \out_o~73_combout  = (!idex_ifaluop_o_3 & (myifout_12 & (!exmem_ifdWEN_o & !exmem_ifdREN_o)))

	.dataa(idex_ifaluop_o_3),
	.datab(myifout_12),
	.datac(exmem_ifdWEN_o),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\out_o~73_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~73 .lut_mask = 16'h0004;
defparam \out_o~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N16
cycloneive_lcell_comb \out_o~74 (
// Equation(s):
// \out_o~74_combout  = (!idex_ifaluop_o_3 & (!exmem_ifdREN_o & (!exmem_ifdWEN_o & myifout_15)))

	.dataa(idex_ifaluop_o_3),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(myifout_15),
	.cin(gnd),
	.combout(\out_o~74_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~74 .lut_mask = 16'h0100;
defparam \out_o~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N18
cycloneive_lcell_comb \out_o~75 (
// Equation(s):
// \out_o~75_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & (!idex_ifaluop_o_3 & myifout_14)))

	.dataa(exmem_ifdWEN_o),
	.datab(exmem_ifdREN_o),
	.datac(idex_ifaluop_o_3),
	.datad(myifout_14),
	.cin(gnd),
	.combout(\out_o~75_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~75 .lut_mask = 16'h0100;
defparam \out_o~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N20
cycloneive_lcell_comb \out_o~76 (
// Equation(s):
// \out_o~76_combout  = (!idex_ifaluop_o_3 & (!exmem_ifdREN_o & (!exmem_ifdWEN_o & myifout_17)))

	.dataa(idex_ifaluop_o_3),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(myifout_17),
	.cin(gnd),
	.combout(\out_o~76_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~76 .lut_mask = 16'h0100;
defparam \out_o~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N6
cycloneive_lcell_comb \out_o~77 (
// Equation(s):
// \out_o~77_combout  = (!exmem_ifdWEN_o & (!idex_ifaluop_o_3 & (!exmem_ifdREN_o & myifout_16)))

	.dataa(exmem_ifdWEN_o),
	.datab(idex_ifaluop_o_3),
	.datac(exmem_ifdREN_o),
	.datad(myifout_16),
	.cin(gnd),
	.combout(\out_o~77_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~77 .lut_mask = 16'h0100;
defparam \out_o~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N16
cycloneive_lcell_comb \out_o~78 (
// Equation(s):
// \out_o~78_combout  = (!idex_ifaluop_o_3 & (!exmem_ifdWEN_o & (myifout_19 & !exmem_ifdREN_o)))

	.dataa(idex_ifaluop_o_3),
	.datab(exmem_ifdWEN_o),
	.datac(myifout_19),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\out_o~78_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~78 .lut_mask = 16'h0010;
defparam \out_o~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N26
cycloneive_lcell_comb \out_o~79 (
// Equation(s):
// \out_o~79_combout  = (!idex_ifaluop_o_3 & (!exmem_ifdREN_o & (!exmem_ifdWEN_o & myifout_18)))

	.dataa(idex_ifaluop_o_3),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(myifout_18),
	.cin(gnd),
	.combout(\out_o~79_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~79 .lut_mask = 16'h0100;
defparam \out_o~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N22
cycloneive_lcell_comb \out_o~80 (
// Equation(s):
// \out_o~80_combout  = (!exmem_ifdREN_o & (!exmem_ifdWEN_o & (!idex_ifaluop_o_3 & myifout_21)))

	.dataa(exmem_ifdREN_o),
	.datab(exmem_ifdWEN_o),
	.datac(idex_ifaluop_o_3),
	.datad(myifout_21),
	.cin(gnd),
	.combout(\out_o~80_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~80 .lut_mask = 16'h0100;
defparam \out_o~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N6
cycloneive_lcell_comb \out_o~81 (
// Equation(s):
// \out_o~81_combout  = (!idex_ifaluop_o_3 & (!exmem_ifdREN_o & (myifout_20 & !exmem_ifdWEN_o)))

	.dataa(idex_ifaluop_o_3),
	.datab(exmem_ifdREN_o),
	.datac(myifout_20),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\out_o~81_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~81 .lut_mask = 16'h0010;
defparam \out_o~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N16
cycloneive_lcell_comb \out_o~82 (
// Equation(s):
// \out_o~82_combout  = (!exmem_ifdREN_o & (!idex_ifaluop_o_3 & (myifout_23 & !exmem_ifdWEN_o)))

	.dataa(exmem_ifdREN_o),
	.datab(idex_ifaluop_o_3),
	.datac(myifout_23),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\out_o~82_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~82 .lut_mask = 16'h0010;
defparam \out_o~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N12
cycloneive_lcell_comb \out_o~83 (
// Equation(s):
// \out_o~83_combout  = (!exmem_ifdREN_o & (!idex_ifaluop_o_3 & (myifout_22 & !exmem_ifdWEN_o)))

	.dataa(exmem_ifdREN_o),
	.datab(idex_ifaluop_o_3),
	.datac(myifout_22),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\out_o~83_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~83 .lut_mask = 16'h0010;
defparam \out_o~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N14
cycloneive_lcell_comb \out_o~84 (
// Equation(s):
// \out_o~84_combout  = (!exmem_ifdREN_o & (!exmem_ifdWEN_o & myifout_25))

	.dataa(exmem_ifdREN_o),
	.datab(gnd),
	.datac(exmem_ifdWEN_o),
	.datad(myifout_25),
	.cin(gnd),
	.combout(\out_o~84_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~84 .lut_mask = 16'h0500;
defparam \out_o~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N0
cycloneive_lcell_comb \out_o~85 (
// Equation(s):
// \out_o~85_combout  = (!exmem_ifdREN_o & (!exmem_ifdWEN_o & myifout_24))

	.dataa(gnd),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(myifout_24),
	.cin(gnd),
	.combout(\out_o~85_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~85 .lut_mask = 16'h0300;
defparam \out_o~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N28
cycloneive_lcell_comb \out_o~86 (
// Equation(s):
// \out_o~86_combout  = (!exmem_ifdREN_o & (!exmem_ifdWEN_o & myifout_27))

	.dataa(exmem_ifdREN_o),
	.datab(gnd),
	.datac(exmem_ifdWEN_o),
	.datad(myifout_27),
	.cin(gnd),
	.combout(\out_o~86_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~86 .lut_mask = 16'h0500;
defparam \out_o~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N28
cycloneive_lcell_comb \out_o~87 (
// Equation(s):
// \out_o~87_combout  = (myifout_26 & (!exmem_ifdWEN_o & !exmem_ifdREN_o))

	.dataa(myifout_26),
	.datab(gnd),
	.datac(exmem_ifdWEN_o),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\out_o~87_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~87 .lut_mask = 16'h000A;
defparam \out_o~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N8
cycloneive_lcell_comb \out_o~88 (
// Equation(s):
// \out_o~88_combout  = (!exmem_ifdREN_o & (!exmem_ifdWEN_o & myifout_29))

	.dataa(gnd),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(myifout_29),
	.cin(gnd),
	.combout(\out_o~88_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~88 .lut_mask = 16'h0300;
defparam \out_o~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N4
cycloneive_lcell_comb \out_o~89 (
// Equation(s):
// \out_o~89_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & myifout_28))

	.dataa(exmem_ifdWEN_o),
	.datab(exmem_ifdREN_o),
	.datac(myifout_28),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_o~89_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~89 .lut_mask = 16'h1010;
defparam \out_o~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N30
cycloneive_lcell_comb \out_o~90 (
// Equation(s):
// \out_o~90_combout  = (!idex_ifaluop_o_3 & (!exmem_ifdREN_o & (!exmem_ifdWEN_o & myifnegative)))

	.dataa(idex_ifaluop_o_3),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(myifnegative),
	.cin(gnd),
	.combout(\out_o~90_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~90 .lut_mask = 16'h0100;
defparam \out_o~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N4
cycloneive_lcell_comb \out_o~91 (
// Equation(s):
// \out_o~91_combout  = (!exmem_ifdREN_o & (!idex_ifaluop_o_3 & (myifout_30 & !exmem_ifdWEN_o)))

	.dataa(exmem_ifdREN_o),
	.datab(idex_ifaluop_o_3),
	.datac(myifout_30),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\out_o~91_combout ),
	.cout());
// synopsys translate_off
defparam \out_o~91 .lut_mask = 16'h0010;
defparam \out_o~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N28
cycloneive_lcell_comb \halt_o~0 (
// Equation(s):
// \halt_o~0_combout  = (idex_ifhalt_o & (!exmem_ifdWEN_o & !exmem_ifdREN_o))

	.dataa(idex_ifhalt_o),
	.datab(gnd),
	.datac(exmem_ifdWEN_o),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\halt_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \halt_o~0 .lut_mask = 16'h000A;
defparam \halt_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N0
cycloneive_lcell_comb \rdat2_o~0 (
// Equation(s):
// \rdat2_o~0_combout  = (always12 & ((fuifrdat2_ow & (fuifrtReplace_0)) # (!fuifrdat2_ow & ((idex_ifrdat2_o_0)))))

	.dataa(fuifrdat2_ow),
	.datab(always12),
	.datac(fuifrtReplace_0),
	.datad(idex_ifrdat2_o_0),
	.cin(gnd),
	.combout(\rdat2_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~0 .lut_mask = 16'hC480;
defparam \rdat2_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N18
cycloneive_lcell_comb \RegDest_o~0 (
// Equation(s):
// \RegDest_o~0_combout  = (idex_ifRegDest_o_1 & (!exmem_ifdREN_o & !exmem_ifdWEN_o))

	.dataa(idex_ifRegDest_o_1),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(gnd),
	.cin(gnd),
	.combout(\RegDest_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \RegDest_o~0 .lut_mask = 16'h0202;
defparam \RegDest_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N20
cycloneive_lcell_comb \rt_o~0 (
// Equation(s):
// \rt_o~0_combout  = (!exmem_ifdREN_o & (idex_ifrt_o_1 & !exmem_ifdWEN_o))

	.dataa(gnd),
	.datab(exmem_ifdREN_o),
	.datac(idex_ifrt_o_1),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\rt_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \rt_o~0 .lut_mask = 16'h0030;
defparam \rt_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N4
cycloneive_lcell_comb \rd_o~0 (
// Equation(s):
// \rd_o~0_combout  = (!exmem_ifdREN_o & (idex_ifrd_o_1 & !exmem_ifdWEN_o))

	.dataa(exmem_ifdREN_o),
	.datab(idex_ifrd_o_1),
	.datac(gnd),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\rd_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \rd_o~0 .lut_mask = 16'h0044;
defparam \rd_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N6
cycloneive_lcell_comb \RegDest_o~1 (
// Equation(s):
// \RegDest_o~1_combout  = (!exmem_ifdREN_o & (idex_ifRegDest_o_0 & !exmem_ifdWEN_o))

	.dataa(gnd),
	.datab(exmem_ifdREN_o),
	.datac(idex_ifRegDest_o_0),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\RegDest_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \RegDest_o~1 .lut_mask = 16'h0030;
defparam \RegDest_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N16
cycloneive_lcell_comb \rt_o~1 (
// Equation(s):
// \rt_o~1_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & idex_ifrt_o_0))

	.dataa(exmem_ifdWEN_o),
	.datab(exmem_ifdREN_o),
	.datac(gnd),
	.datad(idex_ifrt_o_0),
	.cin(gnd),
	.combout(\rt_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \rt_o~1 .lut_mask = 16'h1100;
defparam \rt_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N26
cycloneive_lcell_comb \rd_o~1 (
// Equation(s):
// \rd_o~1_combout  = (!exmem_ifdWEN_o & (idex_ifrd_o_0 & !exmem_ifdREN_o))

	.dataa(exmem_ifdWEN_o),
	.datab(gnd),
	.datac(idex_ifrd_o_0),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\rd_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \rd_o~1 .lut_mask = 16'h0050;
defparam \rd_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N22
cycloneive_lcell_comb \rt_o~2 (
// Equation(s):
// \rt_o~2_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & idex_ifrt_o_3))

	.dataa(exmem_ifdWEN_o),
	.datab(exmem_ifdREN_o),
	.datac(gnd),
	.datad(idex_ifrt_o_3),
	.cin(gnd),
	.combout(\rt_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \rt_o~2 .lut_mask = 16'h1100;
defparam \rt_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N12
cycloneive_lcell_comb \rd_o~2 (
// Equation(s):
// \rd_o~2_combout  = (!exmem_ifdWEN_o & (idex_ifrd_o_3 & !exmem_ifdREN_o))

	.dataa(exmem_ifdWEN_o),
	.datab(idex_ifrd_o_3),
	.datac(gnd),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\rd_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \rd_o~2 .lut_mask = 16'h0044;
defparam \rd_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N8
cycloneive_lcell_comb \rt_o~3 (
// Equation(s):
// \rt_o~3_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & idex_ifrt_o_2))

	.dataa(exmem_ifdWEN_o),
	.datab(exmem_ifdREN_o),
	.datac(gnd),
	.datad(idex_ifrt_o_2),
	.cin(gnd),
	.combout(\rt_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \rt_o~3 .lut_mask = 16'h1100;
defparam \rt_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N10
cycloneive_lcell_comb \rd_o~3 (
// Equation(s):
// \rd_o~3_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & idex_ifrd_o_2))

	.dataa(exmem_ifdWEN_o),
	.datab(exmem_ifdREN_o),
	.datac(gnd),
	.datad(idex_ifrd_o_2),
	.cin(gnd),
	.combout(\rd_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \rd_o~3 .lut_mask = 16'h1100;
defparam \rd_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N26
cycloneive_lcell_comb \regWEN_o~0 (
// Equation(s):
// \regWEN_o~0_combout  = (idex_ifregWEN_o & (!exmem_ifdREN_o & !exmem_ifdWEN_o))

	.dataa(idex_ifregWEN_o),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(gnd),
	.cin(gnd),
	.combout(\regWEN_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \regWEN_o~0 .lut_mask = 16'h0202;
defparam \regWEN_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N30
cycloneive_lcell_comb \rt_o~4 (
// Equation(s):
// \rt_o~4_combout  = (!exmem_ifdREN_o & (!exmem_ifdWEN_o & idex_ifrt_o_4))

	.dataa(gnd),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(idex_ifrt_o_4),
	.cin(gnd),
	.combout(\rt_o~4_combout ),
	.cout());
// synopsys translate_off
defparam \rt_o~4 .lut_mask = 16'h0300;
defparam \rt_o~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N8
cycloneive_lcell_comb \rd_o~4 (
// Equation(s):
// \rd_o~4_combout  = (!exmem_ifdREN_o & (idex_ifrd_o_4 & !exmem_ifdWEN_o))

	.dataa(exmem_ifdREN_o),
	.datab(gnd),
	.datac(idex_ifrd_o_4),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\rd_o~4_combout ),
	.cout());
// synopsys translate_off
defparam \rd_o~4 .lut_mask = 16'h0050;
defparam \rd_o~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N16
cycloneive_lcell_comb \jal_o~0 (
// Equation(s):
// \jal_o~0_combout  = (idex_ifjal_o & (!exmem_ifdREN_o & !exmem_ifdWEN_o))

	.dataa(idex_ifjal_o),
	.datab(exmem_ifdREN_o),
	.datac(gnd),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\jal_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \jal_o~0 .lut_mask = 16'h0022;
defparam \jal_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N26
cycloneive_lcell_comb \lui_o~0 (
// Equation(s):
// \lui_o~0_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & idex_iflui_o))

	.dataa(exmem_ifdWEN_o),
	.datab(exmem_ifdREN_o),
	.datac(idex_iflui_o),
	.datad(gnd),
	.cin(gnd),
	.combout(\lui_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \lui_o~0 .lut_mask = 16'h1010;
defparam \lui_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N18
cycloneive_lcell_comb \next_pc_o~0 (
// Equation(s):
// \next_pc_o~0_combout  = (!exmem_ifdREN_o & (!exmem_ifdWEN_o & idex_ifnext_pc_o_1))

	.dataa(exmem_ifdREN_o),
	.datab(exmem_ifdWEN_o),
	.datac(gnd),
	.datad(idex_ifnext_pc_o_1),
	.cin(gnd),
	.combout(\next_pc_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~0 .lut_mask = 16'h1100;
defparam \next_pc_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N8
cycloneive_lcell_comb \memToReg_o~0 (
// Equation(s):
// \memToReg_o~0_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & idex_ifmemToReg_o))

	.dataa(exmem_ifdWEN_o),
	.datab(gnd),
	.datac(exmem_ifdREN_o),
	.datad(idex_ifmemToReg_o),
	.cin(gnd),
	.combout(\memToReg_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \memToReg_o~0 .lut_mask = 16'h0500;
defparam \memToReg_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N22
cycloneive_lcell_comb \next_pc_o~1 (
// Equation(s):
// \next_pc_o~1_combout  = (!exmem_ifdREN_o & (!exmem_ifdWEN_o & idex_ifnext_pc_o_0))

	.dataa(exmem_ifdREN_o),
	.datab(exmem_ifdWEN_o),
	.datac(gnd),
	.datad(idex_ifnext_pc_o_0),
	.cin(gnd),
	.combout(\next_pc_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~1 .lut_mask = 16'h1100;
defparam \next_pc_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N28
cycloneive_lcell_comb \next_pc_o~2 (
// Equation(s):
// \next_pc_o~2_combout  = (!exmem_ifdREN_o & (idex_ifnext_pc_o_2 & !exmem_ifdWEN_o))

	.dataa(exmem_ifdREN_o),
	.datab(idex_ifnext_pc_o_2),
	.datac(gnd),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\next_pc_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~2 .lut_mask = 16'h0044;
defparam \next_pc_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N16
cycloneive_lcell_comb \next_pc_o~3 (
// Equation(s):
// \next_pc_o~3_combout  = (!exmem_ifdWEN_o & (idex_ifnext_pc_o_4 & !exmem_ifdREN_o))

	.dataa(gnd),
	.datab(exmem_ifdWEN_o),
	.datac(idex_ifnext_pc_o_4),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\next_pc_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~3 .lut_mask = 16'h0030;
defparam \next_pc_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N4
cycloneive_lcell_comb \exmem_if.next_pc_o[4]~feeder (
// Equation(s):
// \exmem_if.next_pc_o[4]~feeder_combout  = \next_pc_o~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\next_pc_o~3_combout ),
	.cin(gnd),
	.combout(\exmem_if.next_pc_o[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \exmem_if.next_pc_o[4]~feeder .lut_mask = 16'hFF00;
defparam \exmem_if.next_pc_o[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N12
cycloneive_lcell_comb \next_pc_o~4 (
// Equation(s):
// \next_pc_o~4_combout  = (!exmem_ifdREN_o & (idex_ifnext_pc_o_3 & !exmem_ifdWEN_o))

	.dataa(exmem_ifdREN_o),
	.datab(idex_ifnext_pc_o_3),
	.datac(gnd),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\next_pc_o~4_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~4 .lut_mask = 16'h0044;
defparam \next_pc_o~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N26
cycloneive_lcell_comb \next_pc_o~5 (
// Equation(s):
// \next_pc_o~5_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & idex_ifnext_pc_o_8))

	.dataa(exmem_ifdWEN_o),
	.datab(exmem_ifdREN_o),
	.datac(gnd),
	.datad(idex_ifnext_pc_o_8),
	.cin(gnd),
	.combout(\next_pc_o~5_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~5 .lut_mask = 16'h1100;
defparam \next_pc_o~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N8
cycloneive_lcell_comb \next_pc_o~6 (
// Equation(s):
// \next_pc_o~6_combout  = (!exmem_ifdREN_o & (idex_ifnext_pc_o_7 & !exmem_ifdWEN_o))

	.dataa(exmem_ifdREN_o),
	.datab(idex_ifnext_pc_o_7),
	.datac(gnd),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\next_pc_o~6_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~6 .lut_mask = 16'h0044;
defparam \next_pc_o~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N30
cycloneive_lcell_comb \next_pc_o~7 (
// Equation(s):
// \next_pc_o~7_combout  = (!exmem_ifdWEN_o & (idex_ifnext_pc_o_6 & !exmem_ifdREN_o))

	.dataa(exmem_ifdWEN_o),
	.datab(idex_ifnext_pc_o_6),
	.datac(gnd),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\next_pc_o~7_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~7 .lut_mask = 16'h0044;
defparam \next_pc_o~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N20
cycloneive_lcell_comb \next_pc_o~8 (
// Equation(s):
// \next_pc_o~8_combout  = (idex_ifnext_pc_o_5 & (!exmem_ifdREN_o & !exmem_ifdWEN_o))

	.dataa(idex_ifnext_pc_o_5),
	.datab(exmem_ifdREN_o),
	.datac(gnd),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\next_pc_o~8_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~8 .lut_mask = 16'h0022;
defparam \next_pc_o~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N18
cycloneive_lcell_comb \imm_o~0 (
// Equation(s):
// \imm_o~0_combout  = (!exmem_ifdREN_o & (!exmem_ifdWEN_o & idex_ifimm_o_0))

	.dataa(exmem_ifdREN_o),
	.datab(exmem_ifdWEN_o),
	.datac(gnd),
	.datad(idex_ifimm_o_0),
	.cin(gnd),
	.combout(\imm_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~0 .lut_mask = 16'h1100;
defparam \imm_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N0
cycloneive_lcell_comb \next_pc_o~9 (
// Equation(s):
// \next_pc_o~9_combout  = (idex_ifnext_pc_o_16 & (!exmem_ifdREN_o & !exmem_ifdWEN_o))

	.dataa(gnd),
	.datab(idex_ifnext_pc_o_16),
	.datac(exmem_ifdREN_o),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\next_pc_o~9_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~9 .lut_mask = 16'h000C;
defparam \next_pc_o~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N20
cycloneive_lcell_comb \next_pc_o~10 (
// Equation(s):
// \next_pc_o~10_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & idex_ifnext_pc_o_15))

	.dataa(exmem_ifdWEN_o),
	.datab(exmem_ifdREN_o),
	.datac(gnd),
	.datad(idex_ifnext_pc_o_15),
	.cin(gnd),
	.combout(\next_pc_o~10_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~10 .lut_mask = 16'h1100;
defparam \next_pc_o~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N30
cycloneive_lcell_comb \next_pc_o~11 (
// Equation(s):
// \next_pc_o~11_combout  = (!exmem_ifdREN_o & (idex_ifnext_pc_o_14 & !exmem_ifdWEN_o))

	.dataa(gnd),
	.datab(exmem_ifdREN_o),
	.datac(idex_ifnext_pc_o_14),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\next_pc_o~11_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~11 .lut_mask = 16'h0030;
defparam \next_pc_o~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N14
cycloneive_lcell_comb \next_pc_o~12 (
// Equation(s):
// \next_pc_o~12_combout  = (!exmem_ifdREN_o & (idex_ifnext_pc_o_13 & !exmem_ifdWEN_o))

	.dataa(exmem_ifdREN_o),
	.datab(idex_ifnext_pc_o_13),
	.datac(exmem_ifdWEN_o),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pc_o~12_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~12 .lut_mask = 16'h0404;
defparam \next_pc_o~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N4
cycloneive_lcell_comb \next_pc_o~13 (
// Equation(s):
// \next_pc_o~13_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & idex_ifnext_pc_o_12))

	.dataa(exmem_ifdWEN_o),
	.datab(gnd),
	.datac(exmem_ifdREN_o),
	.datad(idex_ifnext_pc_o_12),
	.cin(gnd),
	.combout(\next_pc_o~13_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~13 .lut_mask = 16'h0500;
defparam \next_pc_o~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N16
cycloneive_lcell_comb \next_pc_o~14 (
// Equation(s):
// \next_pc_o~14_combout  = (!exmem_ifdREN_o & (idex_ifnext_pc_o_11 & !exmem_ifdWEN_o))

	.dataa(exmem_ifdREN_o),
	.datab(gnd),
	.datac(idex_ifnext_pc_o_11),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\next_pc_o~14_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~14 .lut_mask = 16'h0050;
defparam \next_pc_o~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N10
cycloneive_lcell_comb \next_pc_o~15 (
// Equation(s):
// \next_pc_o~15_combout  = (idex_ifnext_pc_o_10 & (!exmem_ifdREN_o & !exmem_ifdWEN_o))

	.dataa(gnd),
	.datab(idex_ifnext_pc_o_10),
	.datac(exmem_ifdREN_o),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\next_pc_o~15_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~15 .lut_mask = 16'h000C;
defparam \next_pc_o~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N30
cycloneive_lcell_comb \next_pc_o~16 (
// Equation(s):
// \next_pc_o~16_combout  = (!exmem_ifdREN_o & (idex_ifnext_pc_o_9 & !exmem_ifdWEN_o))

	.dataa(exmem_ifdREN_o),
	.datab(idex_ifnext_pc_o_9),
	.datac(exmem_ifdWEN_o),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pc_o~16_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~16 .lut_mask = 16'h0404;
defparam \next_pc_o~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N24
cycloneive_lcell_comb \next_pc_o~17 (
// Equation(s):
// \next_pc_o~17_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & idex_ifnext_pc_o_31))

	.dataa(exmem_ifdWEN_o),
	.datab(exmem_ifdREN_o),
	.datac(idex_ifnext_pc_o_31),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pc_o~17_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~17 .lut_mask = 16'h1010;
defparam \next_pc_o~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N14
cycloneive_lcell_comb \imm_o~1 (
// Equation(s):
// \imm_o~1_combout  = (!exmem_ifdWEN_o & (idex_ifimm_o_15 & !exmem_ifdREN_o))

	.dataa(exmem_ifdWEN_o),
	.datab(idex_ifimm_o_15),
	.datac(exmem_ifdREN_o),
	.datad(gnd),
	.cin(gnd),
	.combout(\imm_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~1 .lut_mask = 16'h0404;
defparam \imm_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N22
cycloneive_lcell_comb \next_pc_o~18 (
// Equation(s):
// \next_pc_o~18_combout  = (idex_ifnext_pc_o_29 & (!exmem_ifdREN_o & !exmem_ifdWEN_o))

	.dataa(idex_ifnext_pc_o_29),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pc_o~18_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~18 .lut_mask = 16'h0202;
defparam \next_pc_o~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N20
cycloneive_lcell_comb \imm_o~2 (
// Equation(s):
// \imm_o~2_combout  = (idex_ifimm_o_13 & (!exmem_ifdREN_o & !exmem_ifdWEN_o))

	.dataa(idex_ifimm_o_13),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(gnd),
	.cin(gnd),
	.combout(\imm_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~2 .lut_mask = 16'h0202;
defparam \imm_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N30
cycloneive_lcell_comb \imm_o~3 (
// Equation(s):
// \imm_o~3_combout  = (!exmem_ifdWEN_o & (idex_ifimm_o_14 & !exmem_ifdREN_o))

	.dataa(exmem_ifdWEN_o),
	.datab(idex_ifimm_o_14),
	.datac(gnd),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\imm_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~3 .lut_mask = 16'h0044;
defparam \imm_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N14
cycloneive_lcell_comb \next_pc_o~19 (
// Equation(s):
// \next_pc_o~19_combout  = (idex_ifnext_pc_o_30 & (!exmem_ifdWEN_o & !exmem_ifdREN_o))

	.dataa(gnd),
	.datab(idex_ifnext_pc_o_30),
	.datac(exmem_ifdWEN_o),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\next_pc_o~19_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~19 .lut_mask = 16'h000C;
defparam \next_pc_o~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N22
cycloneive_lcell_comb \imm_o~4 (
// Equation(s):
// \imm_o~4_combout  = (idex_ifimm_o_12 & (!exmem_ifdWEN_o & !exmem_ifdREN_o))

	.dataa(idex_ifimm_o_12),
	.datab(gnd),
	.datac(exmem_ifdWEN_o),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\imm_o~4_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~4 .lut_mask = 16'h000A;
defparam \imm_o~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N26
cycloneive_lcell_comb \next_pc_o~20 (
// Equation(s):
// \next_pc_o~20_combout  = (idex_ifnext_pc_o_28 & (!exmem_ifdREN_o & !exmem_ifdWEN_o))

	.dataa(idex_ifnext_pc_o_28),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pc_o~20_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~20 .lut_mask = 16'h0202;
defparam \next_pc_o~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N12
cycloneive_lcell_comb \imm_o~5 (
// Equation(s):
// \imm_o~5_combout  = (!exmem_ifdREN_o & (!exmem_ifdWEN_o & idex_ifimm_o_10))

	.dataa(exmem_ifdREN_o),
	.datab(exmem_ifdWEN_o),
	.datac(gnd),
	.datad(idex_ifimm_o_10),
	.cin(gnd),
	.combout(\imm_o~5_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~5 .lut_mask = 16'h1100;
defparam \imm_o~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N6
cycloneive_lcell_comb \next_pc_o~21 (
// Equation(s):
// \next_pc_o~21_combout  = (!exmem_ifdREN_o & (idex_ifnext_pc_o_26 & !exmem_ifdWEN_o))

	.dataa(exmem_ifdREN_o),
	.datab(gnd),
	.datac(idex_ifnext_pc_o_26),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\next_pc_o~21_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~21 .lut_mask = 16'h0050;
defparam \next_pc_o~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N4
cycloneive_lcell_comb \next_pc_o~22 (
// Equation(s):
// \next_pc_o~22_combout  = (!exmem_ifdREN_o & (!exmem_ifdWEN_o & idex_ifnext_pc_o_27))

	.dataa(exmem_ifdREN_o),
	.datab(gnd),
	.datac(exmem_ifdWEN_o),
	.datad(idex_ifnext_pc_o_27),
	.cin(gnd),
	.combout(\next_pc_o~22_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~22 .lut_mask = 16'h0500;
defparam \next_pc_o~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N0
cycloneive_lcell_comb \imm_o~6 (
// Equation(s):
// \imm_o~6_combout  = (idex_ifimm_o_11 & (!exmem_ifdREN_o & !exmem_ifdWEN_o))

	.dataa(idex_ifimm_o_11),
	.datab(exmem_ifdREN_o),
	.datac(gnd),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\imm_o~6_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~6 .lut_mask = 16'h0022;
defparam \imm_o~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N30
cycloneive_lcell_comb \next_pc_o~23 (
// Equation(s):
// \next_pc_o~23_combout  = (idex_ifnext_pc_o_25 & (!exmem_ifdWEN_o & !exmem_ifdREN_o))

	.dataa(idex_ifnext_pc_o_25),
	.datab(exmem_ifdWEN_o),
	.datac(gnd),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\next_pc_o~23_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~23 .lut_mask = 16'h0022;
defparam \next_pc_o~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N12
cycloneive_lcell_comb \imm_o~7 (
// Equation(s):
// \imm_o~7_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & idex_ifimm_o_9))

	.dataa(exmem_ifdWEN_o),
	.datab(exmem_ifdREN_o),
	.datac(idex_ifimm_o_9),
	.datad(gnd),
	.cin(gnd),
	.combout(\imm_o~7_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~7 .lut_mask = 16'h1010;
defparam \imm_o~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N20
cycloneive_lcell_comb \imm_o~8 (
// Equation(s):
// \imm_o~8_combout  = (idex_ifimm_o_8 & (!exmem_ifdWEN_o & !exmem_ifdREN_o))

	.dataa(idex_ifimm_o_8),
	.datab(exmem_ifdWEN_o),
	.datac(gnd),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\imm_o~8_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~8 .lut_mask = 16'h0022;
defparam \imm_o~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N20
cycloneive_lcell_comb \next_pc_o~24 (
// Equation(s):
// \next_pc_o~24_combout  = (idex_ifnext_pc_o_24 & (!exmem_ifdWEN_o & !exmem_ifdREN_o))

	.dataa(idex_ifnext_pc_o_24),
	.datab(exmem_ifdWEN_o),
	.datac(gnd),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\next_pc_o~24_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~24 .lut_mask = 16'h0022;
defparam \next_pc_o~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N22
cycloneive_lcell_comb \imm_o~9 (
// Equation(s):
// \imm_o~9_combout  = (!exmem_ifdREN_o & (idex_ifimm_o_6 & !exmem_ifdWEN_o))

	.dataa(gnd),
	.datab(exmem_ifdREN_o),
	.datac(idex_ifimm_o_6),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\imm_o~9_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~9 .lut_mask = 16'h0030;
defparam \imm_o~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N22
cycloneive_lcell_comb \next_pc_o~25 (
// Equation(s):
// \next_pc_o~25_combout  = (idex_ifnext_pc_o_22 & (!exmem_ifdWEN_o & !exmem_ifdREN_o))

	.dataa(idex_ifnext_pc_o_22),
	.datab(gnd),
	.datac(exmem_ifdWEN_o),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\next_pc_o~25_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~25 .lut_mask = 16'h000A;
defparam \next_pc_o~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N4
cycloneive_lcell_comb \next_pc_o~26 (
// Equation(s):
// \next_pc_o~26_combout  = (!exmem_ifdREN_o & (idex_ifnext_pc_o_23 & !exmem_ifdWEN_o))

	.dataa(exmem_ifdREN_o),
	.datab(idex_ifnext_pc_o_23),
	.datac(gnd),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\next_pc_o~26_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~26 .lut_mask = 16'h0044;
defparam \next_pc_o~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N24
cycloneive_lcell_comb \imm_o~10 (
// Equation(s):
// \imm_o~10_combout  = (idex_ifimm_o_7 & (!exmem_ifdWEN_o & !exmem_ifdREN_o))

	.dataa(gnd),
	.datab(idex_ifimm_o_7),
	.datac(exmem_ifdWEN_o),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\imm_o~10_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~10 .lut_mask = 16'h000C;
defparam \imm_o~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N10
cycloneive_lcell_comb \next_pc_o~27 (
// Equation(s):
// \next_pc_o~27_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & idex_ifnext_pc_o_21))

	.dataa(exmem_ifdWEN_o),
	.datab(exmem_ifdREN_o),
	.datac(gnd),
	.datad(idex_ifnext_pc_o_21),
	.cin(gnd),
	.combout(\next_pc_o~27_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~27 .lut_mask = 16'h1100;
defparam \next_pc_o~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N12
cycloneive_lcell_comb \exmem_if.next_pc_o[21]~feeder (
// Equation(s):
// \exmem_if.next_pc_o[21]~feeder_combout  = \next_pc_o~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\next_pc_o~27_combout ),
	.cin(gnd),
	.combout(\exmem_if.next_pc_o[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \exmem_if.next_pc_o[21]~feeder .lut_mask = 16'hFF00;
defparam \exmem_if.next_pc_o[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N28
cycloneive_lcell_comb \imm_o~11 (
// Equation(s):
// \imm_o~11_combout  = (!exmem_ifdREN_o & (idex_ifimm_o_5 & !exmem_ifdWEN_o))

	.dataa(exmem_ifdREN_o),
	.datab(idex_ifimm_o_5),
	.datac(gnd),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\imm_o~11_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~11 .lut_mask = 16'h0044;
defparam \imm_o~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N18
cycloneive_lcell_comb \imm_o~12 (
// Equation(s):
// \imm_o~12_combout  = (idex_ifimm_o_4 & (!exmem_ifdWEN_o & !exmem_ifdREN_o))

	.dataa(idex_ifimm_o_4),
	.datab(exmem_ifdWEN_o),
	.datac(gnd),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\imm_o~12_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~12 .lut_mask = 16'h0022;
defparam \imm_o~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N12
cycloneive_lcell_comb \next_pc_o~28 (
// Equation(s):
// \next_pc_o~28_combout  = (idex_ifnext_pc_o_20 & (!exmem_ifdWEN_o & !exmem_ifdREN_o))

	.dataa(idex_ifnext_pc_o_20),
	.datab(exmem_ifdWEN_o),
	.datac(gnd),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\next_pc_o~28_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~28 .lut_mask = 16'h0022;
defparam \next_pc_o~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N4
cycloneive_lcell_comb \imm_o~13 (
// Equation(s):
// \imm_o~13_combout  = (!exmem_ifdREN_o & (idex_ifimm_o_2 & !exmem_ifdWEN_o))

	.dataa(gnd),
	.datab(exmem_ifdREN_o),
	.datac(idex_ifimm_o_2),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\imm_o~13_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~13 .lut_mask = 16'h0030;
defparam \imm_o~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N18
cycloneive_lcell_comb \next_pc_o~29 (
// Equation(s):
// \next_pc_o~29_combout  = (idex_ifnext_pc_o_18 & (!exmem_ifdREN_o & !exmem_ifdWEN_o))

	.dataa(idex_ifnext_pc_o_18),
	.datab(exmem_ifdREN_o),
	.datac(gnd),
	.datad(exmem_ifdWEN_o),
	.cin(gnd),
	.combout(\next_pc_o~29_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~29 .lut_mask = 16'h0022;
defparam \next_pc_o~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N28
cycloneive_lcell_comb \next_pc_o~30 (
// Equation(s):
// \next_pc_o~30_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & idex_ifnext_pc_o_19))

	.dataa(exmem_ifdWEN_o),
	.datab(exmem_ifdREN_o),
	.datac(idex_ifnext_pc_o_19),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pc_o~30_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~30 .lut_mask = 16'h1010;
defparam \next_pc_o~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N30
cycloneive_lcell_comb \imm_o~14 (
// Equation(s):
// \imm_o~14_combout  = (idex_ifimm_o_3 & (!exmem_ifdWEN_o & !exmem_ifdREN_o))

	.dataa(idex_ifimm_o_3),
	.datab(gnd),
	.datac(exmem_ifdWEN_o),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\imm_o~14_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~14 .lut_mask = 16'h000A;
defparam \imm_o~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N10
cycloneive_lcell_comb \next_pc_o~31 (
// Equation(s):
// \next_pc_o~31_combout  = (!exmem_ifdWEN_o & (idex_ifnext_pc_o_17 & !exmem_ifdREN_o))

	.dataa(gnd),
	.datab(exmem_ifdWEN_o),
	.datac(idex_ifnext_pc_o_17),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\next_pc_o~31_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~31 .lut_mask = 16'h0030;
defparam \next_pc_o~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N24
cycloneive_lcell_comb \imm_o~15 (
// Equation(s):
// \imm_o~15_combout  = (!exmem_ifdWEN_o & (!exmem_ifdREN_o & idex_ifimm_o_1))

	.dataa(exmem_ifdWEN_o),
	.datab(exmem_ifdREN_o),
	.datac(gnd),
	.datad(idex_ifimm_o_1),
	.cin(gnd),
	.combout(\imm_o~15_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~15 .lut_mask = 16'h1100;
defparam \imm_o~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N10
cycloneive_lcell_comb \rdat2_o~1 (
// Equation(s):
// \rdat2_o~1_combout  = (always12 & ((fuifrdat2_ow & ((fuifrtReplace_1))) # (!fuifrdat2_ow & (idex_ifrdat2_o_1))))

	.dataa(always12),
	.datab(idex_ifrdat2_o_1),
	.datac(fuifrtReplace_1),
	.datad(fuifrdat2_ow),
	.cin(gnd),
	.combout(\rdat2_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~1 .lut_mask = 16'hA088;
defparam \rdat2_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N6
cycloneive_lcell_comb \rdat2_o~2 (
// Equation(s):
// \rdat2_o~2_combout  = (always12 & ((fuifrdat2_ow & ((fuifrtReplace_2))) # (!fuifrdat2_ow & (idex_ifrdat2_o_2))))

	.dataa(always12),
	.datab(idex_ifrdat2_o_2),
	.datac(fuifrtReplace_2),
	.datad(fuifrdat2_ow),
	.cin(gnd),
	.combout(\rdat2_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~2 .lut_mask = 16'hA088;
defparam \rdat2_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N18
cycloneive_lcell_comb \rdat2_o~3 (
// Equation(s):
// \rdat2_o~3_combout  = (always12 & ((fuifrdat2_ow & (fuifrtReplace_3)) # (!fuifrdat2_ow & ((idex_ifrdat2_o_3)))))

	.dataa(fuifrdat2_ow),
	.datab(fuifrtReplace_3),
	.datac(always12),
	.datad(idex_ifrdat2_o_3),
	.cin(gnd),
	.combout(\rdat2_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~3 .lut_mask = 16'hD080;
defparam \rdat2_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N12
cycloneive_lcell_comb \rdat2_o~4 (
// Equation(s):
// \rdat2_o~4_combout  = (always12 & ((fuifrdat2_ow & (fuifrtReplace_4)) # (!fuifrdat2_ow & ((idex_ifrdat2_o_4)))))

	.dataa(fuifrtReplace_4),
	.datab(always12),
	.datac(fuifrdat2_ow),
	.datad(idex_ifrdat2_o_4),
	.cin(gnd),
	.combout(\rdat2_o~4_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~4 .lut_mask = 16'h8C80;
defparam \rdat2_o~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N20
cycloneive_lcell_comb \rdat2_o~5 (
// Equation(s):
// \rdat2_o~5_combout  = (always12 & ((fuifrdat2_ow & (fuifrtReplace_5)) # (!fuifrdat2_ow & ((idex_ifrdat2_o_5)))))

	.dataa(fuifrdat2_ow),
	.datab(fuifrtReplace_5),
	.datac(idex_ifrdat2_o_5),
	.datad(always12),
	.cin(gnd),
	.combout(\rdat2_o~5_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~5 .lut_mask = 16'hD800;
defparam \rdat2_o~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N0
cycloneive_lcell_comb \rdat2_o~6 (
// Equation(s):
// \rdat2_o~6_combout  = (always12 & ((fuifrdat2_ow & ((fuifrtReplace_6))) # (!fuifrdat2_ow & (idex_ifrdat2_o_6))))

	.dataa(fuifrdat2_ow),
	.datab(always12),
	.datac(idex_ifrdat2_o_6),
	.datad(fuifrtReplace_6),
	.cin(gnd),
	.combout(\rdat2_o~6_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~6 .lut_mask = 16'hC840;
defparam \rdat2_o~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N18
cycloneive_lcell_comb \rdat2_o~7 (
// Equation(s):
// \rdat2_o~7_combout  = (always12 & ((fuifrdat2_ow & ((fuifrtReplace_7))) # (!fuifrdat2_ow & (idex_ifrdat2_o_7))))

	.dataa(idex_ifrdat2_o_7),
	.datab(fuifrtReplace_7),
	.datac(fuifrdat2_ow),
	.datad(always12),
	.cin(gnd),
	.combout(\rdat2_o~7_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~7 .lut_mask = 16'hCA00;
defparam \rdat2_o~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N26
cycloneive_lcell_comb \rdat2_o~8 (
// Equation(s):
// \rdat2_o~8_combout  = (always12 & ((fuifrdat2_ow & ((fuifrtReplace_8))) # (!fuifrdat2_ow & (idex_ifrdat2_o_8))))

	.dataa(idex_ifrdat2_o_8),
	.datab(fuifrtReplace_8),
	.datac(always12),
	.datad(fuifrdat2_ow),
	.cin(gnd),
	.combout(\rdat2_o~8_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~8 .lut_mask = 16'hC0A0;
defparam \rdat2_o~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N28
cycloneive_lcell_comb \rdat2_o~9 (
// Equation(s):
// \rdat2_o~9_combout  = (always12 & ((fuifrdat2_ow & ((fuifrtReplace_9))) # (!fuifrdat2_ow & (idex_ifrdat2_o_9))))

	.dataa(fuifrdat2_ow),
	.datab(idex_ifrdat2_o_9),
	.datac(always12),
	.datad(fuifrtReplace_9),
	.cin(gnd),
	.combout(\rdat2_o~9_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~9 .lut_mask = 16'hE040;
defparam \rdat2_o~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N18
cycloneive_lcell_comb \rdat2_o~10 (
// Equation(s):
// \rdat2_o~10_combout  = (always12 & ((fuifrdat2_ow & (fuifrtReplace_10)) # (!fuifrdat2_ow & ((idex_ifrdat2_o_10)))))

	.dataa(fuifrtReplace_10),
	.datab(fuifrdat2_ow),
	.datac(always12),
	.datad(idex_ifrdat2_o_10),
	.cin(gnd),
	.combout(\rdat2_o~10_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~10 .lut_mask = 16'hB080;
defparam \rdat2_o~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N24
cycloneive_lcell_comb \rdat2_o~11 (
// Equation(s):
// \rdat2_o~11_combout  = (always12 & ((fuifrdat2_ow & (fuifrtReplace_11)) # (!fuifrdat2_ow & ((idex_ifrdat2_o_11)))))

	.dataa(fuifrdat2_ow),
	.datab(fuifrtReplace_11),
	.datac(always12),
	.datad(idex_ifrdat2_o_11),
	.cin(gnd),
	.combout(\rdat2_o~11_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~11 .lut_mask = 16'hD080;
defparam \rdat2_o~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N28
cycloneive_lcell_comb \rdat2_o~12 (
// Equation(s):
// \rdat2_o~12_combout  = (always12 & ((fuifrdat2_ow & ((fuifrtReplace_12))) # (!fuifrdat2_ow & (idex_ifrdat2_o_12))))

	.dataa(always12),
	.datab(idex_ifrdat2_o_12),
	.datac(fuifrdat2_ow),
	.datad(fuifrtReplace_12),
	.cin(gnd),
	.combout(\rdat2_o~12_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~12 .lut_mask = 16'hA808;
defparam \rdat2_o~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N2
cycloneive_lcell_comb \rdat2_o~13 (
// Equation(s):
// \rdat2_o~13_combout  = (always12 & ((fuifrdat2_ow & (fuifrtReplace_13)) # (!fuifrdat2_ow & ((idex_ifrdat2_o_13)))))

	.dataa(fuifrdat2_ow),
	.datab(fuifrtReplace_13),
	.datac(always12),
	.datad(idex_ifrdat2_o_13),
	.cin(gnd),
	.combout(\rdat2_o~13_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~13 .lut_mask = 16'hD080;
defparam \rdat2_o~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N2
cycloneive_lcell_comb \rdat2_o~14 (
// Equation(s):
// \rdat2_o~14_combout  = (always12 & ((fuifrdat2_ow & (fuifrtReplace_14)) # (!fuifrdat2_ow & ((idex_ifrdat2_o_14)))))

	.dataa(fuifrdat2_ow),
	.datab(fuifrtReplace_14),
	.datac(always12),
	.datad(idex_ifrdat2_o_14),
	.cin(gnd),
	.combout(\rdat2_o~14_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~14 .lut_mask = 16'hD080;
defparam \rdat2_o~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N24
cycloneive_lcell_comb \rdat2_o~15 (
// Equation(s):
// \rdat2_o~15_combout  = (always12 & ((fuifrdat2_ow & (fuifrtReplace_15)) # (!fuifrdat2_ow & ((idex_ifrdat2_o_15)))))

	.dataa(fuifrtReplace_15),
	.datab(always12),
	.datac(idex_ifrdat2_o_15),
	.datad(fuifrdat2_ow),
	.cin(gnd),
	.combout(\rdat2_o~15_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~15 .lut_mask = 16'h88C0;
defparam \rdat2_o~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N20
cycloneive_lcell_comb \rdat2_o~16 (
// Equation(s):
// \rdat2_o~16_combout  = (always12 & ((fuifrdat2_ow & ((fuifrtReplace_16))) # (!fuifrdat2_ow & (idex_ifrdat2_o_16))))

	.dataa(idex_ifrdat2_o_16),
	.datab(always12),
	.datac(fuifrdat2_ow),
	.datad(fuifrtReplace_16),
	.cin(gnd),
	.combout(\rdat2_o~16_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~16 .lut_mask = 16'hC808;
defparam \rdat2_o~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N4
cycloneive_lcell_comb \rdat2_o~17 (
// Equation(s):
// \rdat2_o~17_combout  = (always12 & ((fuifrdat2_ow & ((fuifrtReplace_17))) # (!fuifrdat2_ow & (idex_ifrdat2_o_17))))

	.dataa(always12),
	.datab(idex_ifrdat2_o_17),
	.datac(fuifrdat2_ow),
	.datad(fuifrtReplace_17),
	.cin(gnd),
	.combout(\rdat2_o~17_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~17 .lut_mask = 16'hA808;
defparam \rdat2_o~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N28
cycloneive_lcell_comb \rdat2_o~18 (
// Equation(s):
// \rdat2_o~18_combout  = (always12 & ((fuifrdat2_ow & ((fuifrtReplace_18))) # (!fuifrdat2_ow & (idex_ifrdat2_o_18))))

	.dataa(idex_ifrdat2_o_18),
	.datab(fuifrtReplace_18),
	.datac(fuifrdat2_ow),
	.datad(always12),
	.cin(gnd),
	.combout(\rdat2_o~18_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~18 .lut_mask = 16'hCA00;
defparam \rdat2_o~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N14
cycloneive_lcell_comb \rdat2_o~19 (
// Equation(s):
// \rdat2_o~19_combout  = (always12 & ((fuifrdat2_ow & ((fuifrtReplace_19))) # (!fuifrdat2_ow & (idex_ifrdat2_o_19))))

	.dataa(fuifrdat2_ow),
	.datab(always12),
	.datac(idex_ifrdat2_o_19),
	.datad(fuifrtReplace_19),
	.cin(gnd),
	.combout(\rdat2_o~19_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~19 .lut_mask = 16'hC840;
defparam \rdat2_o~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N2
cycloneive_lcell_comb \rdat2_o~20 (
// Equation(s):
// \rdat2_o~20_combout  = (always12 & ((fuifrdat2_ow & (fuifrtReplace_20)) # (!fuifrdat2_ow & ((idex_ifrdat2_o_20)))))

	.dataa(always12),
	.datab(fuifrdat2_ow),
	.datac(fuifrtReplace_20),
	.datad(idex_ifrdat2_o_20),
	.cin(gnd),
	.combout(\rdat2_o~20_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~20 .lut_mask = 16'hA280;
defparam \rdat2_o~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N22
cycloneive_lcell_comb \rdat2_o~21 (
// Equation(s):
// \rdat2_o~21_combout  = (always12 & ((fuifrdat2_ow & ((fuifrtReplace_21))) # (!fuifrdat2_ow & (idex_ifrdat2_o_21))))

	.dataa(always12),
	.datab(idex_ifrdat2_o_21),
	.datac(fuifrdat2_ow),
	.datad(fuifrtReplace_21),
	.cin(gnd),
	.combout(\rdat2_o~21_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~21 .lut_mask = 16'hA808;
defparam \rdat2_o~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N26
cycloneive_lcell_comb \rdat2_o~22 (
// Equation(s):
// \rdat2_o~22_combout  = (always12 & ((fuifrdat2_ow & ((fuifrtReplace_22))) # (!fuifrdat2_ow & (idex_ifrdat2_o_22))))

	.dataa(fuifrdat2_ow),
	.datab(idex_ifrdat2_o_22),
	.datac(fuifrtReplace_22),
	.datad(always12),
	.cin(gnd),
	.combout(\rdat2_o~22_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~22 .lut_mask = 16'hE400;
defparam \rdat2_o~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N20
cycloneive_lcell_comb \rdat2_o~23 (
// Equation(s):
// \rdat2_o~23_combout  = (always12 & ((fuifrdat2_ow & (fuifrtReplace_23)) # (!fuifrdat2_ow & ((idex_ifrdat2_o_23)))))

	.dataa(fuifrtReplace_23),
	.datab(fuifrdat2_ow),
	.datac(idex_ifrdat2_o_23),
	.datad(always12),
	.cin(gnd),
	.combout(\rdat2_o~23_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~23 .lut_mask = 16'hB800;
defparam \rdat2_o~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N0
cycloneive_lcell_comb \rdat2_o~24 (
// Equation(s):
// \rdat2_o~24_combout  = (always12 & ((fuifrdat2_ow & (fuifrtReplace_24)) # (!fuifrdat2_ow & ((idex_ifrdat2_o_24)))))

	.dataa(fuifrdat2_ow),
	.datab(fuifrtReplace_24),
	.datac(always12),
	.datad(idex_ifrdat2_o_24),
	.cin(gnd),
	.combout(\rdat2_o~24_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~24 .lut_mask = 16'hD080;
defparam \rdat2_o~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N18
cycloneive_lcell_comb \rdat2_o~25 (
// Equation(s):
// \rdat2_o~25_combout  = (always12 & ((fuifrdat2_ow & ((fuifrtReplace_25))) # (!fuifrdat2_ow & (idex_ifrdat2_o_25))))

	.dataa(fuifrdat2_ow),
	.datab(idex_ifrdat2_o_25),
	.datac(fuifrtReplace_25),
	.datad(always12),
	.cin(gnd),
	.combout(\rdat2_o~25_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~25 .lut_mask = 16'hE400;
defparam \rdat2_o~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N24
cycloneive_lcell_comb \rdat2_o~26 (
// Equation(s):
// \rdat2_o~26_combout  = (always12 & ((fuifrdat2_ow & (fuifrtReplace_26)) # (!fuifrdat2_ow & ((idex_ifrdat2_o_26)))))

	.dataa(fuifrdat2_ow),
	.datab(fuifrtReplace_26),
	.datac(idex_ifrdat2_o_26),
	.datad(always12),
	.cin(gnd),
	.combout(\rdat2_o~26_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~26 .lut_mask = 16'hD800;
defparam \rdat2_o~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N22
cycloneive_lcell_comb \rdat2_o~27 (
// Equation(s):
// \rdat2_o~27_combout  = (always12 & ((fuifrdat2_ow & (fuifrtReplace_27)) # (!fuifrdat2_ow & ((idex_ifrdat2_o_27)))))

	.dataa(fuifrdat2_ow),
	.datab(fuifrtReplace_27),
	.datac(always12),
	.datad(idex_ifrdat2_o_27),
	.cin(gnd),
	.combout(\rdat2_o~27_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~27 .lut_mask = 16'hD080;
defparam \rdat2_o~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N14
cycloneive_lcell_comb \rdat2_o~28 (
// Equation(s):
// \rdat2_o~28_combout  = (always12 & ((fuifrdat2_ow & ((fuifrtReplace_28))) # (!fuifrdat2_ow & (idex_ifrdat2_o_28))))

	.dataa(fuifrdat2_ow),
	.datab(idex_ifrdat2_o_28),
	.datac(fuifrtReplace_28),
	.datad(always12),
	.cin(gnd),
	.combout(\rdat2_o~28_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~28 .lut_mask = 16'hE400;
defparam \rdat2_o~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N30
cycloneive_lcell_comb \rdat2_o~29 (
// Equation(s):
// \rdat2_o~29_combout  = (always12 & ((fuifrdat2_ow & ((fuifrtReplace_29))) # (!fuifrdat2_ow & (idex_ifrdat2_o_29))))

	.dataa(always12),
	.datab(idex_ifrdat2_o_29),
	.datac(fuifrtReplace_29),
	.datad(fuifrdat2_ow),
	.cin(gnd),
	.combout(\rdat2_o~29_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~29 .lut_mask = 16'hA088;
defparam \rdat2_o~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N16
cycloneive_lcell_comb \rdat2_o~30 (
// Equation(s):
// \rdat2_o~30_combout  = (always12 & ((fuifrdat2_ow & (fuifrtReplace_30)) # (!fuifrdat2_ow & ((idex_ifrdat2_o_30)))))

	.dataa(fuifrtReplace_30),
	.datab(always12),
	.datac(idex_ifrdat2_o_30),
	.datad(fuifrdat2_ow),
	.cin(gnd),
	.combout(\rdat2_o~30_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~30 .lut_mask = 16'h88C0;
defparam \rdat2_o~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N26
cycloneive_lcell_comb \rdat2_o~31 (
// Equation(s):
// \rdat2_o~31_combout  = (always12 & ((fuifrdat2_ow & (fuifrtReplace_31)) # (!fuifrdat2_ow & ((idex_ifrdat2_o_31)))))

	.dataa(fuifrdat2_ow),
	.datab(fuifrtReplace_31),
	.datac(idex_ifrdat2_o_31),
	.datad(always12),
	.cin(gnd),
	.combout(\rdat2_o~31_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~31 .lut_mask = 16'hD800;
defparam \rdat2_o~31 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module forward_unit (
	idex_ifrt_o_0,
	idex_ifrt_o_1,
	rwMEM,
	rwMEM1,
	idex_ifrt_o_2,
	idex_ifrt_o_3,
	rwMEM2,
	rwMEM3,
	exmem_ifregWEN_o,
	idex_ifrt_o_4,
	rwMEM4,
	always0,
	rwWB,
	rwWB1,
	rwWB2,
	rwWB3,
	memwb_ifregWEN_o,
	rwWB4,
	always01,
	wdat,
	mem_data,
	fuifrtReplace_1,
	idex_ifrs_o_1,
	idex_ifrs_o_0,
	idex_ifrs_o_3,
	idex_ifrs_o_2,
	idex_ifrs_o_4,
	always02,
	always03,
	mem_data1,
	wdat1,
	fuifrtReplace_0,
	wdat2,
	mem_data2,
	wdat3,
	mem_data3,
	wdat4,
	mem_data4,
	fuifrtReplace_2,
	wdat5,
	mem_data5,
	wdat6,
	mem_data6,
	wdat7,
	mem_data7,
	wdat8,
	mem_data8,
	fuifrtReplace_3,
	wdat9,
	mem_data9,
	wdat10,
	mem_data10,
	wdat11,
	mem_data11,
	wdat12,
	mem_data12,
	wdat13,
	mem_data13,
	wdat14,
	mem_data14,
	wdat15,
	mem_data15,
	wdat16,
	mem_data16,
	fuifrtReplace_4,
	wdat17,
	mem_data17,
	wdat18,
	mem_data18,
	wdat19,
	mem_data19,
	wdat20,
	mem_data20,
	wdat21,
	mem_data21,
	wdat22,
	mem_data22,
	wdat23,
	mem_data23,
	wdat24,
	mem_data24,
	wdat25,
	mem_data25,
	wdat26,
	mem_data26,
	wdat27,
	mem_data27,
	wdat28,
	mem_data28,
	wdat29,
	mem_data29,
	wdat30,
	mem_data30,
	wdat31,
	mem_data31,
	fuifrtReplace_31,
	fuifrtReplace_16,
	fuifrtReplace_17,
	fuifrtReplace_18,
	fuifrtReplace_19,
	fuifrtReplace_20,
	fuifrtReplace_21,
	fuifrtReplace_22,
	fuifrtReplace_23,
	fuifrtReplace_24,
	fuifrtReplace_25,
	fuifrtReplace_26,
	fuifrtReplace_5,
	fuifrtReplace_6,
	fuifrtReplace_7,
	fuifrtReplace_8,
	fuifrtReplace_27,
	fuifrtReplace_28,
	fuifrtReplace_29,
	fuifrtReplace_30,
	fuifrtReplace_9,
	fuifrtReplace_14,
	fuifrtReplace_15,
	fuifrtReplace_10,
	fuifrtReplace_11,
	fuifrtReplace_12,
	fuifrtReplace_13,
	fuifrdat2_ow,
	devpor,
	devclrn,
	devoe);
input 	idex_ifrt_o_0;
input 	idex_ifrt_o_1;
input 	rwMEM;
input 	rwMEM1;
input 	idex_ifrt_o_2;
input 	idex_ifrt_o_3;
input 	rwMEM2;
input 	rwMEM3;
input 	exmem_ifregWEN_o;
input 	idex_ifrt_o_4;
input 	rwMEM4;
output 	always0;
input 	rwWB;
input 	rwWB1;
input 	rwWB2;
input 	rwWB3;
input 	memwb_ifregWEN_o;
input 	rwWB4;
output 	always01;
input 	wdat;
input 	mem_data;
output 	fuifrtReplace_1;
input 	idex_ifrs_o_1;
input 	idex_ifrs_o_0;
input 	idex_ifrs_o_3;
input 	idex_ifrs_o_2;
input 	idex_ifrs_o_4;
output 	always02;
output 	always03;
input 	mem_data1;
input 	wdat1;
output 	fuifrtReplace_0;
input 	wdat2;
input 	mem_data2;
input 	wdat3;
input 	mem_data3;
input 	wdat4;
input 	mem_data4;
output 	fuifrtReplace_2;
input 	wdat5;
input 	mem_data5;
input 	wdat6;
input 	mem_data6;
input 	wdat7;
input 	mem_data7;
input 	wdat8;
input 	mem_data8;
output 	fuifrtReplace_3;
input 	wdat9;
input 	mem_data9;
input 	wdat10;
input 	mem_data10;
input 	wdat11;
input 	mem_data11;
input 	wdat12;
input 	mem_data12;
input 	wdat13;
input 	mem_data13;
input 	wdat14;
input 	mem_data14;
input 	wdat15;
input 	mem_data15;
input 	wdat16;
input 	mem_data16;
output 	fuifrtReplace_4;
input 	wdat17;
input 	mem_data17;
input 	wdat18;
input 	mem_data18;
input 	wdat19;
input 	mem_data19;
input 	wdat20;
input 	mem_data20;
input 	wdat21;
input 	mem_data21;
input 	wdat22;
input 	mem_data22;
input 	wdat23;
input 	mem_data23;
input 	wdat24;
input 	mem_data24;
input 	wdat25;
input 	mem_data25;
input 	wdat26;
input 	mem_data26;
input 	wdat27;
input 	mem_data27;
input 	wdat28;
input 	mem_data28;
input 	wdat29;
input 	mem_data29;
input 	wdat30;
input 	mem_data30;
input 	wdat31;
input 	mem_data31;
output 	fuifrtReplace_31;
output 	fuifrtReplace_16;
output 	fuifrtReplace_17;
output 	fuifrtReplace_18;
output 	fuifrtReplace_19;
output 	fuifrtReplace_20;
output 	fuifrtReplace_21;
output 	fuifrtReplace_22;
output 	fuifrtReplace_23;
output 	fuifrtReplace_24;
output 	fuifrtReplace_25;
output 	fuifrtReplace_26;
output 	fuifrtReplace_5;
output 	fuifrtReplace_6;
output 	fuifrtReplace_7;
output 	fuifrtReplace_8;
output 	fuifrtReplace_27;
output 	fuifrtReplace_28;
output 	fuifrtReplace_29;
output 	fuifrtReplace_30;
output 	fuifrtReplace_9;
output 	fuifrtReplace_14;
output 	fuifrtReplace_15;
output 	fuifrtReplace_10;
output 	fuifrtReplace_11;
output 	fuifrtReplace_12;
output 	fuifrtReplace_13;
output 	fuifrdat2_ow;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \always0~0_combout ;
wire \always0~2_combout ;
wire \always0~1_combout ;
wire \always0~6_combout ;
wire \always0~5_combout ;
wire \always0~4_combout ;
wire \fuif.rtReplace[4]~36_combout ;
wire \always0~8_combout ;
wire \always0~9_combout ;
wire \always0~10_combout ;
wire \always0~14_combout ;
wire \always0~12_combout ;
wire \always0~13_combout ;


// Location: LCCOMB_X56_Y31_N8
cycloneive_lcell_comb \always0~3 (
// Equation(s):
// always0 = (\always0~0_combout  & (\always0~2_combout  & \always0~1_combout ))

	.dataa(\always0~0_combout ),
	.datab(gnd),
	.datac(\always0~2_combout ),
	.datad(\always0~1_combout ),
	.cin(gnd),
	.combout(always0),
	.cout());
// synopsys translate_off
defparam \always0~3 .lut_mask = 16'hA000;
defparam \always0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N0
cycloneive_lcell_comb \always0~7 (
// Equation(s):
// always01 = (\always0~6_combout  & (\always0~5_combout  & \always0~4_combout ))

	.dataa(\always0~6_combout ),
	.datab(gnd),
	.datac(\always0~5_combout ),
	.datad(\always0~4_combout ),
	.cin(gnd),
	.combout(always01),
	.cout());
// synopsys translate_off
defparam \always0~7 .lut_mask = 16'hA000;
defparam \always0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N16
cycloneive_lcell_comb \fuif.rtReplace[1]~4 (
// Equation(s):
// fuifrtReplace_1 = (\fuif.rtReplace[4]~36_combout  & ((\wdat~1_combout ) # ((always0 & \mem_data~4_combout )))) # (!\fuif.rtReplace[4]~36_combout  & (((always0 & \mem_data~4_combout ))))

	.dataa(\fuif.rtReplace[4]~36_combout ),
	.datab(wdat),
	.datac(always0),
	.datad(mem_data),
	.cin(gnd),
	.combout(fuifrtReplace_1),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[1]~4 .lut_mask = 16'hF888;
defparam \fuif.rtReplace[1]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N30
cycloneive_lcell_comb \always0~11 (
// Equation(s):
// always02 = (\always0~8_combout  & (\always0~9_combout  & \always0~10_combout ))

	.dataa(gnd),
	.datab(\always0~8_combout ),
	.datac(\always0~9_combout ),
	.datad(\always0~10_combout ),
	.cin(gnd),
	.combout(always02),
	.cout());
// synopsys translate_off
defparam \always0~11 .lut_mask = 16'hC000;
defparam \always0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N8
cycloneive_lcell_comb \always0~15 (
// Equation(s):
// always03 = (\always0~14_combout  & (\always0~12_combout  & \always0~13_combout ))

	.dataa(\always0~14_combout ),
	.datab(\always0~12_combout ),
	.datac(gnd),
	.datad(\always0~13_combout ),
	.cin(gnd),
	.combout(always03),
	.cout());
// synopsys translate_off
defparam \always0~15 .lut_mask = 16'h8800;
defparam \always0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N6
cycloneive_lcell_comb \fuif.rtReplace[0]~5 (
// Equation(s):
// fuifrtReplace_0 = (\wdat~3_combout  & ((\fuif.rtReplace[4]~36_combout ) # ((always0 & \mem_data~6_combout )))) # (!\wdat~3_combout  & (always0 & (\mem_data~6_combout )))

	.dataa(wdat1),
	.datab(always0),
	.datac(mem_data1),
	.datad(\fuif.rtReplace[4]~36_combout ),
	.cin(gnd),
	.combout(fuifrtReplace_0),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[0]~5 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[0]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N14
cycloneive_lcell_comb \fuif.rtReplace[2]~6 (
// Equation(s):
// fuifrtReplace_2 = (\wdat~5_combout  & ((\fuif.rtReplace[4]~36_combout ) # ((\mem_data~8_combout  & always0)))) # (!\wdat~5_combout  & (((\mem_data~8_combout  & always0))))

	.dataa(wdat2),
	.datab(\fuif.rtReplace[4]~36_combout ),
	.datac(mem_data2),
	.datad(always0),
	.cin(gnd),
	.combout(fuifrtReplace_2),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[2]~6 .lut_mask = 16'hF888;
defparam \fuif.rtReplace[2]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N28
cycloneive_lcell_comb \fuif.rtReplace[3]~7 (
// Equation(s):
// fuifrtReplace_3 = (always0 & ((\mem_data~12_combout ) # ((\wdat~9_combout  & \fuif.rtReplace[4]~36_combout )))) # (!always0 & (\wdat~9_combout  & (\fuif.rtReplace[4]~36_combout )))

	.dataa(always0),
	.datab(wdat4),
	.datac(\fuif.rtReplace[4]~36_combout ),
	.datad(mem_data4),
	.cin(gnd),
	.combout(fuifrtReplace_3),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[3]~7 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[3]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N20
cycloneive_lcell_comb \fuif.rtReplace[4]~8 (
// Equation(s):
// fuifrtReplace_4 = (always0 & ((\mem_data~10_combout ) # ((\fuif.rtReplace[4]~36_combout  & \wdat~7_combout )))) # (!always0 & (\fuif.rtReplace[4]~36_combout  & (\wdat~7_combout )))

	.dataa(always0),
	.datab(\fuif.rtReplace[4]~36_combout ),
	.datac(wdat3),
	.datad(mem_data3),
	.cin(gnd),
	.combout(fuifrtReplace_4),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[4]~8 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[4]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N10
cycloneive_lcell_comb \fuif.rtReplace[31]~9 (
// Equation(s):
// fuifrtReplace_31 = (always0 & ((\mem_data~40_combout ) # ((\wdat~37_combout  & \fuif.rtReplace[4]~36_combout )))) # (!always0 & (\wdat~37_combout  & ((\fuif.rtReplace[4]~36_combout ))))

	.dataa(always0),
	.datab(wdat17),
	.datac(mem_data17),
	.datad(\fuif.rtReplace[4]~36_combout ),
	.cin(gnd),
	.combout(fuifrtReplace_31),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[31]~9 .lut_mask = 16'hECA0;
defparam \fuif.rtReplace[31]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N0
cycloneive_lcell_comb \fuif.rtReplace[16]~10 (
// Equation(s):
// fuifrtReplace_16 = (always0 & ((\mem_data~24_combout ) # ((\fuif.rtReplace[4]~36_combout  & \wdat~21_combout )))) # (!always0 & (\fuif.rtReplace[4]~36_combout  & (\wdat~21_combout )))

	.dataa(always0),
	.datab(\fuif.rtReplace[4]~36_combout ),
	.datac(wdat9),
	.datad(mem_data9),
	.cin(gnd),
	.combout(fuifrtReplace_16),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[16]~10 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[16]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N0
cycloneive_lcell_comb \fuif.rtReplace[17]~11 (
// Equation(s):
// fuifrtReplace_17 = (always0 & ((\mem_data~68_combout ) # ((\fuif.rtReplace[4]~36_combout  & \wdat~65_combout )))) # (!always0 & (\fuif.rtReplace[4]~36_combout  & (\wdat~65_combout )))

	.dataa(always0),
	.datab(\fuif.rtReplace[4]~36_combout ),
	.datac(wdat31),
	.datad(mem_data31),
	.cin(gnd),
	.combout(fuifrtReplace_17),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[17]~11 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[17]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N12
cycloneive_lcell_comb \fuif.rtReplace[18]~12 (
// Equation(s):
// fuifrtReplace_18 = (always0 & ((\mem_data~64_combout ) # ((\fuif.rtReplace[4]~36_combout  & \wdat~61_combout )))) # (!always0 & (\fuif.rtReplace[4]~36_combout  & (\wdat~61_combout )))

	.dataa(always0),
	.datab(\fuif.rtReplace[4]~36_combout ),
	.datac(wdat29),
	.datad(mem_data29),
	.cin(gnd),
	.combout(fuifrtReplace_18),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[18]~12 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[18]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N0
cycloneive_lcell_comb \fuif.rtReplace[19]~13 (
// Equation(s):
// fuifrtReplace_19 = (\fuif.rtReplace[4]~36_combout  & ((\wdat~63_combout ) # ((always0 & \mem_data~66_combout )))) # (!\fuif.rtReplace[4]~36_combout  & (always0 & ((\mem_data~66_combout ))))

	.dataa(\fuif.rtReplace[4]~36_combout ),
	.datab(always0),
	.datac(wdat30),
	.datad(mem_data30),
	.cin(gnd),
	.combout(fuifrtReplace_19),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[19]~13 .lut_mask = 16'hECA0;
defparam \fuif.rtReplace[19]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N0
cycloneive_lcell_comb \fuif.rtReplace[20]~14 (
// Equation(s):
// fuifrtReplace_20 = (always0 & ((\mem_data~62_combout ) # ((\wdat~59_combout  & \fuif.rtReplace[4]~36_combout )))) # (!always0 & (\wdat~59_combout  & (\fuif.rtReplace[4]~36_combout )))

	.dataa(always0),
	.datab(wdat28),
	.datac(\fuif.rtReplace[4]~36_combout ),
	.datad(mem_data28),
	.cin(gnd),
	.combout(fuifrtReplace_20),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[20]~14 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[20]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N28
cycloneive_lcell_comb \fuif.rtReplace[21]~15 (
// Equation(s):
// fuifrtReplace_21 = (always0 & ((\mem_data~60_combout ) # ((\wdat~57_combout  & \fuif.rtReplace[4]~36_combout )))) # (!always0 & (\wdat~57_combout  & (\fuif.rtReplace[4]~36_combout )))

	.dataa(always0),
	.datab(wdat27),
	.datac(\fuif.rtReplace[4]~36_combout ),
	.datad(mem_data27),
	.cin(gnd),
	.combout(fuifrtReplace_21),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[21]~15 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[21]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N6
cycloneive_lcell_comb \fuif.rtReplace[22]~16 (
// Equation(s):
// fuifrtReplace_22 = (always0 & ((\mem_data~56_combout ) # ((\wdat~53_combout  & \fuif.rtReplace[4]~36_combout )))) # (!always0 & (\wdat~53_combout  & (\fuif.rtReplace[4]~36_combout )))

	.dataa(always0),
	.datab(wdat25),
	.datac(\fuif.rtReplace[4]~36_combout ),
	.datad(mem_data25),
	.cin(gnd),
	.combout(fuifrtReplace_22),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[22]~16 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[22]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N10
cycloneive_lcell_comb \fuif.rtReplace[23]~17 (
// Equation(s):
// fuifrtReplace_23 = (\wdat~55_combout  & ((\fuif.rtReplace[4]~36_combout ) # ((always0 & \mem_data~58_combout )))) # (!\wdat~55_combout  & (((always0 & \mem_data~58_combout ))))

	.dataa(wdat26),
	.datab(\fuif.rtReplace[4]~36_combout ),
	.datac(always0),
	.datad(mem_data26),
	.cin(gnd),
	.combout(fuifrtReplace_23),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[23]~17 .lut_mask = 16'hF888;
defparam \fuif.rtReplace[23]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N20
cycloneive_lcell_comb \fuif.rtReplace[24]~18 (
// Equation(s):
// fuifrtReplace_24 = (\fuif.rtReplace[4]~36_combout  & ((\wdat~51_combout ) # ((always0 & \mem_data~54_combout )))) # (!\fuif.rtReplace[4]~36_combout  & (always0 & (\mem_data~54_combout )))

	.dataa(\fuif.rtReplace[4]~36_combout ),
	.datab(always0),
	.datac(mem_data24),
	.datad(wdat24),
	.cin(gnd),
	.combout(fuifrtReplace_24),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[24]~18 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[24]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N2
cycloneive_lcell_comb \fuif.rtReplace[25]~19 (
// Equation(s):
// fuifrtReplace_25 = (\wdat~49_combout  & ((\fuif.rtReplace[4]~36_combout ) # ((always0 & \mem_data~52_combout )))) # (!\wdat~49_combout  & (((always0 & \mem_data~52_combout ))))

	.dataa(wdat23),
	.datab(\fuif.rtReplace[4]~36_combout ),
	.datac(always0),
	.datad(mem_data23),
	.cin(gnd),
	.combout(fuifrtReplace_25),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[25]~19 .lut_mask = 16'hF888;
defparam \fuif.rtReplace[25]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N6
cycloneive_lcell_comb \fuif.rtReplace[26]~20 (
// Equation(s):
// fuifrtReplace_26 = (\fuif.rtReplace[4]~36_combout  & ((\wdat~45_combout ) # ((always0 & \mem_data~48_combout )))) # (!\fuif.rtReplace[4]~36_combout  & (((always0 & \mem_data~48_combout ))))

	.dataa(\fuif.rtReplace[4]~36_combout ),
	.datab(wdat21),
	.datac(always0),
	.datad(mem_data21),
	.cin(gnd),
	.combout(fuifrtReplace_26),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[26]~20 .lut_mask = 16'hF888;
defparam \fuif.rtReplace[26]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N24
cycloneive_lcell_comb \fuif.rtReplace[5]~21 (
// Equation(s):
// fuifrtReplace_5 = (\fuif.rtReplace[4]~36_combout  & ((\wdat~17_combout ) # ((always0 & \mem_data~20_combout )))) # (!\fuif.rtReplace[4]~36_combout  & (((always0 & \mem_data~20_combout ))))

	.dataa(\fuif.rtReplace[4]~36_combout ),
	.datab(wdat8),
	.datac(always0),
	.datad(mem_data8),
	.cin(gnd),
	.combout(fuifrtReplace_5),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[5]~21 .lut_mask = 16'hF888;
defparam \fuif.rtReplace[5]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N16
cycloneive_lcell_comb \fuif.rtReplace[6]~22 (
// Equation(s):
// fuifrtReplace_6 = (always0 & ((\mem_data~18_combout ) # ((\wdat~15_combout  & \fuif.rtReplace[4]~36_combout )))) # (!always0 & (\wdat~15_combout  & (\fuif.rtReplace[4]~36_combout )))

	.dataa(always0),
	.datab(wdat7),
	.datac(\fuif.rtReplace[4]~36_combout ),
	.datad(mem_data7),
	.cin(gnd),
	.combout(fuifrtReplace_6),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[6]~22 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[6]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N0
cycloneive_lcell_comb \fuif.rtReplace[7]~23 (
// Equation(s):
// fuifrtReplace_7 = (always0 & ((\mem_data~16_combout ) # ((\wdat~13_combout  & \fuif.rtReplace[4]~36_combout )))) # (!always0 & (\wdat~13_combout  & ((\fuif.rtReplace[4]~36_combout ))))

	.dataa(always0),
	.datab(wdat6),
	.datac(mem_data6),
	.datad(\fuif.rtReplace[4]~36_combout ),
	.cin(gnd),
	.combout(fuifrtReplace_7),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[7]~23 .lut_mask = 16'hECA0;
defparam \fuif.rtReplace[7]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N28
cycloneive_lcell_comb \fuif.rtReplace[8]~24 (
// Equation(s):
// fuifrtReplace_8 = (always0 & ((\mem_data~14_combout ) # ((\wdat~11_combout  & \fuif.rtReplace[4]~36_combout )))) # (!always0 & (\wdat~11_combout  & (\fuif.rtReplace[4]~36_combout )))

	.dataa(always0),
	.datab(wdat5),
	.datac(\fuif.rtReplace[4]~36_combout ),
	.datad(mem_data5),
	.cin(gnd),
	.combout(fuifrtReplace_8),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[8]~24 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[8]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N18
cycloneive_lcell_comb \fuif.rtReplace[27]~25 (
// Equation(s):
// fuifrtReplace_27 = (\fuif.rtReplace[4]~36_combout  & ((\wdat~47_combout ) # ((always0 & \mem_data~50_combout )))) # (!\fuif.rtReplace[4]~36_combout  & (((always0 & \mem_data~50_combout ))))

	.dataa(\fuif.rtReplace[4]~36_combout ),
	.datab(wdat22),
	.datac(always0),
	.datad(mem_data22),
	.cin(gnd),
	.combout(fuifrtReplace_27),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[27]~25 .lut_mask = 16'hF888;
defparam \fuif.rtReplace[27]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N16
cycloneive_lcell_comb \fuif.rtReplace[28]~26 (
// Equation(s):
// fuifrtReplace_28 = (\fuif.rtReplace[4]~36_combout  & ((\wdat~43_combout ) # ((always0 & \mem_data~46_combout )))) # (!\fuif.rtReplace[4]~36_combout  & (((always0 & \mem_data~46_combout ))))

	.dataa(\fuif.rtReplace[4]~36_combout ),
	.datab(wdat20),
	.datac(always0),
	.datad(mem_data20),
	.cin(gnd),
	.combout(fuifrtReplace_28),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[28]~26 .lut_mask = 16'hF888;
defparam \fuif.rtReplace[28]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N16
cycloneive_lcell_comb \fuif.rtReplace[29]~27 (
// Equation(s):
// fuifrtReplace_29 = (\fuif.rtReplace[4]~36_combout  & ((\wdat~39_combout ) # ((always0 & \mem_data~42_combout )))) # (!\fuif.rtReplace[4]~36_combout  & (((always0 & \mem_data~42_combout ))))

	.dataa(\fuif.rtReplace[4]~36_combout ),
	.datab(wdat18),
	.datac(always0),
	.datad(mem_data18),
	.cin(gnd),
	.combout(fuifrtReplace_29),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[29]~27 .lut_mask = 16'hF888;
defparam \fuif.rtReplace[29]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N28
cycloneive_lcell_comb \fuif.rtReplace[30]~28 (
// Equation(s):
// fuifrtReplace_30 = (\fuif.rtReplace[4]~36_combout  & ((\wdat~41_combout ) # ((always0 & \mem_data~44_combout )))) # (!\fuif.rtReplace[4]~36_combout  & (always0 & ((\mem_data~44_combout ))))

	.dataa(\fuif.rtReplace[4]~36_combout ),
	.datab(always0),
	.datac(wdat19),
	.datad(mem_data19),
	.cin(gnd),
	.combout(fuifrtReplace_30),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[30]~28 .lut_mask = 16'hECA0;
defparam \fuif.rtReplace[30]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N28
cycloneive_lcell_comb \fuif.rtReplace[9]~29 (
// Equation(s):
// fuifrtReplace_9 = (always0 & ((\mem_data~38_combout ) # ((\fuif.rtReplace[4]~36_combout  & \wdat~35_combout )))) # (!always0 & (\fuif.rtReplace[4]~36_combout  & (\wdat~35_combout )))

	.dataa(always0),
	.datab(\fuif.rtReplace[4]~36_combout ),
	.datac(wdat16),
	.datad(mem_data16),
	.cin(gnd),
	.combout(fuifrtReplace_9),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[9]~29 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[9]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N0
cycloneive_lcell_comb \fuif.rtReplace[14]~30 (
// Equation(s):
// fuifrtReplace_14 = (always0 & ((\mem_data~28_combout ) # ((\wdat~25_combout  & \fuif.rtReplace[4]~36_combout )))) # (!always0 & (\wdat~25_combout  & (\fuif.rtReplace[4]~36_combout )))

	.dataa(always0),
	.datab(wdat11),
	.datac(\fuif.rtReplace[4]~36_combout ),
	.datad(mem_data11),
	.cin(gnd),
	.combout(fuifrtReplace_14),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[14]~30 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[14]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N18
cycloneive_lcell_comb \fuif.rtReplace[15]~31 (
// Equation(s):
// fuifrtReplace_15 = (always0 & ((\mem_data~26_combout ) # ((\fuif.rtReplace[4]~36_combout  & \wdat~23_combout )))) # (!always0 & (\fuif.rtReplace[4]~36_combout  & (\wdat~23_combout )))

	.dataa(always0),
	.datab(\fuif.rtReplace[4]~36_combout ),
	.datac(wdat10),
	.datad(mem_data10),
	.cin(gnd),
	.combout(fuifrtReplace_15),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[15]~31 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[15]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N28
cycloneive_lcell_comb \fuif.rtReplace[10]~32 (
// Equation(s):
// fuifrtReplace_10 = (always0 & ((\mem_data~36_combout ) # ((\wdat~33_combout  & \fuif.rtReplace[4]~36_combout )))) # (!always0 & (\wdat~33_combout  & (\fuif.rtReplace[4]~36_combout )))

	.dataa(always0),
	.datab(wdat15),
	.datac(\fuif.rtReplace[4]~36_combout ),
	.datad(mem_data15),
	.cin(gnd),
	.combout(fuifrtReplace_10),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[10]~32 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[10]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N12
cycloneive_lcell_comb \fuif.rtReplace[11]~33 (
// Equation(s):
// fuifrtReplace_11 = (\fuif.rtReplace[4]~36_combout  & ((\wdat~31_combout ) # ((always0 & \mem_data~34_combout )))) # (!\fuif.rtReplace[4]~36_combout  & (((always0 & \mem_data~34_combout ))))

	.dataa(\fuif.rtReplace[4]~36_combout ),
	.datab(wdat14),
	.datac(always0),
	.datad(mem_data14),
	.cin(gnd),
	.combout(fuifrtReplace_11),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[11]~33 .lut_mask = 16'hF888;
defparam \fuif.rtReplace[11]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N22
cycloneive_lcell_comb \fuif.rtReplace[12]~34 (
// Equation(s):
// fuifrtReplace_12 = (\fuif.rtReplace[4]~36_combout  & ((\wdat~29_combout ) # ((always0 & \mem_data~32_combout )))) # (!\fuif.rtReplace[4]~36_combout  & (always0 & ((\mem_data~32_combout ))))

	.dataa(\fuif.rtReplace[4]~36_combout ),
	.datab(always0),
	.datac(wdat13),
	.datad(mem_data13),
	.cin(gnd),
	.combout(fuifrtReplace_12),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[12]~34 .lut_mask = 16'hECA0;
defparam \fuif.rtReplace[12]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N10
cycloneive_lcell_comb \fuif.rtReplace[13]~35 (
// Equation(s):
// fuifrtReplace_13 = (always0 & ((\mem_data~30_combout ) # ((\wdat~27_combout  & \fuif.rtReplace[4]~36_combout )))) # (!always0 & (\wdat~27_combout  & (\fuif.rtReplace[4]~36_combout )))

	.dataa(always0),
	.datab(wdat12),
	.datac(\fuif.rtReplace[4]~36_combout ),
	.datad(mem_data12),
	.cin(gnd),
	.combout(fuifrtReplace_13),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[13]~35 .lut_mask = 16'hEAC0;
defparam \fuif.rtReplace[13]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N12
cycloneive_lcell_comb \fuif.rdat2_ow~0 (
// Equation(s):
// fuifrdat2_ow = (always0) # ((\always0~6_combout  & (\always0~5_combout  & \always0~4_combout )))

	.dataa(\always0~6_combout ),
	.datab(always0),
	.datac(\always0~5_combout ),
	.datad(\always0~4_combout ),
	.cin(gnd),
	.combout(fuifrdat2_ow),
	.cout());
// synopsys translate_off
defparam \fuif.rdat2_ow~0 .lut_mask = 16'hECCC;
defparam \fuif.rdat2_ow~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N26
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// \always0~0_combout  = (idex_ifrt_o_1 & (\rwMEM~0_combout  & (\rwMEM~1_combout  $ (!idex_ifrt_o_0)))) # (!idex_ifrt_o_1 & (!\rwMEM~0_combout  & (\rwMEM~1_combout  $ (!idex_ifrt_o_0))))

	.dataa(idex_ifrt_o_1),
	.datab(rwMEM1),
	.datac(idex_ifrt_o_0),
	.datad(rwMEM),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'h8241;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N22
cycloneive_lcell_comb \always0~2 (
// Equation(s):
// \always0~2_combout  = (exmem_ifregWEN_o & (\rwMEM~4_combout  $ (!idex_ifrt_o_4)))

	.dataa(exmem_ifregWEN_o),
	.datab(rwMEM4),
	.datac(idex_ifrt_o_4),
	.datad(gnd),
	.cin(gnd),
	.combout(\always0~2_combout ),
	.cout());
// synopsys translate_off
defparam \always0~2 .lut_mask = 16'h8282;
defparam \always0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N24
cycloneive_lcell_comb \always0~1 (
// Equation(s):
// \always0~1_combout  = (\rwMEM~2_combout  & (idex_ifrt_o_3 & (idex_ifrt_o_2 $ (!\rwMEM~3_combout )))) # (!\rwMEM~2_combout  & (!idex_ifrt_o_3 & (idex_ifrt_o_2 $ (!\rwMEM~3_combout ))))

	.dataa(rwMEM2),
	.datab(idex_ifrt_o_3),
	.datac(idex_ifrt_o_2),
	.datad(rwMEM3),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
// synopsys translate_off
defparam \always0~1 .lut_mask = 16'h9009;
defparam \always0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N6
cycloneive_lcell_comb \always0~6 (
// Equation(s):
// \always0~6_combout  = (memwb_ifregWEN_o & (idex_ifrt_o_4 $ (!\rwWB~4_combout )))

	.dataa(gnd),
	.datab(idex_ifrt_o_4),
	.datac(memwb_ifregWEN_o),
	.datad(rwWB4),
	.cin(gnd),
	.combout(\always0~6_combout ),
	.cout());
// synopsys translate_off
defparam \always0~6 .lut_mask = 16'hC030;
defparam \always0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N30
cycloneive_lcell_comb \always0~5 (
// Equation(s):
// \always0~5_combout  = (idex_ifrt_o_2 & (\rwWB~3_combout  & (\rwWB~2_combout  $ (!idex_ifrt_o_3)))) # (!idex_ifrt_o_2 & (!\rwWB~3_combout  & (\rwWB~2_combout  $ (!idex_ifrt_o_3))))

	.dataa(idex_ifrt_o_2),
	.datab(rwWB2),
	.datac(idex_ifrt_o_3),
	.datad(rwWB3),
	.cin(gnd),
	.combout(\always0~5_combout ),
	.cout());
// synopsys translate_off
defparam \always0~5 .lut_mask = 16'h8241;
defparam \always0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N28
cycloneive_lcell_comb \always0~4 (
// Equation(s):
// \always0~4_combout  = (\rwWB~0_combout  & (idex_ifrt_o_1 & (idex_ifrt_o_0 $ (!\rwWB~1_combout )))) # (!\rwWB~0_combout  & (!idex_ifrt_o_1 & (idex_ifrt_o_0 $ (!\rwWB~1_combout ))))

	.dataa(rwWB),
	.datab(idex_ifrt_o_0),
	.datac(idex_ifrt_o_1),
	.datad(rwWB1),
	.cin(gnd),
	.combout(\always0~4_combout ),
	.cout());
// synopsys translate_off
defparam \always0~4 .lut_mask = 16'h8421;
defparam \always0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N2
cycloneive_lcell_comb \fuif.rtReplace[4]~36 (
// Equation(s):
// \fuif.rtReplace[4]~36_combout  = (\always0~6_combout  & (!always0 & (\always0~5_combout  & \always0~4_combout )))

	.dataa(\always0~6_combout ),
	.datab(always0),
	.datac(\always0~5_combout ),
	.datad(\always0~4_combout ),
	.cin(gnd),
	.combout(\fuif.rtReplace[4]~36_combout ),
	.cout());
// synopsys translate_off
defparam \fuif.rtReplace[4]~36 .lut_mask = 16'h2000;
defparam \fuif.rtReplace[4]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N18
cycloneive_lcell_comb \always0~8 (
// Equation(s):
// \always0~8_combout  = (idex_ifrs_o_0 & (\rwWB~1_combout  & (\rwWB~0_combout  $ (!idex_ifrs_o_1)))) # (!idex_ifrs_o_0 & (!\rwWB~1_combout  & (\rwWB~0_combout  $ (!idex_ifrs_o_1))))

	.dataa(idex_ifrs_o_0),
	.datab(rwWB1),
	.datac(rwWB),
	.datad(idex_ifrs_o_1),
	.cin(gnd),
	.combout(\always0~8_combout ),
	.cout());
// synopsys translate_off
defparam \always0~8 .lut_mask = 16'h9009;
defparam \always0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N22
cycloneive_lcell_comb \always0~9 (
// Equation(s):
// \always0~9_combout  = (\rwWB~2_combout  & (idex_ifrs_o_3 & (\rwWB~3_combout  $ (!idex_ifrs_o_2)))) # (!\rwWB~2_combout  & (!idex_ifrs_o_3 & (\rwWB~3_combout  $ (!idex_ifrs_o_2))))

	.dataa(rwWB2),
	.datab(rwWB3),
	.datac(idex_ifrs_o_3),
	.datad(idex_ifrs_o_2),
	.cin(gnd),
	.combout(\always0~9_combout ),
	.cout());
// synopsys translate_off
defparam \always0~9 .lut_mask = 16'h8421;
defparam \always0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N16
cycloneive_lcell_comb \always0~10 (
// Equation(s):
// \always0~10_combout  = (memwb_ifregWEN_o & (\rwWB~4_combout  $ (!idex_ifrs_o_4)))

	.dataa(rwWB4),
	.datab(gnd),
	.datac(memwb_ifregWEN_o),
	.datad(idex_ifrs_o_4),
	.cin(gnd),
	.combout(\always0~10_combout ),
	.cout());
// synopsys translate_off
defparam \always0~10 .lut_mask = 16'hA050;
defparam \always0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N12
cycloneive_lcell_comb \always0~14 (
// Equation(s):
// \always0~14_combout  = (exmem_ifregWEN_o & (idex_ifrs_o_4 $ (!\rwMEM~4_combout )))

	.dataa(idex_ifrs_o_4),
	.datab(rwMEM4),
	.datac(exmem_ifregWEN_o),
	.datad(gnd),
	.cin(gnd),
	.combout(\always0~14_combout ),
	.cout());
// synopsys translate_off
defparam \always0~14 .lut_mask = 16'h9090;
defparam \always0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N20
cycloneive_lcell_comb \always0~12 (
// Equation(s):
// \always0~12_combout  = (\rwMEM~1_combout  & (idex_ifrs_o_0 & (idex_ifrs_o_1 $ (!\rwMEM~0_combout )))) # (!\rwMEM~1_combout  & (!idex_ifrs_o_0 & (idex_ifrs_o_1 $ (!\rwMEM~0_combout ))))

	.dataa(rwMEM1),
	.datab(idex_ifrs_o_0),
	.datac(idex_ifrs_o_1),
	.datad(rwMEM),
	.cin(gnd),
	.combout(\always0~12_combout ),
	.cout());
// synopsys translate_off
defparam \always0~12 .lut_mask = 16'h9009;
defparam \always0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N18
cycloneive_lcell_comb \always0~13 (
// Equation(s):
// \always0~13_combout  = (\rwMEM~3_combout  & (idex_ifrs_o_2 & (idex_ifrs_o_3 $ (!\rwMEM~2_combout )))) # (!\rwMEM~3_combout  & (!idex_ifrs_o_2 & (idex_ifrs_o_3 $ (!\rwMEM~2_combout ))))

	.dataa(rwMEM3),
	.datab(idex_ifrs_o_3),
	.datac(rwMEM2),
	.datad(idex_ifrs_o_2),
	.cin(gnd),
	.combout(\always0~13_combout ),
	.cout());
// synopsys translate_off
defparam \always0~13 .lut_mask = 16'h8241;
defparam \always0~13 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module hazard_unit (
	exmem_ifdWEN_o,
	exmem_ifdREN_o,
	rwMEM,
	rwMEM1,
	rwMEM2,
	rwMEM3,
	exmem_ifregWEN_o,
	rwMEM4,
	myifout_1,
	idex_ifjumpSel_o_1,
	idex_ifjumpSel_o_0,
	idex_ifinstr_o_31,
	idex_ifinstr_o_30,
	idex_ifinstr_o_27,
	idex_ifinstr_o_26,
	idex_ifinstr_o_28,
	ifid_ifinstr_o_17,
	ifid_ifinstr_o_16,
	ifid_ifinstr_o_19,
	ifid_ifinstr_o_18,
	ifid_ifinstr_o_20,
	ifid_ifinstr_o_22,
	ifid_ifinstr_o_21,
	ifid_ifinstr_o_24,
	ifid_ifinstr_o_23,
	ifid_ifinstr_o_25,
	huiffreeze,
	idex_ifbne_o,
	Equal10,
	Equal101,
	flush,
	idex_ifPCSel_o,
	huifflush,
	devpor,
	devclrn,
	devoe);
input 	exmem_ifdWEN_o;
input 	exmem_ifdREN_o;
input 	rwMEM;
input 	rwMEM1;
input 	rwMEM2;
input 	rwMEM3;
input 	exmem_ifregWEN_o;
input 	rwMEM4;
input 	myifout_1;
input 	idex_ifjumpSel_o_1;
input 	idex_ifjumpSel_o_0;
input 	idex_ifinstr_o_31;
input 	idex_ifinstr_o_30;
input 	idex_ifinstr_o_27;
input 	idex_ifinstr_o_26;
input 	idex_ifinstr_o_28;
input 	ifid_ifinstr_o_17;
input 	ifid_ifinstr_o_16;
input 	ifid_ifinstr_o_19;
input 	ifid_ifinstr_o_18;
input 	ifid_ifinstr_o_20;
input 	ifid_ifinstr_o_22;
input 	ifid_ifinstr_o_21;
input 	ifid_ifinstr_o_24;
input 	ifid_ifinstr_o_23;
input 	ifid_ifinstr_o_25;
output 	huiffreeze;
input 	idex_ifbne_o;
input 	Equal10;
input 	Equal101;
output 	flush;
input 	idex_ifPCSel_o;
output 	huifflush;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Equal2~1_combout ;
wire \Equal2~0_combout ;
wire \Equal2~2_combout ;
wire \Equal3~1_combout ;
wire \Equal3~0_combout ;
wire \Equal3~2_combout ;
wire \huif.freeze~1_combout ;
wire \huif.freeze~0_combout ;


// Location: LCCOMB_X57_Y27_N18
cycloneive_lcell_comb \huif.freeze~2 (
// Equation(s):
// huiffreeze = (\huif.freeze~1_combout  & (\huif.freeze~0_combout  & ((\Equal2~2_combout ) # (\Equal3~2_combout ))))

	.dataa(\Equal2~2_combout ),
	.datab(\Equal3~2_combout ),
	.datac(\huif.freeze~1_combout ),
	.datad(\huif.freeze~0_combout ),
	.cin(gnd),
	.combout(huiffreeze),
	.cout());
// synopsys translate_off
defparam \huif.freeze~2 .lut_mask = 16'hE000;
defparam \huif.freeze~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N10
cycloneive_lcell_comb \flush~0 (
// Equation(s):
// flush = idex_ifbne_o $ (((!myifout_1 & (Equal101 & Equal10))))

	.dataa(myifout_1),
	.datab(idex_ifbne_o),
	.datac(Equal101),
	.datad(Equal10),
	.cin(gnd),
	.combout(flush),
	.cout());
// synopsys translate_off
defparam \flush~0 .lut_mask = 16'h9CCC;
defparam \flush~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N0
cycloneive_lcell_comb \huif.flush~0 (
// Equation(s):
// huifflush = (idex_ifjumpSel_o_0 & (((idex_ifPCSel_o & flush)) # (!idex_ifjumpSel_o_1))) # (!idex_ifjumpSel_o_0 & (((idex_ifjumpSel_o_1))))

	.dataa(idex_ifjumpSel_o_0),
	.datab(idex_ifPCSel_o),
	.datac(idex_ifjumpSel_o_1),
	.datad(flush),
	.cin(gnd),
	.combout(huifflush),
	.cout());
// synopsys translate_off
defparam \huif.flush~0 .lut_mask = 16'hDA5A;
defparam \huif.flush~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N8
cycloneive_lcell_comb \Equal2~1 (
// Equation(s):
// \Equal2~1_combout  = (\rwMEM~3_combout  & (ifid_ifinstr_o_18 & (\rwMEM~2_combout  $ (!ifid_ifinstr_o_19)))) # (!\rwMEM~3_combout  & (!ifid_ifinstr_o_18 & (\rwMEM~2_combout  $ (!ifid_ifinstr_o_19))))

	.dataa(rwMEM3),
	.datab(rwMEM2),
	.datac(ifid_ifinstr_o_18),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~1 .lut_mask = 16'h8421;
defparam \Equal2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N0
cycloneive_lcell_comb \Equal2~0 (
// Equation(s):
// \Equal2~0_combout  = (\rwMEM~1_combout  & (ifid_ifinstr_o_16 & (\rwMEM~0_combout  $ (!ifid_ifinstr_o_17)))) # (!\rwMEM~1_combout  & (!ifid_ifinstr_o_16 & (\rwMEM~0_combout  $ (!ifid_ifinstr_o_17))))

	.dataa(rwMEM1),
	.datab(rwMEM),
	.datac(ifid_ifinstr_o_17),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~0 .lut_mask = 16'h8241;
defparam \Equal2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N26
cycloneive_lcell_comb \Equal2~2 (
// Equation(s):
// \Equal2~2_combout  = (\Equal2~1_combout  & (\Equal2~0_combout  & (\rwMEM~4_combout  $ (!ifid_ifinstr_o_20))))

	.dataa(rwMEM4),
	.datab(ifid_ifinstr_o_20),
	.datac(\Equal2~1_combout ),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(\Equal2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~2 .lut_mask = 16'h9000;
defparam \Equal2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N2
cycloneive_lcell_comb \Equal3~1 (
// Equation(s):
// \Equal3~1_combout  = (\rwMEM~3_combout  & (ifid_ifinstr_o_23 & (\rwMEM~2_combout  $ (!ifid_ifinstr_o_24)))) # (!\rwMEM~3_combout  & (!ifid_ifinstr_o_23 & (\rwMEM~2_combout  $ (!ifid_ifinstr_o_24))))

	.dataa(rwMEM3),
	.datab(rwMEM2),
	.datac(ifid_ifinstr_o_23),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Equal3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~1 .lut_mask = 16'h8421;
defparam \Equal3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N16
cycloneive_lcell_comb \Equal3~0 (
// Equation(s):
// \Equal3~0_combout  = (\rwMEM~1_combout  & (ifid_ifinstr_o_21 & (\rwMEM~0_combout  $ (!ifid_ifinstr_o_22)))) # (!\rwMEM~1_combout  & (!ifid_ifinstr_o_21 & (\rwMEM~0_combout  $ (!ifid_ifinstr_o_22))))

	.dataa(rwMEM1),
	.datab(rwMEM),
	.datac(ifid_ifinstr_o_21),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Equal3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~0 .lut_mask = 16'h8421;
defparam \Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N28
cycloneive_lcell_comb \Equal3~2 (
// Equation(s):
// \Equal3~2_combout  = (\Equal3~1_combout  & (\Equal3~0_combout  & (\rwMEM~4_combout  $ (!ifid_ifinstr_o_25))))

	.dataa(rwMEM4),
	.datab(\Equal3~1_combout ),
	.datac(ifid_ifinstr_o_25),
	.datad(\Equal3~0_combout ),
	.cin(gnd),
	.combout(\Equal3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~2 .lut_mask = 16'h8400;
defparam \Equal3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N14
cycloneive_lcell_comb \huif.freeze~1 (
// Equation(s):
// \huif.freeze~1_combout  = (!idex_ifinstr_o_28 & (exmem_ifregWEN_o & (idex_ifinstr_o_27 & idex_ifinstr_o_26)))

	.dataa(idex_ifinstr_o_28),
	.datab(exmem_ifregWEN_o),
	.datac(idex_ifinstr_o_27),
	.datad(idex_ifinstr_o_26),
	.cin(gnd),
	.combout(\huif.freeze~1_combout ),
	.cout());
// synopsys translate_off
defparam \huif.freeze~1 .lut_mask = 16'h4000;
defparam \huif.freeze~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N20
cycloneive_lcell_comb \huif.freeze~0 (
// Equation(s):
// \huif.freeze~0_combout  = (!idex_ifinstr_o_30 & (idex_ifinstr_o_31 & (!exmem_ifdWEN_o & !exmem_ifdREN_o)))

	.dataa(idex_ifinstr_o_30),
	.datab(idex_ifinstr_o_31),
	.datac(exmem_ifdWEN_o),
	.datad(exmem_ifdREN_o),
	.cin(gnd),
	.combout(\huif.freeze~0_combout ),
	.cout());
// synopsys translate_off
defparam \huif.freeze~0 .lut_mask = 16'h0004;
defparam \huif.freeze~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module id_ex (
	idex_ifaluop_o_1,
	idex_ifrt_o_0,
	idex_ifrt_o_1,
	idex_ifrt_o_2,
	idex_ifrt_o_3,
	idex_ifrt_o_4,
	idex_ifALUSel_o_1,
	idex_ifALUSel_o_0,
	idex_ifimm_o_1,
	idex_ifshamt_o_1,
	idex_ifrdat2_o_1,
	idex_ifrdat1_o_1,
	idex_ifrs_o_1,
	idex_ifrs_o_0,
	idex_ifrs_o_3,
	idex_ifrs_o_2,
	idex_ifrs_o_4,
	idex_ifimm_o_0,
	idex_ifshamt_o_0,
	idex_ifrdat2_o_0,
	idex_ifrdat1_o_0,
	idex_ifaluop_o_2,
	idex_ifrdat1_o_2,
	idex_ifrdat1_o_4,
	idex_ifrdat1_o_3,
	idex_ifimm_o_2,
	idex_ifshamt_o_2,
	idex_ifrdat2_o_2,
	idex_ifrdat1_o_8,
	idex_ifrdat1_o_7,
	idex_ifrdat1_o_6,
	idex_ifrdat1_o_5,
	idex_ifrdat2_o_3,
	idex_ifimm_o_3,
	idex_ifshamt_o_3,
	idex_ifrdat1_o_16,
	idex_ifrdat1_o_15,
	idex_ifrdat1_o_14,
	idex_ifrdat1_o_13,
	idex_ifrdat1_o_12,
	idex_ifrdat1_o_11,
	idex_ifrdat1_o_10,
	idex_ifrdat1_o_9,
	idex_ifrdat2_o_4,
	idex_ifimm_o_4,
	idex_ifshamt_o_4,
	idex_ifrdat1_o_31,
	idex_ifrdat1_o_29,
	idex_ifrdat1_o_30,
	idex_ifrdat1_o_28,
	idex_ifrdat1_o_26,
	idex_ifrdat1_o_27,
	idex_ifrdat1_o_25,
	idex_ifrdat1_o_24,
	idex_ifrdat1_o_22,
	idex_ifrdat1_o_23,
	idex_ifrdat1_o_21,
	idex_ifrdat1_o_20,
	idex_ifrdat1_o_18,
	idex_ifrdat1_o_19,
	idex_ifrdat1_o_17,
	idex_ifimm_o_15,
	idex_ifrdat2_o_31,
	idex_ifrdat2_o_16,
	idex_ifrdat2_o_17,
	idex_ifrdat2_o_18,
	idex_ifrdat2_o_19,
	idex_ifrdat2_o_20,
	idex_ifrdat2_o_21,
	idex_ifrdat2_o_22,
	idex_ifrdat2_o_23,
	idex_ifrdat2_o_24,
	idex_ifrdat2_o_25,
	idex_ifrdat2_o_26,
	idex_ifrdat2_o_5,
	idex_ifimm_o_5,
	idex_ifrdat2_o_6,
	idex_ifimm_o_6,
	idex_ifrdat2_o_7,
	idex_ifimm_o_7,
	idex_ifrdat2_o_8,
	idex_ifimm_o_8,
	idex_ifrdat2_o_27,
	idex_ifrdat2_o_28,
	idex_ifrdat2_o_29,
	idex_ifrdat2_o_30,
	idex_ifrdat2_o_9,
	idex_ifimm_o_9,
	idex_ifrdat2_o_14,
	idex_ifimm_o_14,
	idex_ifrdat2_o_15,
	idex_ifrdat2_o_10,
	idex_ifimm_o_10,
	idex_ifrdat2_o_11,
	idex_ifimm_o_11,
	idex_ifrdat2_o_12,
	idex_ifimm_o_12,
	idex_ifrdat2_o_13,
	idex_ifimm_o_13,
	idex_ifaluop_o_0,
	idex_ifaluop_o_3,
	idex_ifdWEN_o,
	idex_ifdREN_o,
	idex_ifnext_pc_o_1,
	idex_ifjumpSel_o_1,
	idex_ifjumpSel_o_0,
	always1,
	idex_ifinstr_o_31,
	idex_ifinstr_o_30,
	idex_ifinstr_o_27,
	idex_ifinstr_o_26,
	idex_ifinstr_o_28,
	ifid_ifinstr_o_17,
	ifid_ifinstr_o_16,
	ifid_ifinstr_o_19,
	ifid_ifinstr_o_18,
	ifid_ifinstr_o_20,
	ifid_ifinstr_o_22,
	ifid_ifinstr_o_21,
	ifid_ifinstr_o_24,
	ifid_ifinstr_o_23,
	ifid_ifinstr_o_25,
	huiffreeze,
	idex_ifbne_o,
	idex_ifPCSel_o,
	huifflush,
	idex_ifnext_pc_o_0,
	idex_ifnext_pc_o_3,
	idex_ifnext_pc_o_2,
	idex_ifimm_26_o_1,
	idex_ifimm_26_o_0,
	idex_ifnext_pc_o_5,
	idex_ifnext_pc_o_4,
	idex_ifimm_26_o_3,
	idex_ifimm_26_o_2,
	idex_ifnext_pc_o_7,
	idex_ifnext_pc_o_6,
	idex_ifimm_26_o_5,
	idex_ifimm_26_o_4,
	idex_ifnext_pc_o_9,
	idex_ifnext_pc_o_8,
	idex_ifimm_26_o_7,
	idex_ifimm_26_o_6,
	idex_ifnext_pc_o_11,
	idex_ifnext_pc_o_10,
	idex_ifimm_26_o_9,
	idex_ifimm_26_o_8,
	idex_ifnext_pc_o_13,
	idex_ifnext_pc_o_12,
	idex_ifimm_26_o_11,
	idex_ifimm_26_o_10,
	idex_ifnext_pc_o_15,
	idex_ifnext_pc_o_14,
	idex_ifimm_26_o_13,
	idex_ifimm_26_o_12,
	idex_ifnext_pc_o_17,
	idex_ifnext_pc_o_16,
	idex_ifimm_26_o_15,
	idex_ifimm_26_o_14,
	idex_ifnext_pc_o_19,
	idex_ifnext_pc_o_18,
	idex_ifimm_26_o_17,
	idex_ifimm_26_o_16,
	idex_ifnext_pc_o_21,
	idex_ifnext_pc_o_20,
	idex_ifimm_26_o_19,
	idex_ifimm_26_o_18,
	idex_ifnext_pc_o_23,
	idex_ifnext_pc_o_22,
	idex_ifimm_26_o_21,
	idex_ifimm_26_o_20,
	idex_ifnext_pc_o_25,
	idex_ifnext_pc_o_24,
	idex_ifimm_26_o_23,
	idex_ifimm_26_o_22,
	idex_ifnext_pc_o_27,
	idex_ifnext_pc_o_26,
	idex_ifimm_26_o_25,
	idex_ifimm_26_o_24,
	idex_ifnext_pc_o_29,
	idex_ifnext_pc_o_28,
	idex_ifnext_pc_o_31,
	idex_ifnext_pc_o_30,
	idex_ifhalt_o,
	ifid_ifinstr_o_26,
	ifid_ifinstr_o_31,
	ifid_ifinstr_o_27,
	ifid_ifinstr_o_28,
	ifid_ifinstr_o_30,
	ifid_ifinstr_o_5,
	ifid_ifinstr_o_4,
	always0,
	ifid_ifinstr_o_29,
	ifid_ifinstr_o_1,
	ifid_ifinstr_o_3,
	ifid_ifinstr_o_2,
	idex_ifRegDest_o_1,
	idex_ifrd_o_1,
	idex_ifRegDest_o_0,
	idex_ifrd_o_0,
	idex_ifrd_o_3,
	idex_ifrd_o_2,
	idex_ifregWEN_o,
	idex_ifrd_o_4,
	cuifregWEN,
	Equal0,
	ifid_ifinstr_o_0,
	Equal3,
	Equal2,
	idex_ifjal_o,
	idex_iflui_o,
	idex_ifmemToReg_o,
	ifid_ifinstr_o_7,
	Mux62,
	Mux621,
	Mux30,
	Mux301,
	ifid_ifinstr_o_6,
	Mux63,
	Mux631,
	Mux31,
	Mux311,
	Equal10,
	Mux29,
	Mux291,
	Mux27,
	Mux271,
	Mux28,
	Mux281,
	ifid_ifinstr_o_8,
	Mux61,
	Mux611,
	Mux23,
	Mux231,
	Mux24,
	Mux241,
	Mux25,
	Mux251,
	Mux26,
	Mux261,
	Mux60,
	Mux601,
	ifid_ifinstr_o_9,
	Mux15,
	Mux151,
	Mux16,
	Mux161,
	Mux17,
	Mux171,
	Mux18,
	Mux181,
	Mux19,
	Mux191,
	Mux20,
	Mux201,
	Mux21,
	Mux211,
	Mux22,
	Mux221,
	Mux59,
	Mux591,
	ifid_ifinstr_o_10,
	Mux0,
	Mux01,
	Mux2,
	Mux210,
	Mux1,
	Mux11,
	Mux3,
	Mux32,
	Mux5,
	Mux51,
	Mux4,
	Mux41,
	Mux6,
	Mux64,
	Mux7,
	Mux71,
	Mux9,
	Mux91,
	Mux8,
	Mux81,
	Mux10,
	Mux101,
	Mux111,
	Mux112,
	Mux13,
	Mux131,
	Mux12,
	Mux121,
	Mux14,
	Mux141,
	ifid_ifinstr_o_15,
	Mux321,
	Mux322,
	Mux47,
	Mux471,
	Mux46,
	Mux461,
	Mux45,
	Mux451,
	Mux44,
	Mux441,
	Mux43,
	Mux431,
	Mux42,
	Mux421,
	Mux411,
	Mux412,
	Mux40,
	Mux401,
	Mux39,
	Mux391,
	Mux38,
	Mux381,
	Mux37,
	Mux371,
	Mux58,
	Mux581,
	Mux57,
	Mux571,
	Mux56,
	Mux561,
	Mux55,
	Mux551,
	Mux36,
	Mux361,
	Mux35,
	Mux351,
	Mux34,
	Mux341,
	Mux33,
	Mux331,
	Mux54,
	Mux541,
	Mux49,
	Mux491,
	ifid_ifinstr_o_14,
	Mux48,
	Mux481,
	Mux53,
	Mux531,
	Mux52,
	Mux521,
	ifid_ifinstr_o_11,
	Mux511,
	Mux512,
	ifid_ifinstr_o_12,
	Mux50,
	Mux501,
	ifid_ifinstr_o_13,
	Equal14,
	Equal21,
	Equal01,
	ifid_ifnext_pc_o_1,
	Equal5,
	ifid_ifnext_pc_o_0,
	ifid_ifnext_pc_o_3,
	ifid_ifnext_pc_o_2,
	ifid_ifnext_pc_o_5,
	ifid_ifnext_pc_o_4,
	ifid_ifnext_pc_o_7,
	ifid_ifnext_pc_o_6,
	ifid_ifnext_pc_o_9,
	ifid_ifnext_pc_o_8,
	ifid_ifnext_pc_o_11,
	ifid_ifnext_pc_o_10,
	ifid_ifnext_pc_o_13,
	ifid_ifnext_pc_o_12,
	ifid_ifnext_pc_o_15,
	ifid_ifnext_pc_o_14,
	ifid_ifnext_pc_o_17,
	ifid_ifnext_pc_o_16,
	ifid_ifnext_pc_o_19,
	ifid_ifnext_pc_o_18,
	ifid_ifnext_pc_o_21,
	ifid_ifnext_pc_o_20,
	ifid_ifnext_pc_o_23,
	ifid_ifnext_pc_o_22,
	ifid_ifnext_pc_o_25,
	ifid_ifnext_pc_o_24,
	ifid_ifnext_pc_o_27,
	ifid_ifnext_pc_o_26,
	ifid_ifnext_pc_o_29,
	ifid_ifnext_pc_o_28,
	ifid_ifnext_pc_o_31,
	ifid_ifnext_pc_o_30,
	cuifregWEN1,
	Equal1,
	CPUCLK,
	nRST,
	devpor,
	devclrn,
	devoe);
output 	idex_ifaluop_o_1;
output 	idex_ifrt_o_0;
output 	idex_ifrt_o_1;
output 	idex_ifrt_o_2;
output 	idex_ifrt_o_3;
output 	idex_ifrt_o_4;
output 	idex_ifALUSel_o_1;
output 	idex_ifALUSel_o_0;
output 	idex_ifimm_o_1;
output 	idex_ifshamt_o_1;
output 	idex_ifrdat2_o_1;
output 	idex_ifrdat1_o_1;
output 	idex_ifrs_o_1;
output 	idex_ifrs_o_0;
output 	idex_ifrs_o_3;
output 	idex_ifrs_o_2;
output 	idex_ifrs_o_4;
output 	idex_ifimm_o_0;
output 	idex_ifshamt_o_0;
output 	idex_ifrdat2_o_0;
output 	idex_ifrdat1_o_0;
output 	idex_ifaluop_o_2;
output 	idex_ifrdat1_o_2;
output 	idex_ifrdat1_o_4;
output 	idex_ifrdat1_o_3;
output 	idex_ifimm_o_2;
output 	idex_ifshamt_o_2;
output 	idex_ifrdat2_o_2;
output 	idex_ifrdat1_o_8;
output 	idex_ifrdat1_o_7;
output 	idex_ifrdat1_o_6;
output 	idex_ifrdat1_o_5;
output 	idex_ifrdat2_o_3;
output 	idex_ifimm_o_3;
output 	idex_ifshamt_o_3;
output 	idex_ifrdat1_o_16;
output 	idex_ifrdat1_o_15;
output 	idex_ifrdat1_o_14;
output 	idex_ifrdat1_o_13;
output 	idex_ifrdat1_o_12;
output 	idex_ifrdat1_o_11;
output 	idex_ifrdat1_o_10;
output 	idex_ifrdat1_o_9;
output 	idex_ifrdat2_o_4;
output 	idex_ifimm_o_4;
output 	idex_ifshamt_o_4;
output 	idex_ifrdat1_o_31;
output 	idex_ifrdat1_o_29;
output 	idex_ifrdat1_o_30;
output 	idex_ifrdat1_o_28;
output 	idex_ifrdat1_o_26;
output 	idex_ifrdat1_o_27;
output 	idex_ifrdat1_o_25;
output 	idex_ifrdat1_o_24;
output 	idex_ifrdat1_o_22;
output 	idex_ifrdat1_o_23;
output 	idex_ifrdat1_o_21;
output 	idex_ifrdat1_o_20;
output 	idex_ifrdat1_o_18;
output 	idex_ifrdat1_o_19;
output 	idex_ifrdat1_o_17;
output 	idex_ifimm_o_15;
output 	idex_ifrdat2_o_31;
output 	idex_ifrdat2_o_16;
output 	idex_ifrdat2_o_17;
output 	idex_ifrdat2_o_18;
output 	idex_ifrdat2_o_19;
output 	idex_ifrdat2_o_20;
output 	idex_ifrdat2_o_21;
output 	idex_ifrdat2_o_22;
output 	idex_ifrdat2_o_23;
output 	idex_ifrdat2_o_24;
output 	idex_ifrdat2_o_25;
output 	idex_ifrdat2_o_26;
output 	idex_ifrdat2_o_5;
output 	idex_ifimm_o_5;
output 	idex_ifrdat2_o_6;
output 	idex_ifimm_o_6;
output 	idex_ifrdat2_o_7;
output 	idex_ifimm_o_7;
output 	idex_ifrdat2_o_8;
output 	idex_ifimm_o_8;
output 	idex_ifrdat2_o_27;
output 	idex_ifrdat2_o_28;
output 	idex_ifrdat2_o_29;
output 	idex_ifrdat2_o_30;
output 	idex_ifrdat2_o_9;
output 	idex_ifimm_o_9;
output 	idex_ifrdat2_o_14;
output 	idex_ifimm_o_14;
output 	idex_ifrdat2_o_15;
output 	idex_ifrdat2_o_10;
output 	idex_ifimm_o_10;
output 	idex_ifrdat2_o_11;
output 	idex_ifimm_o_11;
output 	idex_ifrdat2_o_12;
output 	idex_ifimm_o_12;
output 	idex_ifrdat2_o_13;
output 	idex_ifimm_o_13;
output 	idex_ifaluop_o_0;
output 	idex_ifaluop_o_3;
output 	idex_ifdWEN_o;
output 	idex_ifdREN_o;
output 	idex_ifnext_pc_o_1;
output 	idex_ifjumpSel_o_1;
output 	idex_ifjumpSel_o_0;
input 	always1;
output 	idex_ifinstr_o_31;
output 	idex_ifinstr_o_30;
output 	idex_ifinstr_o_27;
output 	idex_ifinstr_o_26;
output 	idex_ifinstr_o_28;
input 	ifid_ifinstr_o_17;
input 	ifid_ifinstr_o_16;
input 	ifid_ifinstr_o_19;
input 	ifid_ifinstr_o_18;
input 	ifid_ifinstr_o_20;
input 	ifid_ifinstr_o_22;
input 	ifid_ifinstr_o_21;
input 	ifid_ifinstr_o_24;
input 	ifid_ifinstr_o_23;
input 	ifid_ifinstr_o_25;
input 	huiffreeze;
output 	idex_ifbne_o;
output 	idex_ifPCSel_o;
input 	huifflush;
output 	idex_ifnext_pc_o_0;
output 	idex_ifnext_pc_o_3;
output 	idex_ifnext_pc_o_2;
output 	idex_ifimm_26_o_1;
output 	idex_ifimm_26_o_0;
output 	idex_ifnext_pc_o_5;
output 	idex_ifnext_pc_o_4;
output 	idex_ifimm_26_o_3;
output 	idex_ifimm_26_o_2;
output 	idex_ifnext_pc_o_7;
output 	idex_ifnext_pc_o_6;
output 	idex_ifimm_26_o_5;
output 	idex_ifimm_26_o_4;
output 	idex_ifnext_pc_o_9;
output 	idex_ifnext_pc_o_8;
output 	idex_ifimm_26_o_7;
output 	idex_ifimm_26_o_6;
output 	idex_ifnext_pc_o_11;
output 	idex_ifnext_pc_o_10;
output 	idex_ifimm_26_o_9;
output 	idex_ifimm_26_o_8;
output 	idex_ifnext_pc_o_13;
output 	idex_ifnext_pc_o_12;
output 	idex_ifimm_26_o_11;
output 	idex_ifimm_26_o_10;
output 	idex_ifnext_pc_o_15;
output 	idex_ifnext_pc_o_14;
output 	idex_ifimm_26_o_13;
output 	idex_ifimm_26_o_12;
output 	idex_ifnext_pc_o_17;
output 	idex_ifnext_pc_o_16;
output 	idex_ifimm_26_o_15;
output 	idex_ifimm_26_o_14;
output 	idex_ifnext_pc_o_19;
output 	idex_ifnext_pc_o_18;
output 	idex_ifimm_26_o_17;
output 	idex_ifimm_26_o_16;
output 	idex_ifnext_pc_o_21;
output 	idex_ifnext_pc_o_20;
output 	idex_ifimm_26_o_19;
output 	idex_ifimm_26_o_18;
output 	idex_ifnext_pc_o_23;
output 	idex_ifnext_pc_o_22;
output 	idex_ifimm_26_o_21;
output 	idex_ifimm_26_o_20;
output 	idex_ifnext_pc_o_25;
output 	idex_ifnext_pc_o_24;
output 	idex_ifimm_26_o_23;
output 	idex_ifimm_26_o_22;
output 	idex_ifnext_pc_o_27;
output 	idex_ifnext_pc_o_26;
output 	idex_ifimm_26_o_25;
output 	idex_ifimm_26_o_24;
output 	idex_ifnext_pc_o_29;
output 	idex_ifnext_pc_o_28;
output 	idex_ifnext_pc_o_31;
output 	idex_ifnext_pc_o_30;
output 	idex_ifhalt_o;
input 	ifid_ifinstr_o_26;
input 	ifid_ifinstr_o_31;
input 	ifid_ifinstr_o_27;
input 	ifid_ifinstr_o_28;
input 	ifid_ifinstr_o_30;
input 	ifid_ifinstr_o_5;
input 	ifid_ifinstr_o_4;
input 	always0;
input 	ifid_ifinstr_o_29;
input 	ifid_ifinstr_o_1;
input 	ifid_ifinstr_o_3;
input 	ifid_ifinstr_o_2;
output 	idex_ifRegDest_o_1;
output 	idex_ifrd_o_1;
output 	idex_ifRegDest_o_0;
output 	idex_ifrd_o_0;
output 	idex_ifrd_o_3;
output 	idex_ifrd_o_2;
output 	idex_ifregWEN_o;
output 	idex_ifrd_o_4;
input 	cuifregWEN;
input 	Equal0;
input 	ifid_ifinstr_o_0;
input 	Equal3;
input 	Equal2;
output 	idex_ifjal_o;
output 	idex_iflui_o;
output 	idex_ifmemToReg_o;
input 	ifid_ifinstr_o_7;
input 	Mux62;
input 	Mux621;
input 	Mux30;
input 	Mux301;
input 	ifid_ifinstr_o_6;
input 	Mux63;
input 	Mux631;
input 	Mux31;
input 	Mux311;
input 	Equal10;
input 	Mux29;
input 	Mux291;
input 	Mux27;
input 	Mux271;
input 	Mux28;
input 	Mux281;
input 	ifid_ifinstr_o_8;
input 	Mux61;
input 	Mux611;
input 	Mux23;
input 	Mux231;
input 	Mux24;
input 	Mux241;
input 	Mux25;
input 	Mux251;
input 	Mux26;
input 	Mux261;
input 	Mux60;
input 	Mux601;
input 	ifid_ifinstr_o_9;
input 	Mux15;
input 	Mux151;
input 	Mux16;
input 	Mux161;
input 	Mux17;
input 	Mux171;
input 	Mux18;
input 	Mux181;
input 	Mux19;
input 	Mux191;
input 	Mux20;
input 	Mux201;
input 	Mux21;
input 	Mux211;
input 	Mux22;
input 	Mux221;
input 	Mux59;
input 	Mux591;
input 	ifid_ifinstr_o_10;
input 	Mux0;
input 	Mux01;
input 	Mux2;
input 	Mux210;
input 	Mux1;
input 	Mux11;
input 	Mux3;
input 	Mux32;
input 	Mux5;
input 	Mux51;
input 	Mux4;
input 	Mux41;
input 	Mux6;
input 	Mux64;
input 	Mux7;
input 	Mux71;
input 	Mux9;
input 	Mux91;
input 	Mux8;
input 	Mux81;
input 	Mux10;
input 	Mux101;
input 	Mux111;
input 	Mux112;
input 	Mux13;
input 	Mux131;
input 	Mux12;
input 	Mux121;
input 	Mux14;
input 	Mux141;
input 	ifid_ifinstr_o_15;
input 	Mux321;
input 	Mux322;
input 	Mux47;
input 	Mux471;
input 	Mux46;
input 	Mux461;
input 	Mux45;
input 	Mux451;
input 	Mux44;
input 	Mux441;
input 	Mux43;
input 	Mux431;
input 	Mux42;
input 	Mux421;
input 	Mux411;
input 	Mux412;
input 	Mux40;
input 	Mux401;
input 	Mux39;
input 	Mux391;
input 	Mux38;
input 	Mux381;
input 	Mux37;
input 	Mux371;
input 	Mux58;
input 	Mux581;
input 	Mux57;
input 	Mux571;
input 	Mux56;
input 	Mux561;
input 	Mux55;
input 	Mux551;
input 	Mux36;
input 	Mux361;
input 	Mux35;
input 	Mux351;
input 	Mux34;
input 	Mux341;
input 	Mux33;
input 	Mux331;
input 	Mux54;
input 	Mux541;
input 	Mux49;
input 	Mux491;
input 	ifid_ifinstr_o_14;
input 	Mux48;
input 	Mux481;
input 	Mux53;
input 	Mux531;
input 	Mux52;
input 	Mux521;
input 	ifid_ifinstr_o_11;
input 	Mux511;
input 	Mux512;
input 	ifid_ifinstr_o_12;
input 	Mux50;
input 	Mux501;
input 	ifid_ifinstr_o_13;
input 	Equal14;
input 	Equal21;
input 	Equal01;
input 	ifid_ifnext_pc_o_1;
input 	Equal5;
input 	ifid_ifnext_pc_o_0;
input 	ifid_ifnext_pc_o_3;
input 	ifid_ifnext_pc_o_2;
input 	ifid_ifnext_pc_o_5;
input 	ifid_ifnext_pc_o_4;
input 	ifid_ifnext_pc_o_7;
input 	ifid_ifnext_pc_o_6;
input 	ifid_ifnext_pc_o_9;
input 	ifid_ifnext_pc_o_8;
input 	ifid_ifnext_pc_o_11;
input 	ifid_ifnext_pc_o_10;
input 	ifid_ifnext_pc_o_13;
input 	ifid_ifnext_pc_o_12;
input 	ifid_ifnext_pc_o_15;
input 	ifid_ifnext_pc_o_14;
input 	ifid_ifnext_pc_o_17;
input 	ifid_ifnext_pc_o_16;
input 	ifid_ifnext_pc_o_19;
input 	ifid_ifnext_pc_o_18;
input 	ifid_ifnext_pc_o_21;
input 	ifid_ifnext_pc_o_20;
input 	ifid_ifnext_pc_o_23;
input 	ifid_ifnext_pc_o_22;
input 	ifid_ifnext_pc_o_25;
input 	ifid_ifnext_pc_o_24;
input 	ifid_ifnext_pc_o_27;
input 	ifid_ifnext_pc_o_26;
input 	ifid_ifnext_pc_o_29;
input 	ifid_ifnext_pc_o_28;
input 	ifid_ifnext_pc_o_31;
input 	ifid_ifnext_pc_o_30;
input 	cuifregWEN1;
input 	Equal1;
input 	CPUCLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \aluop_o~1_combout ;
wire \aluop_o~7_combout ;
wire \aluop_o~10_combout ;
wire \aluop_o~11_combout ;
wire \aluop_o~15_combout ;
wire \aluop_o~0_combout ;
wire \always0~0_combout ;
wire \aluop_o~2_combout ;
wire \aluop_o~3_combout ;
wire \aluop_o~4_combout ;
wire \aluop_o~5_combout ;
wire \idex_if.rt_o[4]~0_combout ;
wire \imm_26_o~0_combout ;
wire \imm_26_o~1_combout ;
wire \imm_26_o~2_combout ;
wire \imm_26_o~3_combout ;
wire \imm_26_o~4_combout ;
wire \idex_if.rt_o[4]~feeder_combout ;
wire \ALUSel_o~0_combout ;
wire \ALUSel_o~1_combout ;
wire \ALUSel_o~3_combout ;
wire \ALUSel_o~2_combout ;
wire \ALUSel_o~4_combout ;
wire \imm_o~0_combout ;
wire \imm_o~1_combout ;
wire \rdat2_o~0_combout ;
wire \rdat2_o~1_combout ;
wire \rdat1_o~0_combout ;
wire \rdat1_o~1_combout ;
wire \imm_26_o~5_combout ;
wire \idex_if.rs_o[1]~feeder_combout ;
wire \imm_26_o~6_combout ;
wire \imm_26_o~7_combout ;
wire \imm_26_o~8_combout ;
wire \idex_if.rs_o[2]~feeder_combout ;
wire \imm_26_o~9_combout ;
wire \idex_if.rs_o[4]~feeder_combout ;
wire \imm_o~2_combout ;
wire \imm_o~3_combout ;
wire \rdat2_o~2_combout ;
wire \rdat2_o~3_combout ;
wire \rdat1_o~2_combout ;
wire \rdat1_o~3_combout ;
wire \aluop_o~8_combout ;
wire \aluop_o~6_combout ;
wire \aluop_o~9_combout ;
wire \rdat1_o~4_combout ;
wire \rdat1_o~5_combout ;
wire \rdat1_o~6_combout ;
wire \rdat1_o~7_combout ;
wire \rdat1_o~8_combout ;
wire \rdat1_o~9_combout ;
wire \imm_o~4_combout ;
wire \idex_if.imm_o[2]~feeder_combout ;
wire \imm_o~5_combout ;
wire \idex_if.shamt_o[2]~feeder_combout ;
wire \rdat2_o~4_combout ;
wire \rdat2_o~5_combout ;
wire \rdat1_o~10_combout ;
wire \rdat1_o~11_combout ;
wire \rdat1_o~12_combout ;
wire \rdat1_o~13_combout ;
wire \rdat1_o~14_combout ;
wire \rdat1_o~15_combout ;
wire \rdat1_o~16_combout ;
wire \rdat1_o~17_combout ;
wire \rdat2_o~6_combout ;
wire \rdat2_o~7_combout ;
wire \imm_o~6_combout ;
wire \imm_o~7_combout ;
wire \rdat1_o~18_combout ;
wire \rdat1_o~19_combout ;
wire \rdat1_o~20_combout ;
wire \rdat1_o~21_combout ;
wire \rdat1_o~22_combout ;
wire \rdat1_o~23_combout ;
wire \rdat1_o~24_combout ;
wire \rdat1_o~25_combout ;
wire \rdat1_o~26_combout ;
wire \rdat1_o~27_combout ;
wire \rdat1_o~28_combout ;
wire \rdat1_o~29_combout ;
wire \rdat1_o~30_combout ;
wire \rdat1_o~31_combout ;
wire \rdat1_o~32_combout ;
wire \rdat1_o~33_combout ;
wire \rdat2_o~8_combout ;
wire \rdat2_o~9_combout ;
wire \imm_o~8_combout ;
wire \imm_o~9_combout ;
wire \rdat1_o~34_combout ;
wire \rdat1_o~35_combout ;
wire \rdat1_o~36_combout ;
wire \rdat1_o~37_combout ;
wire \rdat1_o~38_combout ;
wire \rdat1_o~39_combout ;
wire \rdat1_o~40_combout ;
wire \rdat1_o~41_combout ;
wire \rdat1_o~42_combout ;
wire \rdat1_o~43_combout ;
wire \rdat1_o~44_combout ;
wire \rdat1_o~45_combout ;
wire \rdat1_o~46_combout ;
wire \rdat1_o~47_combout ;
wire \rdat1_o~48_combout ;
wire \rdat1_o~49_combout ;
wire \rdat1_o~50_combout ;
wire \rdat1_o~51_combout ;
wire \rdat1_o~52_combout ;
wire \rdat1_o~53_combout ;
wire \rdat1_o~54_combout ;
wire \rdat1_o~55_combout ;
wire \rdat1_o~56_combout ;
wire \rdat1_o~57_combout ;
wire \rdat1_o~58_combout ;
wire \rdat1_o~59_combout ;
wire \rdat1_o~60_combout ;
wire \rdat1_o~61_combout ;
wire \rdat1_o~62_combout ;
wire \rdat1_o~63_combout ;
wire \imm_o~10_combout ;
wire \idex_if.imm_o[15]~feeder_combout ;
wire \rdat2_o~10_combout ;
wire \rdat2_o~11_combout ;
wire \rdat2_o~12_combout ;
wire \rdat2_o~13_combout ;
wire \rdat2_o~14_combout ;
wire \rdat2_o~15_combout ;
wire \rdat2_o~16_combout ;
wire \rdat2_o~17_combout ;
wire \rdat2_o~18_combout ;
wire \rdat2_o~19_combout ;
wire \rdat2_o~20_combout ;
wire \rdat2_o~21_combout ;
wire \rdat2_o~22_combout ;
wire \rdat2_o~23_combout ;
wire \rdat2_o~24_combout ;
wire \rdat2_o~25_combout ;
wire \rdat2_o~26_combout ;
wire \rdat2_o~27_combout ;
wire \rdat2_o~28_combout ;
wire \rdat2_o~29_combout ;
wire \rdat2_o~30_combout ;
wire \rdat2_o~31_combout ;
wire \rdat2_o~32_combout ;
wire \rdat2_o~33_combout ;
wire \rdat2_o~34_combout ;
wire \rdat2_o~35_combout ;
wire \imm_o~11_combout ;
wire \rdat2_o~36_combout ;
wire \rdat2_o~37_combout ;
wire \rdat2_o~38_combout ;
wire \rdat2_o~39_combout ;
wire \rdat2_o~40_combout ;
wire \rdat2_o~41_combout ;
wire \rdat2_o~42_combout ;
wire \rdat2_o~43_combout ;
wire \rdat2_o~44_combout ;
wire \rdat2_o~45_combout ;
wire \rdat2_o~46_combout ;
wire \rdat2_o~47_combout ;
wire \rdat2_o~48_combout ;
wire \rdat2_o~49_combout ;
wire \rdat2_o~50_combout ;
wire \rdat2_o~51_combout ;
wire \rdat2_o~52_combout ;
wire \rdat2_o~53_combout ;
wire \imm_o~12_combout ;
wire \idex_if.imm_o[14]~feeder_combout ;
wire \rdat2_o~54_combout ;
wire \rdat2_o~55_combout ;
wire \rdat2_o~56_combout ;
wire \rdat2_o~57_combout ;
wire \rdat2_o~58_combout ;
wire \rdat2_o~59_combout ;
wire \imm_o~13_combout ;
wire \idex_if.imm_o[11]~feeder_combout ;
wire \rdat2_o~60_combout ;
wire \rdat2_o~61_combout ;
wire \imm_o~14_combout ;
wire \rdat2_o~62_combout ;
wire \rdat2_o~63_combout ;
wire \imm_o~15_combout ;
wire \aluop_o~12_combout ;
wire \aluop_o~13_combout ;
wire \aluop_o~14_combout ;
wire \aluop_o~16_combout ;
wire \aluop_o~17_combout ;
wire \aluop_o~18_combout ;
wire \aluop_o~19_combout ;
wire \aluop_o~20_combout ;
wire \instr_o~0_combout ;
wire \dWEN_o~0_combout ;
wire \dREN_o~0_combout ;
wire \next_pc_o~0_combout ;
wire \jumpSel_o~2_combout ;
wire \jumpSel_o~3_combout ;
wire \bne_o~0_combout ;
wire \jumpSel_o~5_combout ;
wire \jumpSel_o~4_combout ;
wire \instr_o~1_combout ;
wire \instr_o~2_combout ;
wire \instr_o~3_combout ;
wire \instr_o~4_combout ;
wire \bne_o~1_combout ;
wire \PCSel_o~0_combout ;
wire \PCSel_o~1_combout ;
wire \next_pc_o~1_combout ;
wire \next_pc_o~2_combout ;
wire \next_pc_o~3_combout ;
wire \next_pc_o~4_combout ;
wire \next_pc_o~5_combout ;
wire \next_pc_o~6_combout ;
wire \next_pc_o~7_combout ;
wire \next_pc_o~8_combout ;
wire \next_pc_o~9_combout ;
wire \next_pc_o~10_combout ;
wire \next_pc_o~11_combout ;
wire \next_pc_o~12_combout ;
wire \next_pc_o~13_combout ;
wire \next_pc_o~14_combout ;
wire \next_pc_o~15_combout ;
wire \next_pc_o~16_combout ;
wire \next_pc_o~17_combout ;
wire \next_pc_o~18_combout ;
wire \next_pc_o~19_combout ;
wire \next_pc_o~20_combout ;
wire \next_pc_o~21_combout ;
wire \next_pc_o~22_combout ;
wire \next_pc_o~23_combout ;
wire \next_pc_o~24_combout ;
wire \next_pc_o~25_combout ;
wire \next_pc_o~26_combout ;
wire \next_pc_o~27_combout ;
wire \next_pc_o~28_combout ;
wire \next_pc_o~29_combout ;
wire \next_pc_o~30_combout ;
wire \next_pc_o~31_combout ;
wire \lui_o~2_combout ;
wire \halt_o~0_combout ;
wire \RegDest_o~0_combout ;
wire \RegDest_o~1_combout ;
wire \idex_if.rd_o[1]~feeder_combout ;
wire \RegDest_o~2_combout ;
wire \RegDest_o~3_combout ;
wire \idex_if.rd_o[2]~feeder_combout ;
wire \regWEN_o~0_combout ;
wire \jal_o~0_combout ;
wire \lui_o~3_combout ;


// Location: LCCOMB_X60_Y26_N30
cycloneive_lcell_comb \aluop_o~1 (
// Equation(s):
// \aluop_o~1_combout  = (ifid_ifinstr_o_27 & (((ifid_ifinstr_o_29)))) # (!ifid_ifinstr_o_27 & ((ifid_ifinstr_o_28 & ((!ifid_ifinstr_o_29))) # (!ifid_ifinstr_o_28 & ((always0) # (ifid_ifinstr_o_29)))))

	.dataa(always0),
	.datab(ifid_ifinstr_o_27),
	.datac(ifid_ifinstr_o_28),
	.datad(ifid_ifinstr_o_29),
	.cin(gnd),
	.combout(\aluop_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~1 .lut_mask = 16'hCF32;
defparam \aluop_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N10
cycloneive_lcell_comb \aluop_o~7 (
// Equation(s):
// \aluop_o~7_combout  = (((ifid_ifinstr_o_2) # (!ifid_ifinstr_o_0)) # (!ifid_ifinstr_o_1)) # (!ifid_ifinstr_o_5)

	.dataa(ifid_ifinstr_o_5),
	.datab(ifid_ifinstr_o_1),
	.datac(ifid_ifinstr_o_2),
	.datad(ifid_ifinstr_o_0),
	.cin(gnd),
	.combout(\aluop_o~7_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~7 .lut_mask = 16'hF7FF;
defparam \aluop_o~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N12
cycloneive_lcell_comb \aluop_o~10 (
// Equation(s):
// \aluop_o~10_combout  = (ifid_ifinstr_o_2 & (ifid_ifinstr_o_5 & ((ifid_ifinstr_o_0)))) # (!ifid_ifinstr_o_2 & (ifid_ifinstr_o_1 & ((ifid_ifinstr_o_5) # (!ifid_ifinstr_o_0))))

	.dataa(ifid_ifinstr_o_5),
	.datab(ifid_ifinstr_o_1),
	.datac(ifid_ifinstr_o_2),
	.datad(ifid_ifinstr_o_0),
	.cin(gnd),
	.combout(\aluop_o~10_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~10 .lut_mask = 16'hA80C;
defparam \aluop_o~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N22
cycloneive_lcell_comb \aluop_o~11 (
// Equation(s):
// \aluop_o~11_combout  = (ifid_ifinstr_o_3 & (ifid_ifinstr_o_0 & (Equal14))) # (!ifid_ifinstr_o_3 & (((\aluop_o~10_combout ))))

	.dataa(ifid_ifinstr_o_0),
	.datab(Equal14),
	.datac(ifid_ifinstr_o_3),
	.datad(\aluop_o~10_combout ),
	.cin(gnd),
	.combout(\aluop_o~11_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~11 .lut_mask = 16'h8F80;
defparam \aluop_o~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N30
cycloneive_lcell_comb \aluop_o~15 (
// Equation(s):
// \aluop_o~15_combout  = (!Equal10 & ((ifid_ifinstr_o_3) # ((ifid_ifinstr_o_2) # (!always0))))

	.dataa(ifid_ifinstr_o_3),
	.datab(Equal10),
	.datac(ifid_ifinstr_o_2),
	.datad(always0),
	.cin(gnd),
	.combout(\aluop_o~15_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~15 .lut_mask = 16'h3233;
defparam \aluop_o~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y31_N17
dffeas \idex_if.aluop_o[1] (
	.clk(CPUCLK),
	.d(\aluop_o~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifaluop_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.aluop_o[1] .is_wysiwyg = "true";
defparam \idex_if.aluop_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N27
dffeas \idex_if.rt_o[0] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_26_o~0_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrt_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rt_o[0] .is_wysiwyg = "true";
defparam \idex_if.rt_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N29
dffeas \idex_if.rt_o[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_26_o~1_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrt_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rt_o[1] .is_wysiwyg = "true";
defparam \idex_if.rt_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N25
dffeas \idex_if.rt_o[2] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_26_o~2_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrt_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rt_o[2] .is_wysiwyg = "true";
defparam \idex_if.rt_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N31
dffeas \idex_if.rt_o[3] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_26_o~3_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrt_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rt_o[3] .is_wysiwyg = "true";
defparam \idex_if.rt_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N19
dffeas \idex_if.rt_o[4] (
	.clk(CPUCLK),
	.d(\idex_if.rt_o[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrt_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rt_o[4] .is_wysiwyg = "true";
defparam \idex_if.rt_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N11
dffeas \idex_if.ALUSel_o[1] (
	.clk(CPUCLK),
	.d(\ALUSel_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifALUSel_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.ALUSel_o[1] .is_wysiwyg = "true";
defparam \idex_if.ALUSel_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N17
dffeas \idex_if.ALUSel_o[0] (
	.clk(CPUCLK),
	.d(\ALUSel_o~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifALUSel_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.ALUSel_o[0] .is_wysiwyg = "true";
defparam \idex_if.ALUSel_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N9
dffeas \idex_if.imm_o[1] (
	.clk(CPUCLK),
	.d(\imm_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_o[1] .is_wysiwyg = "true";
defparam \idex_if.imm_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N3
dffeas \idex_if.shamt_o[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~1_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifshamt_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.shamt_o[1] .is_wysiwyg = "true";
defparam \idex_if.shamt_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N25
dffeas \idex_if.rdat2_o[1] (
	.clk(CPUCLK),
	.d(\rdat2_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[1] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N5
dffeas \idex_if.rdat1_o[1] (
	.clk(CPUCLK),
	.d(\rdat1_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[1] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N5
dffeas \idex_if.rs_o[1] (
	.clk(CPUCLK),
	.d(\idex_if.rs_o[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrs_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rs_o[1] .is_wysiwyg = "true";
defparam \idex_if.rs_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N31
dffeas \idex_if.rs_o[0] (
	.clk(CPUCLK),
	.d(\imm_26_o~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrs_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rs_o[0] .is_wysiwyg = "true";
defparam \idex_if.rs_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N9
dffeas \idex_if.rs_o[3] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_26_o~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrs_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rs_o[3] .is_wysiwyg = "true";
defparam \idex_if.rs_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N21
dffeas \idex_if.rs_o[2] (
	.clk(CPUCLK),
	.d(\idex_if.rs_o[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrs_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rs_o[2] .is_wysiwyg = "true";
defparam \idex_if.rs_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N7
dffeas \idex_if.rs_o[4] (
	.clk(CPUCLK),
	.d(\idex_if.rs_o[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrs_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rs_o[4] .is_wysiwyg = "true";
defparam \idex_if.rs_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N21
dffeas \idex_if.imm_o[0] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~2_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_o[0] .is_wysiwyg = "true";
defparam \idex_if.imm_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N1
dffeas \idex_if.shamt_o[0] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~3_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifshamt_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.shamt_o[0] .is_wysiwyg = "true";
defparam \idex_if.shamt_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N9
dffeas \idex_if.rdat2_o[0] (
	.clk(CPUCLK),
	.d(\rdat2_o~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[0] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y31_N25
dffeas \idex_if.rdat1_o[0] (
	.clk(CPUCLK),
	.d(\rdat1_o~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[0] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N19
dffeas \idex_if.aluop_o[2] (
	.clk(CPUCLK),
	.d(\aluop_o~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifaluop_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.aluop_o[2] .is_wysiwyg = "true";
defparam \idex_if.aluop_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N29
dffeas \idex_if.rdat1_o[2] (
	.clk(CPUCLK),
	.d(\rdat1_o~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[2] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N15
dffeas \idex_if.rdat1_o[4] (
	.clk(CPUCLK),
	.d(\rdat1_o~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[4] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N13
dffeas \idex_if.rdat1_o[3] (
	.clk(CPUCLK),
	.d(\rdat1_o~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[3] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N7
dffeas \idex_if.imm_o[2] (
	.clk(CPUCLK),
	.d(\idex_if.imm_o[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_o[2] .is_wysiwyg = "true";
defparam \idex_if.imm_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N25
dffeas \idex_if.shamt_o[2] (
	.clk(CPUCLK),
	.d(\idex_if.shamt_o[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifshamt_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.shamt_o[2] .is_wysiwyg = "true";
defparam \idex_if.shamt_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N1
dffeas \idex_if.rdat2_o[2] (
	.clk(CPUCLK),
	.d(\rdat2_o~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[2] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y30_N1
dffeas \idex_if.rdat1_o[8] (
	.clk(CPUCLK),
	.d(\rdat1_o~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_8),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[8] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y30_N3
dffeas \idex_if.rdat1_o[7] (
	.clk(CPUCLK),
	.d(\rdat1_o~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_7),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[7] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N21
dffeas \idex_if.rdat1_o[6] (
	.clk(CPUCLK),
	.d(\rdat1_o~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_6),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[6] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N7
dffeas \idex_if.rdat1_o[5] (
	.clk(CPUCLK),
	.d(\rdat1_o~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_5),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[5] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N7
dffeas \idex_if.rdat2_o[3] (
	.clk(CPUCLK),
	.d(\rdat2_o~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[3] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y27_N1
dffeas \idex_if.imm_o[3] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~6_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_o[3] .is_wysiwyg = "true";
defparam \idex_if.imm_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N7
dffeas \idex_if.shamt_o[3] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifshamt_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.shamt_o[3] .is_wysiwyg = "true";
defparam \idex_if.shamt_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y28_N25
dffeas \idex_if.rdat1_o[16] (
	.clk(CPUCLK),
	.d(\rdat1_o~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_16),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[16] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N11
dffeas \idex_if.rdat1_o[15] (
	.clk(CPUCLK),
	.d(\rdat1_o~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_15),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[15] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y28_N19
dffeas \idex_if.rdat1_o[14] (
	.clk(CPUCLK),
	.d(\rdat1_o~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_14),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[14] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N7
dffeas \idex_if.rdat1_o[13] (
	.clk(CPUCLK),
	.d(\rdat1_o~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_13),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[13] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y32_N1
dffeas \idex_if.rdat1_o[12] (
	.clk(CPUCLK),
	.d(\rdat1_o~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_12),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[12] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y32_N31
dffeas \idex_if.rdat1_o[11] (
	.clk(CPUCLK),
	.d(\rdat1_o~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_11),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[11] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y31_N25
dffeas \idex_if.rdat1_o[10] (
	.clk(CPUCLK),
	.d(\rdat1_o~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_10),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[10] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N25
dffeas \idex_if.rdat1_o[9] (
	.clk(CPUCLK),
	.d(\rdat1_o~33_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_9),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[9] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N13
dffeas \idex_if.rdat2_o[4] (
	.clk(CPUCLK),
	.d(\rdat2_o~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[4] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N25
dffeas \idex_if.imm_o[4] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_o[4] .is_wysiwyg = "true";
defparam \idex_if.imm_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N11
dffeas \idex_if.shamt_o[4] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifshamt_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.shamt_o[4] .is_wysiwyg = "true";
defparam \idex_if.shamt_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y27_N1
dffeas \idex_if.rdat1_o[31] (
	.clk(CPUCLK),
	.d(\rdat1_o~35_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_31),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[31] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y27_N15
dffeas \idex_if.rdat1_o[29] (
	.clk(CPUCLK),
	.d(\rdat1_o~37_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_29),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[29] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N9
dffeas \idex_if.rdat1_o[30] (
	.clk(CPUCLK),
	.d(\rdat1_o~39_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_30),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[30] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N19
dffeas \idex_if.rdat1_o[28] (
	.clk(CPUCLK),
	.d(\rdat1_o~41_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_28),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[28] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N19
dffeas \idex_if.rdat1_o[26] (
	.clk(CPUCLK),
	.d(\rdat1_o~43_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_26),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[26] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N21
dffeas \idex_if.rdat1_o[27] (
	.clk(CPUCLK),
	.d(\rdat1_o~45_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_27),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[27] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N29
dffeas \idex_if.rdat1_o[25] (
	.clk(CPUCLK),
	.d(\rdat1_o~47_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_25),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[25] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N1
dffeas \idex_if.rdat1_o[24] (
	.clk(CPUCLK),
	.d(\rdat1_o~49_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_24),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[24] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N9
dffeas \idex_if.rdat1_o[22] (
	.clk(CPUCLK),
	.d(\rdat1_o~51_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_22),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[22] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N31
dffeas \idex_if.rdat1_o[23] (
	.clk(CPUCLK),
	.d(\rdat1_o~53_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_23),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[23] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N13
dffeas \idex_if.rdat1_o[21] (
	.clk(CPUCLK),
	.d(\rdat1_o~55_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_21),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[21] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y31_N31
dffeas \idex_if.rdat1_o[20] (
	.clk(CPUCLK),
	.d(\rdat1_o~57_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_20),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[20] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y29_N17
dffeas \idex_if.rdat1_o[18] (
	.clk(CPUCLK),
	.d(\rdat1_o~59_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_18),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[18] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y29_N15
dffeas \idex_if.rdat1_o[19] (
	.clk(CPUCLK),
	.d(\rdat1_o~61_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_19),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[19] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y31_N3
dffeas \idex_if.rdat1_o[17] (
	.clk(CPUCLK),
	.d(\rdat1_o~63_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat1_o_17),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat1_o[17] .is_wysiwyg = "true";
defparam \idex_if.rdat1_o[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N29
dffeas \idex_if.imm_o[15] (
	.clk(CPUCLK),
	.d(\idex_if.imm_o[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_o_15),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_o[15] .is_wysiwyg = "true";
defparam \idex_if.imm_o[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y31_N29
dffeas \idex_if.rdat2_o[31] (
	.clk(CPUCLK),
	.d(\rdat2_o~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_31),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[31] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N13
dffeas \idex_if.rdat2_o[16] (
	.clk(CPUCLK),
	.d(\rdat2_o~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_16),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[16] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y27_N21
dffeas \idex_if.rdat2_o[17] (
	.clk(CPUCLK),
	.d(\rdat2_o~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_17),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[17] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y27_N25
dffeas \idex_if.rdat2_o[18] (
	.clk(CPUCLK),
	.d(\rdat2_o~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_18),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[18] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N1
dffeas \idex_if.rdat2_o[19] (
	.clk(CPUCLK),
	.d(\rdat2_o~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_19),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[19] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N21
dffeas \idex_if.rdat2_o[20] (
	.clk(CPUCLK),
	.d(\rdat2_o~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_20),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[20] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N3
dffeas \idex_if.rdat2_o[21] (
	.clk(CPUCLK),
	.d(\rdat2_o~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_21),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[21] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N25
dffeas \idex_if.rdat2_o[22] (
	.clk(CPUCLK),
	.d(\rdat2_o~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_22),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[22] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N11
dffeas \idex_if.rdat2_o[23] (
	.clk(CPUCLK),
	.d(\rdat2_o~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_23),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[23] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N31
dffeas \idex_if.rdat2_o[24] (
	.clk(CPUCLK),
	.d(\rdat2_o~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_24),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[24] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N17
dffeas \idex_if.rdat2_o[25] (
	.clk(CPUCLK),
	.d(\rdat2_o~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_25),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[25] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N13
dffeas \idex_if.rdat2_o[26] (
	.clk(CPUCLK),
	.d(\rdat2_o~33_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_26),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[26] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y28_N1
dffeas \idex_if.rdat2_o[5] (
	.clk(CPUCLK),
	.d(\rdat2_o~35_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_5),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[5] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y36_N27
dffeas \idex_if.imm_o[5] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~11_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_o_5),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_o[5] .is_wysiwyg = "true";
defparam \idex_if.imm_o[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y28_N15
dffeas \idex_if.rdat2_o[6] (
	.clk(CPUCLK),
	.d(\rdat2_o~37_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_6),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[6] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N29
dffeas \idex_if.imm_o[6] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~3_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_o_6),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_o[6] .is_wysiwyg = "true";
defparam \idex_if.imm_o[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y29_N5
dffeas \idex_if.rdat2_o[7] (
	.clk(CPUCLK),
	.d(\rdat2_o~39_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_7),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[7] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N15
dffeas \idex_if.imm_o[7] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~1_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_o_7),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_o[7] .is_wysiwyg = "true";
defparam \idex_if.imm_o[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y29_N3
dffeas \idex_if.rdat2_o[8] (
	.clk(CPUCLK),
	.d(\rdat2_o~41_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_8),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[8] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N11
dffeas \idex_if.imm_o[8] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~5_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_o_8),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_o[8] .is_wysiwyg = "true";
defparam \idex_if.imm_o[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N23
dffeas \idex_if.rdat2_o[27] (
	.clk(CPUCLK),
	.d(\rdat2_o~43_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_27),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[27] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N7
dffeas \idex_if.rdat2_o[28] (
	.clk(CPUCLK),
	.d(\rdat2_o~45_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_28),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[28] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N21
dffeas \idex_if.rdat2_o[29] (
	.clk(CPUCLK),
	.d(\rdat2_o~47_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_29),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[29] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N23
dffeas \idex_if.rdat2_o[30] (
	.clk(CPUCLK),
	.d(\rdat2_o~49_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_30),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[30] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N17
dffeas \idex_if.rdat2_o[9] (
	.clk(CPUCLK),
	.d(\rdat2_o~51_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_9),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[9] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N11
dffeas \idex_if.imm_o[9] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~7_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_o_9),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_o[9] .is_wysiwyg = "true";
defparam \idex_if.imm_o[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N11
dffeas \idex_if.rdat2_o[14] (
	.clk(CPUCLK),
	.d(\rdat2_o~53_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_14),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[14] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N25
dffeas \idex_if.imm_o[14] (
	.clk(CPUCLK),
	.d(\idex_if.imm_o[14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_o_14),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_o[14] .is_wysiwyg = "true";
defparam \idex_if.imm_o[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N27
dffeas \idex_if.rdat2_o[15] (
	.clk(CPUCLK),
	.d(\rdat2_o~55_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_15),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[15] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y32_N13
dffeas \idex_if.rdat2_o[10] (
	.clk(CPUCLK),
	.d(\rdat2_o~57_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_10),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[10] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N5
dffeas \idex_if.imm_o[10] (
	.clk(CPUCLK),
	.d(\imm_o~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_o_10),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_o[10] .is_wysiwyg = "true";
defparam \idex_if.imm_o[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N1
dffeas \idex_if.rdat2_o[11] (
	.clk(CPUCLK),
	.d(\rdat2_o~59_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_11),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[11] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N15
dffeas \idex_if.imm_o[11] (
	.clk(CPUCLK),
	.d(\idex_if.imm_o[11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_o_11),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_o[11] .is_wysiwyg = "true";
defparam \idex_if.imm_o[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N23
dffeas \idex_if.rdat2_o[12] (
	.clk(CPUCLK),
	.d(\rdat2_o~61_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_12),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[12] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N5
dffeas \idex_if.imm_o[12] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~14_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_o_12),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_o[12] .is_wysiwyg = "true";
defparam \idex_if.imm_o[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N25
dffeas \idex_if.rdat2_o[13] (
	.clk(CPUCLK),
	.d(\rdat2_o~63_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrdat2_o_13),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rdat2_o[13] .is_wysiwyg = "true";
defparam \idex_if.rdat2_o[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N29
dffeas \idex_if.imm_o[13] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~15_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_o_13),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_o[13] .is_wysiwyg = "true";
defparam \idex_if.imm_o[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N19
dffeas \idex_if.aluop_o[0] (
	.clk(CPUCLK),
	.d(\aluop_o~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifaluop_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.aluop_o[0] .is_wysiwyg = "true";
defparam \idex_if.aluop_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y27_N15
dffeas \idex_if.aluop_o[3] (
	.clk(CPUCLK),
	.d(\aluop_o~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifaluop_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.aluop_o[3] .is_wysiwyg = "true";
defparam \idex_if.aluop_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N27
dffeas \idex_if.dWEN_o (
	.clk(CPUCLK),
	.d(\dWEN_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifdWEN_o),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.dWEN_o .is_wysiwyg = "true";
defparam \idex_if.dWEN_o .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N9
dffeas \idex_if.dREN_o (
	.clk(CPUCLK),
	.d(\dREN_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifdREN_o),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.dREN_o .is_wysiwyg = "true";
defparam \idex_if.dREN_o .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y28_N13
dffeas \idex_if.next_pc_o[1] (
	.clk(CPUCLK),
	.d(\next_pc_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[1] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y27_N17
dffeas \idex_if.jumpSel_o[1] (
	.clk(CPUCLK),
	.d(\jumpSel_o~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifjumpSel_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.jumpSel_o[1] .is_wysiwyg = "true";
defparam \idex_if.jumpSel_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N27
dffeas \idex_if.jumpSel_o[0] (
	.clk(CPUCLK),
	.d(\jumpSel_o~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifjumpSel_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.jumpSel_o[0] .is_wysiwyg = "true";
defparam \idex_if.jumpSel_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y27_N1
dffeas \idex_if.instr_o[31] (
	.clk(CPUCLK),
	.d(\instr_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifinstr_o_31),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.instr_o[31] .is_wysiwyg = "true";
defparam \idex_if.instr_o[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N23
dffeas \idex_if.instr_o[30] (
	.clk(CPUCLK),
	.d(\instr_o~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifinstr_o_30),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.instr_o[30] .is_wysiwyg = "true";
defparam \idex_if.instr_o[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N19
dffeas \idex_if.instr_o[27] (
	.clk(CPUCLK),
	.d(\instr_o~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifinstr_o_27),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.instr_o[27] .is_wysiwyg = "true";
defparam \idex_if.instr_o[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N17
dffeas \idex_if.instr_o[26] (
	.clk(CPUCLK),
	.d(\instr_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifinstr_o_26),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.instr_o[26] .is_wysiwyg = "true";
defparam \idex_if.instr_o[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N15
dffeas \idex_if.instr_o[28] (
	.clk(CPUCLK),
	.d(\instr_o~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifinstr_o_28),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.instr_o[28] .is_wysiwyg = "true";
defparam \idex_if.instr_o[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N1
dffeas \idex_if.bne_o (
	.clk(CPUCLK),
	.d(\bne_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifbne_o),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.bne_o .is_wysiwyg = "true";
defparam \idex_if.bne_o .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y27_N21
dffeas \idex_if.PCSel_o (
	.clk(CPUCLK),
	.d(\PCSel_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifPCSel_o),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.PCSel_o .is_wysiwyg = "true";
defparam \idex_if.PCSel_o .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y32_N25
dffeas \idex_if.next_pc_o[0] (
	.clk(CPUCLK),
	.d(\next_pc_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[0] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N27
dffeas \idex_if.next_pc_o[3] (
	.clk(CPUCLK),
	.d(\next_pc_o~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[3] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N13
dffeas \idex_if.next_pc_o[2] (
	.clk(CPUCLK),
	.d(\next_pc_o~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[2] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N21
dffeas \idex_if.imm_26_o[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~0_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[1] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N31
dffeas \idex_if.imm_26_o[0] (
	.clk(CPUCLK),
	.d(\imm_o~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[0] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N23
dffeas \idex_if.next_pc_o[5] (
	.clk(CPUCLK),
	.d(\next_pc_o~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_5),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[5] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N17
dffeas \idex_if.next_pc_o[4] (
	.clk(CPUCLK),
	.d(\next_pc_o~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[4] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y27_N27
dffeas \idex_if.imm_26_o[3] (
	.clk(CPUCLK),
	.d(\imm_o~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[3] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N17
dffeas \idex_if.imm_26_o[2] (
	.clk(CPUCLK),
	.d(\imm_o~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[2] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y27_N13
dffeas \idex_if.next_pc_o[7] (
	.clk(CPUCLK),
	.d(\next_pc_o~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_7),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[7] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y27_N3
dffeas \idex_if.next_pc_o[6] (
	.clk(CPUCLK),
	.d(\next_pc_o~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_6),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[6] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y36_N23
dffeas \idex_if.imm_26_o[5] (
	.clk(CPUCLK),
	.d(\imm_o~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_5),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[5] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N23
dffeas \idex_if.imm_26_o[4] (
	.clk(CPUCLK),
	.d(\imm_o~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[4] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y29_N29
dffeas \idex_if.next_pc_o[9] (
	.clk(CPUCLK),
	.d(\next_pc_o~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_9),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[9] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y31_N15
dffeas \idex_if.next_pc_o[8] (
	.clk(CPUCLK),
	.d(\next_pc_o~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_8),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[8] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N23
dffeas \idex_if.imm_26_o[7] (
	.clk(CPUCLK),
	.d(\imm_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_7),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[7] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N5
dffeas \idex_if.imm_26_o[6] (
	.clk(CPUCLK),
	.d(\imm_o~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_6),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[6] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N11
dffeas \idex_if.next_pc_o[11] (
	.clk(CPUCLK),
	.d(\next_pc_o~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_11),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[11] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N13
dffeas \idex_if.next_pc_o[10] (
	.clk(CPUCLK),
	.d(\next_pc_o~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_10),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[10] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N27
dffeas \idex_if.imm_26_o[9] (
	.clk(CPUCLK),
	.d(\imm_o~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_9),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[9] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N23
dffeas \idex_if.imm_26_o[8] (
	.clk(CPUCLK),
	.d(\imm_o~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_8),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[8] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N29
dffeas \idex_if.next_pc_o[13] (
	.clk(CPUCLK),
	.d(\next_pc_o~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_13),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[13] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N29
dffeas \idex_if.next_pc_o[12] (
	.clk(CPUCLK),
	.d(\next_pc_o~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_12),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[12] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N21
dffeas \idex_if.imm_26_o[11] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~13_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_11),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[11] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N3
dffeas \idex_if.imm_26_o[10] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~9_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_10),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[10] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N21
dffeas \idex_if.next_pc_o[15] (
	.clk(CPUCLK),
	.d(\next_pc_o~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_15),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[15] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N7
dffeas \idex_if.next_pc_o[14] (
	.clk(CPUCLK),
	.d(\next_pc_o~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_14),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[14] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N1
dffeas \idex_if.imm_26_o[13] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~15_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_13),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[13] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N19
dffeas \idex_if.imm_26_o[12] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~14_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_12),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[12] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N31
dffeas \idex_if.next_pc_o[17] (
	.clk(CPUCLK),
	.d(\next_pc_o~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_17),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[17] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y29_N17
dffeas \idex_if.next_pc_o[16] (
	.clk(CPUCLK),
	.d(\next_pc_o~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_16),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[16] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N27
dffeas \idex_if.imm_26_o[15] (
	.clk(CPUCLK),
	.d(\imm_o~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_15),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[15] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N5
dffeas \idex_if.imm_26_o[14] (
	.clk(CPUCLK),
	.d(\imm_o~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_14),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[14] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y27_N5
dffeas \idex_if.next_pc_o[19] (
	.clk(CPUCLK),
	.d(\next_pc_o~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_19),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[19] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N11
dffeas \idex_if.next_pc_o[18] (
	.clk(CPUCLK),
	.d(\next_pc_o~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_18),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[18] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y31_N21
dffeas \idex_if.imm_26_o[17] (
	.clk(CPUCLK),
	.d(\imm_26_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_17),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[17] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N11
dffeas \idex_if.imm_26_o[16] (
	.clk(CPUCLK),
	.d(\imm_26_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_16),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[16] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N11
dffeas \idex_if.next_pc_o[21] (
	.clk(CPUCLK),
	.d(\next_pc_o~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_21),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[21] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N29
dffeas \idex_if.next_pc_o[20] (
	.clk(CPUCLK),
	.d(\next_pc_o~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_20),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[20] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y31_N7
dffeas \idex_if.imm_26_o[19] (
	.clk(CPUCLK),
	.d(\imm_26_o~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_19),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[19] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N17
dffeas \idex_if.imm_26_o[18] (
	.clk(CPUCLK),
	.d(\imm_26_o~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_18),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[18] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N3
dffeas \idex_if.next_pc_o[23] (
	.clk(CPUCLK),
	.d(\next_pc_o~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_23),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[23] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N27
dffeas \idex_if.next_pc_o[22] (
	.clk(CPUCLK),
	.d(\next_pc_o~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_22),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[22] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N29
dffeas \idex_if.imm_26_o[21] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_26_o~6_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_21),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[21] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N9
dffeas \idex_if.imm_26_o[20] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_26_o~4_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_20),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[20] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N1
dffeas \idex_if.next_pc_o[25] (
	.clk(CPUCLK),
	.d(\next_pc_o~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_25),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[25] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N29
dffeas \idex_if.next_pc_o[24] (
	.clk(CPUCLK),
	.d(\next_pc_o~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_24),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[24] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N11
dffeas \idex_if.imm_26_o[23] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_26_o~8_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_23),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[23] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N3
dffeas \idex_if.imm_26_o[22] (
	.clk(CPUCLK),
	.d(\imm_26_o~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_22),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[22] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N7
dffeas \idex_if.next_pc_o[27] (
	.clk(CPUCLK),
	.d(\next_pc_o~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_27),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[27] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N7
dffeas \idex_if.next_pc_o[26] (
	.clk(CPUCLK),
	.d(\next_pc_o~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_26),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[26] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N25
dffeas \idex_if.imm_26_o[25] (
	.clk(CPUCLK),
	.d(\imm_26_o~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_25),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[25] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N27
dffeas \idex_if.imm_26_o[24] (
	.clk(CPUCLK),
	.d(\imm_26_o~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifimm_26_o_24),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.imm_26_o[24] .is_wysiwyg = "true";
defparam \idex_if.imm_26_o[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N11
dffeas \idex_if.next_pc_o[29] (
	.clk(CPUCLK),
	.d(\next_pc_o~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_29),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[29] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y28_N23
dffeas \idex_if.next_pc_o[28] (
	.clk(CPUCLK),
	.d(\next_pc_o~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_28),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[28] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N21
dffeas \idex_if.next_pc_o[31] (
	.clk(CPUCLK),
	.d(\next_pc_o~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_31),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[31] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N27
dffeas \idex_if.next_pc_o[30] (
	.clk(CPUCLK),
	.d(\next_pc_o~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifnext_pc_o_30),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.next_pc_o[30] .is_wysiwyg = "true";
defparam \idex_if.next_pc_o[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N13
dffeas \idex_if.halt_o (
	.clk(CPUCLK),
	.d(\halt_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifhalt_o),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.halt_o .is_wysiwyg = "true";
defparam \idex_if.halt_o .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N7
dffeas \idex_if.RegDest_o[1] (
	.clk(CPUCLK),
	.d(\RegDest_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifRegDest_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.RegDest_o[1] .is_wysiwyg = "true";
defparam \idex_if.RegDest_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N17
dffeas \idex_if.rd_o[1] (
	.clk(CPUCLK),
	.d(\idex_if.rd_o[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrd_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rd_o[1] .is_wysiwyg = "true";
defparam \idex_if.rd_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y27_N11
dffeas \idex_if.RegDest_o[0] (
	.clk(CPUCLK),
	.d(\RegDest_o~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifRegDest_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.RegDest_o[0] .is_wysiwyg = "true";
defparam \idex_if.RegDest_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N5
dffeas \idex_if.rd_o[0] (
	.clk(CPUCLK),
	.d(\imm_o~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrd_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rd_o[0] .is_wysiwyg = "true";
defparam \idex_if.rd_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N17
dffeas \idex_if.rd_o[3] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~12_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrd_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rd_o[3] .is_wysiwyg = "true";
defparam \idex_if.rd_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N19
dffeas \idex_if.rd_o[2] (
	.clk(CPUCLK),
	.d(\idex_if.rd_o[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrd_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rd_o[2] .is_wysiwyg = "true";
defparam \idex_if.rd_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N11
dffeas \idex_if.regWEN_o (
	.clk(CPUCLK),
	.d(\regWEN_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifregWEN_o),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.regWEN_o .is_wysiwyg = "true";
defparam \idex_if.regWEN_o .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N9
dffeas \idex_if.rd_o[4] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\imm_o~10_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifrd_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.rd_o[4] .is_wysiwyg = "true";
defparam \idex_if.rd_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y27_N25
dffeas \idex_if.jal_o (
	.clk(CPUCLK),
	.d(\jal_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifjal_o),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.jal_o .is_wysiwyg = "true";
defparam \idex_if.jal_o .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N11
dffeas \idex_if.lui_o (
	.clk(CPUCLK),
	.d(\lui_o~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_iflui_o),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.lui_o .is_wysiwyg = "true";
defparam \idex_if.lui_o .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N29
dffeas \idex_if.memToReg_o (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(\dREN_o~0_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\idex_if.rt_o[4]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(idex_ifmemToReg_o),
	.prn(vcc));
// synopsys translate_off
defparam \idex_if.memToReg_o .is_wysiwyg = "true";
defparam \idex_if.memToReg_o .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N4
cycloneive_lcell_comb \aluop_o~0 (
// Equation(s):
// \aluop_o~0_combout  = (ifid_ifinstr_o_26 & (ifid_ifinstr_o_31 & (!ifid_ifinstr_o_28 & ifid_ifinstr_o_27)))

	.dataa(ifid_ifinstr_o_26),
	.datab(ifid_ifinstr_o_31),
	.datac(ifid_ifinstr_o_28),
	.datad(ifid_ifinstr_o_27),
	.cin(gnd),
	.combout(\aluop_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~0 .lut_mask = 16'h0800;
defparam \aluop_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N24
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// \always0~0_combout  = (huiffreeze) # ((always13 & huifflush))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(gnd),
	.datad(huifflush),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'hEECC;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N18
cycloneive_lcell_comb \aluop_o~2 (
// Equation(s):
// \aluop_o~2_combout  = (!ifid_ifinstr_o_26 & ((ifid_ifinstr_o_3 & (!ifid_ifinstr_o_2 & ifid_ifinstr_o_1)) # (!ifid_ifinstr_o_3 & ((ifid_ifinstr_o_1) # (!ifid_ifinstr_o_2)))))

	.dataa(ifid_ifinstr_o_3),
	.datab(ifid_ifinstr_o_26),
	.datac(ifid_ifinstr_o_2),
	.datad(ifid_ifinstr_o_1),
	.cin(gnd),
	.combout(\aluop_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~2 .lut_mask = 16'h1301;
defparam \aluop_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N0
cycloneive_lcell_comb \aluop_o~3 (
// Equation(s):
// \aluop_o~3_combout  = (ifid_ifinstr_o_28 & (((!ifid_ifinstr_o_29)) # (!ifid_ifinstr_o_26))) # (!ifid_ifinstr_o_28 & (((\aluop_o~2_combout ) # (ifid_ifinstr_o_29))))

	.dataa(ifid_ifinstr_o_26),
	.datab(\aluop_o~2_combout ),
	.datac(ifid_ifinstr_o_28),
	.datad(ifid_ifinstr_o_29),
	.cin(gnd),
	.combout(\aluop_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~3 .lut_mask = 16'h5FFC;
defparam \aluop_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N22
cycloneive_lcell_comb \aluop_o~4 (
// Equation(s):
// \aluop_o~4_combout  = (\aluop_o~1_combout  & (!ifid_ifinstr_o_31 & \aluop_o~3_combout ))

	.dataa(\aluop_o~1_combout ),
	.datab(ifid_ifinstr_o_31),
	.datac(gnd),
	.datad(\aluop_o~3_combout ),
	.cin(gnd),
	.combout(\aluop_o~4_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~4 .lut_mask = 16'h2200;
defparam \aluop_o~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N16
cycloneive_lcell_comb \aluop_o~5 (
// Equation(s):
// \aluop_o~5_combout  = (!ifid_ifinstr_o_30 & (!\always0~0_combout  & ((\aluop_o~0_combout ) # (\aluop_o~4_combout ))))

	.dataa(ifid_ifinstr_o_30),
	.datab(\aluop_o~0_combout ),
	.datac(\always0~0_combout ),
	.datad(\aluop_o~4_combout ),
	.cin(gnd),
	.combout(\aluop_o~5_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~5 .lut_mask = 16'h0504;
defparam \aluop_o~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N28
cycloneive_lcell_comb \idex_if.rt_o[4]~0 (
// Equation(s):
// \idex_if.rt_o[4]~0_combout  = (huiffreeze) # (always13)

	.dataa(gnd),
	.datab(huiffreeze),
	.datac(gnd),
	.datad(always1),
	.cin(gnd),
	.combout(\idex_if.rt_o[4]~0_combout ),
	.cout());
// synopsys translate_off
defparam \idex_if.rt_o[4]~0 .lut_mask = 16'hFFCC;
defparam \idex_if.rt_o[4]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N10
cycloneive_lcell_comb \imm_26_o~0 (
// Equation(s):
// \imm_26_o~0_combout  = (ifid_ifinstr_o_16 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(ifid_ifinstr_o_16),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\imm_26_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \imm_26_o~0 .lut_mask = 16'h040C;
defparam \imm_26_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N20
cycloneive_lcell_comb \imm_26_o~1 (
// Equation(s):
// \imm_26_o~1_combout  = (!huiffreeze & (ifid_ifinstr_o_17 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(huifflush),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\imm_26_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \imm_26_o~1 .lut_mask = 16'h1500;
defparam \imm_26_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N16
cycloneive_lcell_comb \imm_26_o~2 (
// Equation(s):
// \imm_26_o~2_combout  = (ifid_ifinstr_o_18 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(ifid_ifinstr_o_18),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\imm_26_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \imm_26_o~2 .lut_mask = 16'h040C;
defparam \imm_26_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N6
cycloneive_lcell_comb \imm_26_o~3 (
// Equation(s):
// \imm_26_o~3_combout  = (!huiffreeze & (ifid_ifinstr_o_19 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(huifflush),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\imm_26_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \imm_26_o~3 .lut_mask = 16'h1500;
defparam \imm_26_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N30
cycloneive_lcell_comb \imm_26_o~4 (
// Equation(s):
// \imm_26_o~4_combout  = (ifid_ifinstr_o_20 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(ifid_ifinstr_o_20),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\imm_26_o~4_combout ),
	.cout());
// synopsys translate_off
defparam \imm_26_o~4 .lut_mask = 16'h040C;
defparam \imm_26_o~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N18
cycloneive_lcell_comb \idex_if.rt_o[4]~feeder (
// Equation(s):
// \idex_if.rt_o[4]~feeder_combout  = \imm_26_o~4_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\imm_26_o~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\idex_if.rt_o[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \idex_if.rt_o[4]~feeder .lut_mask = 16'hF0F0;
defparam \idex_if.rt_o[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N18
cycloneive_lcell_comb \ALUSel_o~0 (
// Equation(s):
// \ALUSel_o~0_combout  = (cuifregWEN & (((!ifid_ifinstr_o_26 & ifid_ifinstr_o_28)) # (!ifid_ifinstr_o_27)))

	.dataa(ifid_ifinstr_o_26),
	.datab(ifid_ifinstr_o_27),
	.datac(ifid_ifinstr_o_28),
	.datad(cuifregWEN),
	.cin(gnd),
	.combout(\ALUSel_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSel_o~0 .lut_mask = 16'h7300;
defparam \ALUSel_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N10
cycloneive_lcell_comb \ALUSel_o~1 (
// Equation(s):
// \ALUSel_o~1_combout  = (!ifid_ifinstr_o_30 & (!\always0~0_combout  & ((\aluop_o~0_combout ) # (\ALUSel_o~0_combout ))))

	.dataa(ifid_ifinstr_o_30),
	.datab(\aluop_o~0_combout ),
	.datac(\always0~0_combout ),
	.datad(\ALUSel_o~0_combout ),
	.cin(gnd),
	.combout(\ALUSel_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSel_o~1 .lut_mask = 16'h0504;
defparam \ALUSel_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N6
cycloneive_lcell_comb \ALUSel_o~3 (
// Equation(s):
// \ALUSel_o~3_combout  = (ifid_ifinstr_o_29 & ((ifid_ifinstr_o_27 & ((!ifid_ifinstr_o_28) # (!ifid_ifinstr_o_26))) # (!ifid_ifinstr_o_27 & ((ifid_ifinstr_o_28)))))

	.dataa(ifid_ifinstr_o_26),
	.datab(ifid_ifinstr_o_27),
	.datac(ifid_ifinstr_o_28),
	.datad(ifid_ifinstr_o_29),
	.cin(gnd),
	.combout(\ALUSel_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSel_o~3 .lut_mask = 16'h7C00;
defparam \ALUSel_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N2
cycloneive_lcell_comb \ALUSel_o~2 (
// Equation(s):
// \ALUSel_o~2_combout  = (!ifid_ifinstr_o_3 & (Equal3 & Equal2))

	.dataa(ifid_ifinstr_o_3),
	.datab(Equal3),
	.datac(Equal2),
	.datad(gnd),
	.cin(gnd),
	.combout(\ALUSel_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSel_o~2 .lut_mask = 16'h4040;
defparam \ALUSel_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N16
cycloneive_lcell_comb \ALUSel_o~4 (
// Equation(s):
// \ALUSel_o~4_combout  = (Equal0 & (!\always0~0_combout  & ((\ALUSel_o~3_combout ) # (\ALUSel_o~2_combout ))))

	.dataa(Equal0),
	.datab(\ALUSel_o~3_combout ),
	.datac(\ALUSel_o~2_combout ),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\ALUSel_o~4_combout ),
	.cout());
// synopsys translate_off
defparam \ALUSel_o~4 .lut_mask = 16'h00A8;
defparam \ALUSel_o~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N8
cycloneive_lcell_comb \imm_o~0 (
// Equation(s):
// \imm_o~0_combout  = (!huiffreeze & (ifid_ifinstr_o_1 & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(ifid_ifinstr_o_1),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\imm_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~0 .lut_mask = 16'h0444;
defparam \imm_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N22
cycloneive_lcell_comb \imm_o~1 (
// Equation(s):
// \imm_o~1_combout  = (!huiffreeze & (ifid_ifinstr_o_7 & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(ifid_ifinstr_o_7),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\imm_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~1 .lut_mask = 16'h0444;
defparam \imm_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N28
cycloneive_lcell_comb \rdat2_o~0 (
// Equation(s):
// \rdat2_o~0_combout  = (ifid_ifinstr_o_20 & (Mux62)) # (!ifid_ifinstr_o_20 & ((Mux621)))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_20),
	.datac(Mux62),
	.datad(Mux621),
	.cin(gnd),
	.combout(\rdat2_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~0 .lut_mask = 16'hF3C0;
defparam \rdat2_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N24
cycloneive_lcell_comb \rdat2_o~1 (
// Equation(s):
// \rdat2_o~1_combout  = (!huiffreeze & (\rdat2_o~0_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat2_o~0_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~1 .lut_mask = 16'h1030;
defparam \rdat2_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N18
cycloneive_lcell_comb \rdat1_o~0 (
// Equation(s):
// \rdat1_o~0_combout  = (ifid_ifinstr_o_25 & ((Mux30))) # (!ifid_ifinstr_o_25 & (Mux301))

	.dataa(ifid_ifinstr_o_25),
	.datab(Mux301),
	.datac(gnd),
	.datad(Mux30),
	.cin(gnd),
	.combout(\rdat1_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~0 .lut_mask = 16'hEE44;
defparam \rdat1_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N4
cycloneive_lcell_comb \rdat1_o~1 (
// Equation(s):
// \rdat1_o~1_combout  = (!huiffreeze & (\rdat1_o~0_combout  & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(\rdat1_o~0_combout ),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\rdat1_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~1 .lut_mask = 16'h0444;
defparam \rdat1_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N2
cycloneive_lcell_comb \imm_26_o~5 (
// Equation(s):
// \imm_26_o~5_combout  = (ifid_ifinstr_o_22 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(ifid_ifinstr_o_22),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\imm_26_o~5_combout ),
	.cout());
// synopsys translate_off
defparam \imm_26_o~5 .lut_mask = 16'h040C;
defparam \imm_26_o~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N4
cycloneive_lcell_comb \idex_if.rs_o[1]~feeder (
// Equation(s):
// \idex_if.rs_o[1]~feeder_combout  = \imm_26_o~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\imm_26_o~5_combout ),
	.cin(gnd),
	.combout(\idex_if.rs_o[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \idex_if.rs_o[1]~feeder .lut_mask = 16'hFF00;
defparam \idex_if.rs_o[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N30
cycloneive_lcell_comb \imm_26_o~6 (
// Equation(s):
// \imm_26_o~6_combout  = (!huiffreeze & (ifid_ifinstr_o_21 & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(ifid_ifinstr_o_21),
	.datad(huifflush),
	.cin(gnd),
	.combout(\imm_26_o~6_combout ),
	.cout());
// synopsys translate_off
defparam \imm_26_o~6 .lut_mask = 16'h1030;
defparam \imm_26_o~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N26
cycloneive_lcell_comb \imm_26_o~7 (
// Equation(s):
// \imm_26_o~7_combout  = (ifid_ifinstr_o_24 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(ifid_ifinstr_o_24),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\imm_26_o~7_combout ),
	.cout());
// synopsys translate_off
defparam \imm_26_o~7 .lut_mask = 16'h040C;
defparam \imm_26_o~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N4
cycloneive_lcell_comb \imm_26_o~8 (
// Equation(s):
// \imm_26_o~8_combout  = (ifid_ifinstr_o_23 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(ifid_ifinstr_o_23),
	.datab(huiffreeze),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\imm_26_o~8_combout ),
	.cout());
// synopsys translate_off
defparam \imm_26_o~8 .lut_mask = 16'h0222;
defparam \imm_26_o~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N20
cycloneive_lcell_comb \idex_if.rs_o[2]~feeder (
// Equation(s):
// \idex_if.rs_o[2]~feeder_combout  = \imm_26_o~8_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\imm_26_o~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\idex_if.rs_o[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \idex_if.rs_o[2]~feeder .lut_mask = 16'hF0F0;
defparam \idex_if.rs_o[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N24
cycloneive_lcell_comb \imm_26_o~9 (
// Equation(s):
// \imm_26_o~9_combout  = (!huiffreeze & (ifid_ifinstr_o_25 & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(ifid_ifinstr_o_25),
	.datad(huifflush),
	.cin(gnd),
	.combout(\imm_26_o~9_combout ),
	.cout());
// synopsys translate_off
defparam \imm_26_o~9 .lut_mask = 16'h1030;
defparam \imm_26_o~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N6
cycloneive_lcell_comb \idex_if.rs_o[4]~feeder (
// Equation(s):
// \idex_if.rs_o[4]~feeder_combout  = \imm_26_o~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\imm_26_o~9_combout ),
	.cin(gnd),
	.combout(\idex_if.rs_o[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \idex_if.rs_o[4]~feeder .lut_mask = 16'hFF00;
defparam \idex_if.rs_o[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N30
cycloneive_lcell_comb \imm_o~2 (
// Equation(s):
// \imm_o~2_combout  = (ifid_ifinstr_o_0 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(ifid_ifinstr_o_0),
	.datab(always1),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\imm_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~2 .lut_mask = 16'h020A;
defparam \imm_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N4
cycloneive_lcell_comb \imm_o~3 (
// Equation(s):
// \imm_o~3_combout  = (!huiffreeze & (ifid_ifinstr_o_6 & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(ifid_ifinstr_o_6),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\imm_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~3 .lut_mask = 16'h0444;
defparam \imm_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N12
cycloneive_lcell_comb \rdat2_o~2 (
// Equation(s):
// \rdat2_o~2_combout  = (ifid_ifinstr_o_20 & (Mux63)) # (!ifid_ifinstr_o_20 & ((Mux631)))

	.dataa(Mux63),
	.datab(ifid_ifinstr_o_20),
	.datac(gnd),
	.datad(Mux631),
	.cin(gnd),
	.combout(\rdat2_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~2 .lut_mask = 16'hBB88;
defparam \rdat2_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N8
cycloneive_lcell_comb \rdat2_o~3 (
// Equation(s):
// \rdat2_o~3_combout  = (!huiffreeze & (\rdat2_o~2_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat2_o~2_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~3 .lut_mask = 16'h1030;
defparam \rdat2_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N12
cycloneive_lcell_comb \rdat1_o~2 (
// Equation(s):
// \rdat1_o~2_combout  = (ifid_ifinstr_o_25 & ((Mux31))) # (!ifid_ifinstr_o_25 & (Mux311))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_25),
	.datac(Mux311),
	.datad(Mux31),
	.cin(gnd),
	.combout(\rdat1_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~2 .lut_mask = 16'hFC30;
defparam \rdat1_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N24
cycloneive_lcell_comb \rdat1_o~3 (
// Equation(s):
// \rdat1_o~3_combout  = (\rdat1_o~2_combout  & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(\rdat1_o~2_combout ),
	.datab(always1),
	.datac(huifflush),
	.datad(huiffreeze),
	.cin(gnd),
	.combout(\rdat1_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~3 .lut_mask = 16'h002A;
defparam \rdat1_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N16
cycloneive_lcell_comb \aluop_o~8 (
// Equation(s):
// \aluop_o~8_combout  = (\aluop_o~7_combout  & (Equal2 & Equal10))

	.dataa(\aluop_o~7_combout ),
	.datab(gnd),
	.datac(Equal2),
	.datad(Equal10),
	.cin(gnd),
	.combout(\aluop_o~8_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~8 .lut_mask = 16'hA000;
defparam \aluop_o~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N16
cycloneive_lcell_comb \aluop_o~6 (
// Equation(s):
// \aluop_o~6_combout  = (ifid_ifinstr_o_28 & (ifid_ifinstr_o_29 & ((!ifid_ifinstr_o_27) # (!ifid_ifinstr_o_26))))

	.dataa(ifid_ifinstr_o_26),
	.datab(ifid_ifinstr_o_27),
	.datac(ifid_ifinstr_o_28),
	.datad(ifid_ifinstr_o_29),
	.cin(gnd),
	.combout(\aluop_o~6_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~6 .lut_mask = 16'h7000;
defparam \aluop_o~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N18
cycloneive_lcell_comb \aluop_o~9 (
// Equation(s):
// \aluop_o~9_combout  = (Equal0 & (!\always0~0_combout  & ((\aluop_o~8_combout ) # (\aluop_o~6_combout ))))

	.dataa(\aluop_o~8_combout ),
	.datab(\aluop_o~6_combout ),
	.datac(Equal0),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\aluop_o~9_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~9 .lut_mask = 16'h00E0;
defparam \aluop_o~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N4
cycloneive_lcell_comb \rdat1_o~4 (
// Equation(s):
// \rdat1_o~4_combout  = (ifid_ifinstr_o_25 & ((Mux29))) # (!ifid_ifinstr_o_25 & (Mux291))

	.dataa(Mux291),
	.datab(ifid_ifinstr_o_25),
	.datac(gnd),
	.datad(Mux29),
	.cin(gnd),
	.combout(\rdat1_o~4_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~4 .lut_mask = 16'hEE22;
defparam \rdat1_o~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N28
cycloneive_lcell_comb \rdat1_o~5 (
// Equation(s):
// \rdat1_o~5_combout  = (!huiffreeze & (\rdat1_o~4_combout  & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(\rdat1_o~4_combout ),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\rdat1_o~5_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~5 .lut_mask = 16'h0444;
defparam \rdat1_o~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N8
cycloneive_lcell_comb \rdat1_o~6 (
// Equation(s):
// \rdat1_o~6_combout  = (ifid_ifinstr_o_25 & ((Mux27))) # (!ifid_ifinstr_o_25 & (Mux271))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_25),
	.datac(Mux271),
	.datad(Mux27),
	.cin(gnd),
	.combout(\rdat1_o~6_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~6 .lut_mask = 16'hFC30;
defparam \rdat1_o~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N14
cycloneive_lcell_comb \rdat1_o~7 (
// Equation(s):
// \rdat1_o~7_combout  = (!huiffreeze & (\rdat1_o~6_combout  & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(\rdat1_o~6_combout ),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\rdat1_o~7_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~7 .lut_mask = 16'h0444;
defparam \rdat1_o~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N2
cycloneive_lcell_comb \rdat1_o~8 (
// Equation(s):
// \rdat1_o~8_combout  = (ifid_ifinstr_o_25 & (Mux28)) # (!ifid_ifinstr_o_25 & ((Mux281)))

	.dataa(ifid_ifinstr_o_25),
	.datab(gnd),
	.datac(Mux28),
	.datad(Mux281),
	.cin(gnd),
	.combout(\rdat1_o~8_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~8 .lut_mask = 16'hF5A0;
defparam \rdat1_o~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N12
cycloneive_lcell_comb \rdat1_o~9 (
// Equation(s):
// \rdat1_o~9_combout  = (!huiffreeze & (\rdat1_o~8_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(huifflush),
	.datad(\rdat1_o~8_combout ),
	.cin(gnd),
	.combout(\rdat1_o~9_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~9 .lut_mask = 16'h1500;
defparam \rdat1_o~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N16
cycloneive_lcell_comb \imm_o~4 (
// Equation(s):
// \imm_o~4_combout  = (!huiffreeze & (ifid_ifinstr_o_2 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(ifid_ifinstr_o_2),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\imm_o~4_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~4 .lut_mask = 16'h0444;
defparam \imm_o~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N6
cycloneive_lcell_comb \idex_if.imm_o[2]~feeder (
// Equation(s):
// \idex_if.imm_o[2]~feeder_combout  = \imm_o~4_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\imm_o~4_combout ),
	.cin(gnd),
	.combout(\idex_if.imm_o[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \idex_if.imm_o[2]~feeder .lut_mask = 16'hFF00;
defparam \idex_if.imm_o[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N22
cycloneive_lcell_comb \imm_o~5 (
// Equation(s):
// \imm_o~5_combout  = (!huiffreeze & (ifid_ifinstr_o_8 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(ifid_ifinstr_o_8),
	.datad(huifflush),
	.cin(gnd),
	.combout(\imm_o~5_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~5 .lut_mask = 16'h1050;
defparam \imm_o~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N24
cycloneive_lcell_comb \idex_if.shamt_o[2]~feeder (
// Equation(s):
// \idex_if.shamt_o[2]~feeder_combout  = \imm_o~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\imm_o~5_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\idex_if.shamt_o[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \idex_if.shamt_o[2]~feeder .lut_mask = 16'hF0F0;
defparam \idex_if.shamt_o[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N14
cycloneive_lcell_comb \rdat2_o~4 (
// Equation(s):
// \rdat2_o~4_combout  = (ifid_ifinstr_o_20 & (Mux61)) # (!ifid_ifinstr_o_20 & ((Mux611)))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_20),
	.datac(Mux61),
	.datad(Mux611),
	.cin(gnd),
	.combout(\rdat2_o~4_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~4 .lut_mask = 16'hF3C0;
defparam \rdat2_o~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N0
cycloneive_lcell_comb \rdat2_o~5 (
// Equation(s):
// \rdat2_o~5_combout  = (\rdat2_o~4_combout  & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(\rdat2_o~4_combout ),
	.datac(huifflush),
	.datad(huiffreeze),
	.cin(gnd),
	.combout(\rdat2_o~5_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~5 .lut_mask = 16'h004C;
defparam \rdat2_o~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N30
cycloneive_lcell_comb \rdat1_o~10 (
// Equation(s):
// \rdat1_o~10_combout  = (ifid_ifinstr_o_25 & (Mux23)) # (!ifid_ifinstr_o_25 & ((Mux231)))

	.dataa(ifid_ifinstr_o_25),
	.datab(gnd),
	.datac(Mux23),
	.datad(Mux231),
	.cin(gnd),
	.combout(\rdat1_o~10_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~10 .lut_mask = 16'hF5A0;
defparam \rdat1_o~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N0
cycloneive_lcell_comb \rdat1_o~11 (
// Equation(s):
// \rdat1_o~11_combout  = (!huiffreeze & (\rdat1_o~10_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(\rdat1_o~10_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~11_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~11 .lut_mask = 16'h1050;
defparam \rdat1_o~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N26
cycloneive_lcell_comb \rdat1_o~12 (
// Equation(s):
// \rdat1_o~12_combout  = (ifid_ifinstr_o_25 & ((Mux24))) # (!ifid_ifinstr_o_25 & (Mux241))

	.dataa(ifid_ifinstr_o_25),
	.datab(gnd),
	.datac(Mux241),
	.datad(Mux24),
	.cin(gnd),
	.combout(\rdat1_o~12_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~12 .lut_mask = 16'hFA50;
defparam \rdat1_o~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N2
cycloneive_lcell_comb \rdat1_o~13 (
// Equation(s):
// \rdat1_o~13_combout  = (!huiffreeze & (\rdat1_o~12_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(\rdat1_o~12_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~13_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~13 .lut_mask = 16'h1050;
defparam \rdat1_o~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N14
cycloneive_lcell_comb \rdat1_o~14 (
// Equation(s):
// \rdat1_o~14_combout  = (ifid_ifinstr_o_25 & ((Mux25))) # (!ifid_ifinstr_o_25 & (Mux251))

	.dataa(ifid_ifinstr_o_25),
	.datab(gnd),
	.datac(Mux251),
	.datad(Mux25),
	.cin(gnd),
	.combout(\rdat1_o~14_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~14 .lut_mask = 16'hFA50;
defparam \rdat1_o~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N20
cycloneive_lcell_comb \rdat1_o~15 (
// Equation(s):
// \rdat1_o~15_combout  = (!huiffreeze & (\rdat1_o~14_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(\rdat1_o~14_combout ),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~15_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~15 .lut_mask = 16'h0444;
defparam \rdat1_o~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N12
cycloneive_lcell_comb \rdat1_o~16 (
// Equation(s):
// \rdat1_o~16_combout  = (ifid_ifinstr_o_25 & ((Mux26))) # (!ifid_ifinstr_o_25 & (Mux261))

	.dataa(ifid_ifinstr_o_25),
	.datab(gnd),
	.datac(Mux261),
	.datad(Mux26),
	.cin(gnd),
	.combout(\rdat1_o~16_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~16 .lut_mask = 16'hFA50;
defparam \rdat1_o~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N6
cycloneive_lcell_comb \rdat1_o~17 (
// Equation(s):
// \rdat1_o~17_combout  = (\rdat1_o~16_combout  & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(\rdat1_o~16_combout ),
	.datab(always1),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~17_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~17 .lut_mask = 16'h020A;
defparam \rdat1_o~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N22
cycloneive_lcell_comb \rdat2_o~6 (
// Equation(s):
// \rdat2_o~6_combout  = (ifid_ifinstr_o_20 & ((Mux60))) # (!ifid_ifinstr_o_20 & (Mux601))

	.dataa(ifid_ifinstr_o_20),
	.datab(Mux601),
	.datac(Mux60),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdat2_o~6_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~6 .lut_mask = 16'hE4E4;
defparam \rdat2_o~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N6
cycloneive_lcell_comb \rdat2_o~7 (
// Equation(s):
// \rdat2_o~7_combout  = (!huiffreeze & (\rdat2_o~6_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(\rdat2_o~6_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~7_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~7 .lut_mask = 16'h1050;
defparam \rdat2_o~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N26
cycloneive_lcell_comb \imm_o~6 (
// Equation(s):
// \imm_o~6_combout  = (!huiffreeze & (ifid_ifinstr_o_3 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(huifflush),
	.datad(ifid_ifinstr_o_3),
	.cin(gnd),
	.combout(\imm_o~6_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~6 .lut_mask = 16'h1500;
defparam \imm_o~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N26
cycloneive_lcell_comb \imm_o~7 (
// Equation(s):
// \imm_o~7_combout  = (!huiffreeze & (ifid_ifinstr_o_9 & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(ifid_ifinstr_o_9),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\imm_o~7_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~7 .lut_mask = 16'h0444;
defparam \imm_o~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N8
cycloneive_lcell_comb \rdat1_o~18 (
// Equation(s):
// \rdat1_o~18_combout  = (ifid_ifinstr_o_25 & ((Mux15))) # (!ifid_ifinstr_o_25 & (Mux151))

	.dataa(ifid_ifinstr_o_25),
	.datab(gnd),
	.datac(Mux151),
	.datad(Mux15),
	.cin(gnd),
	.combout(\rdat1_o~18_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~18 .lut_mask = 16'hFA50;
defparam \rdat1_o~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N24
cycloneive_lcell_comb \rdat1_o~19 (
// Equation(s):
// \rdat1_o~19_combout  = (\rdat1_o~18_combout  & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(\rdat1_o~18_combout ),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~19_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~19 .lut_mask = 16'h040C;
defparam \rdat1_o~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N28
cycloneive_lcell_comb \rdat1_o~20 (
// Equation(s):
// \rdat1_o~20_combout  = (ifid_ifinstr_o_25 & ((Mux16))) # (!ifid_ifinstr_o_25 & (Mux161))

	.dataa(ifid_ifinstr_o_25),
	.datab(gnd),
	.datac(Mux161),
	.datad(Mux16),
	.cin(gnd),
	.combout(\rdat1_o~20_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~20 .lut_mask = 16'hFA50;
defparam \rdat1_o~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N10
cycloneive_lcell_comb \rdat1_o~21 (
// Equation(s):
// \rdat1_o~21_combout  = (!huiffreeze & (\rdat1_o~20_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat1_o~20_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~21_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~21 .lut_mask = 16'h1030;
defparam \rdat1_o~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N4
cycloneive_lcell_comb \rdat1_o~22 (
// Equation(s):
// \rdat1_o~22_combout  = (ifid_ifinstr_o_25 & (Mux17)) # (!ifid_ifinstr_o_25 & ((Mux171)))

	.dataa(Mux17),
	.datab(gnd),
	.datac(ifid_ifinstr_o_25),
	.datad(Mux171),
	.cin(gnd),
	.combout(\rdat1_o~22_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~22 .lut_mask = 16'hAFA0;
defparam \rdat1_o~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N18
cycloneive_lcell_comb \rdat1_o~23 (
// Equation(s):
// \rdat1_o~23_combout  = (!huiffreeze & (\rdat1_o~22_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat1_o~22_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~23_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~23 .lut_mask = 16'h1030;
defparam \rdat1_o~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N18
cycloneive_lcell_comb \rdat1_o~24 (
// Equation(s):
// \rdat1_o~24_combout  = (ifid_ifinstr_o_25 & ((Mux18))) # (!ifid_ifinstr_o_25 & (Mux181))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_25),
	.datac(Mux181),
	.datad(Mux18),
	.cin(gnd),
	.combout(\rdat1_o~24_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~24 .lut_mask = 16'hFC30;
defparam \rdat1_o~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N6
cycloneive_lcell_comb \rdat1_o~25 (
// Equation(s):
// \rdat1_o~25_combout  = (\rdat1_o~24_combout  & (!huiffreeze & ((!always13) # (!huifflush))))

	.dataa(\rdat1_o~24_combout ),
	.datab(huiffreeze),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\rdat1_o~25_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~25 .lut_mask = 16'h0222;
defparam \rdat1_o~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N4
cycloneive_lcell_comb \rdat1_o~26 (
// Equation(s):
// \rdat1_o~26_combout  = (ifid_ifinstr_o_25 & (Mux19)) # (!ifid_ifinstr_o_25 & ((Mux191)))

	.dataa(ifid_ifinstr_o_25),
	.datab(Mux19),
	.datac(Mux191),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdat1_o~26_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~26 .lut_mask = 16'hD8D8;
defparam \rdat1_o~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N0
cycloneive_lcell_comb \rdat1_o~27 (
// Equation(s):
// \rdat1_o~27_combout  = (\rdat1_o~26_combout  & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(\rdat1_o~26_combout ),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~27_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~27 .lut_mask = 16'h040C;
defparam \rdat1_o~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N2
cycloneive_lcell_comb \rdat1_o~28 (
// Equation(s):
// \rdat1_o~28_combout  = (ifid_ifinstr_o_25 & ((Mux20))) # (!ifid_ifinstr_o_25 & (Mux201))

	.dataa(gnd),
	.datab(Mux201),
	.datac(ifid_ifinstr_o_25),
	.datad(Mux20),
	.cin(gnd),
	.combout(\rdat1_o~28_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~28 .lut_mask = 16'hFC0C;
defparam \rdat1_o~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N30
cycloneive_lcell_comb \rdat1_o~29 (
// Equation(s):
// \rdat1_o~29_combout  = (\rdat1_o~28_combout  & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(\rdat1_o~28_combout ),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~29_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~29 .lut_mask = 16'h040C;
defparam \rdat1_o~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N14
cycloneive_lcell_comb \rdat1_o~30 (
// Equation(s):
// \rdat1_o~30_combout  = (ifid_ifinstr_o_25 & (Mux21)) # (!ifid_ifinstr_o_25 & ((Mux211)))

	.dataa(Mux21),
	.datab(Mux211),
	.datac(gnd),
	.datad(ifid_ifinstr_o_25),
	.cin(gnd),
	.combout(\rdat1_o~30_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~30 .lut_mask = 16'hAACC;
defparam \rdat1_o~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N24
cycloneive_lcell_comb \rdat1_o~31 (
// Equation(s):
// \rdat1_o~31_combout  = (!huiffreeze & (\rdat1_o~30_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat1_o~30_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~31_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~31 .lut_mask = 16'h1030;
defparam \rdat1_o~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N16
cycloneive_lcell_comb \rdat1_o~32 (
// Equation(s):
// \rdat1_o~32_combout  = (ifid_ifinstr_o_25 & ((Mux22))) # (!ifid_ifinstr_o_25 & (Mux221))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_25),
	.datac(Mux221),
	.datad(Mux22),
	.cin(gnd),
	.combout(\rdat1_o~32_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~32 .lut_mask = 16'hFC30;
defparam \rdat1_o~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N24
cycloneive_lcell_comb \rdat1_o~33 (
// Equation(s):
// \rdat1_o~33_combout  = (!huiffreeze & (\rdat1_o~32_combout  & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(\rdat1_o~32_combout ),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\rdat1_o~33_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~33 .lut_mask = 16'h0444;
defparam \rdat1_o~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N28
cycloneive_lcell_comb \rdat2_o~8 (
// Equation(s):
// \rdat2_o~8_combout  = (ifid_ifinstr_o_20 & ((Mux59))) # (!ifid_ifinstr_o_20 & (Mux591))

	.dataa(gnd),
	.datab(Mux591),
	.datac(ifid_ifinstr_o_20),
	.datad(Mux59),
	.cin(gnd),
	.combout(\rdat2_o~8_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~8 .lut_mask = 16'hFC0C;
defparam \rdat2_o~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N12
cycloneive_lcell_comb \rdat2_o~9 (
// Equation(s):
// \rdat2_o~9_combout  = (!huiffreeze & (\rdat2_o~8_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat2_o~8_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~9_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~9 .lut_mask = 16'h1030;
defparam \rdat2_o~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N22
cycloneive_lcell_comb \imm_o~8 (
// Equation(s):
// \imm_o~8_combout  = (!huiffreeze & (ifid_ifinstr_o_4 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(ifid_ifinstr_o_4),
	.datad(huifflush),
	.cin(gnd),
	.combout(\imm_o~8_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~8 .lut_mask = 16'h1050;
defparam \imm_o~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N4
cycloneive_lcell_comb \imm_o~9 (
// Equation(s):
// \imm_o~9_combout  = (ifid_ifinstr_o_10 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(ifid_ifinstr_o_10),
	.datac(huifflush),
	.datad(huiffreeze),
	.cin(gnd),
	.combout(\imm_o~9_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~9 .lut_mask = 16'h004C;
defparam \imm_o~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N8
cycloneive_lcell_comb \rdat1_o~34 (
// Equation(s):
// \rdat1_o~34_combout  = (ifid_ifinstr_o_25 & (Mux0)) # (!ifid_ifinstr_o_25 & ((Mux01)))

	.dataa(ifid_ifinstr_o_25),
	.datab(gnd),
	.datac(Mux0),
	.datad(Mux01),
	.cin(gnd),
	.combout(\rdat1_o~34_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~34 .lut_mask = 16'hF5A0;
defparam \rdat1_o~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N0
cycloneive_lcell_comb \rdat1_o~35 (
// Equation(s):
// \rdat1_o~35_combout  = (!huiffreeze & (\rdat1_o~34_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat1_o~34_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~35_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~35 .lut_mask = 16'h1030;
defparam \rdat1_o~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N4
cycloneive_lcell_comb \rdat1_o~36 (
// Equation(s):
// \rdat1_o~36_combout  = (ifid_ifinstr_o_25 & ((Mux2))) # (!ifid_ifinstr_o_25 & (Mux210))

	.dataa(ifid_ifinstr_o_25),
	.datab(gnd),
	.datac(Mux210),
	.datad(Mux2),
	.cin(gnd),
	.combout(\rdat1_o~36_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~36 .lut_mask = 16'hFA50;
defparam \rdat1_o~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N14
cycloneive_lcell_comb \rdat1_o~37 (
// Equation(s):
// \rdat1_o~37_combout  = (!huiffreeze & (\rdat1_o~36_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat1_o~36_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~37_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~37 .lut_mask = 16'h1030;
defparam \rdat1_o~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N12
cycloneive_lcell_comb \rdat1_o~38 (
// Equation(s):
// \rdat1_o~38_combout  = (ifid_ifinstr_o_25 & ((Mux1))) # (!ifid_ifinstr_o_25 & (Mux11))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_25),
	.datac(Mux11),
	.datad(Mux1),
	.cin(gnd),
	.combout(\rdat1_o~38_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~38 .lut_mask = 16'hFC30;
defparam \rdat1_o~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N8
cycloneive_lcell_comb \rdat1_o~39 (
// Equation(s):
// \rdat1_o~39_combout  = (\rdat1_o~38_combout  & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(\rdat1_o~38_combout ),
	.datab(huiffreeze),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~39_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~39 .lut_mask = 16'h0222;
defparam \rdat1_o~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N26
cycloneive_lcell_comb \rdat1_o~40 (
// Equation(s):
// \rdat1_o~40_combout  = (ifid_ifinstr_o_25 & ((Mux3))) # (!ifid_ifinstr_o_25 & (Mux32))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_25),
	.datac(Mux32),
	.datad(Mux3),
	.cin(gnd),
	.combout(\rdat1_o~40_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~40 .lut_mask = 16'hFC30;
defparam \rdat1_o~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N18
cycloneive_lcell_comb \rdat1_o~41 (
// Equation(s):
// \rdat1_o~41_combout  = (\rdat1_o~40_combout  & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(\rdat1_o~40_combout ),
	.datab(huiffreeze),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~41_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~41 .lut_mask = 16'h0222;
defparam \rdat1_o~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N20
cycloneive_lcell_comb \rdat1_o~42 (
// Equation(s):
// \rdat1_o~42_combout  = (ifid_ifinstr_o_25 & ((Mux5))) # (!ifid_ifinstr_o_25 & (Mux51))

	.dataa(ifid_ifinstr_o_25),
	.datab(gnd),
	.datac(Mux51),
	.datad(Mux5),
	.cin(gnd),
	.combout(\rdat1_o~42_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~42 .lut_mask = 16'hFA50;
defparam \rdat1_o~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N18
cycloneive_lcell_comb \rdat1_o~43 (
// Equation(s):
// \rdat1_o~43_combout  = (!huiffreeze & (\rdat1_o~42_combout  & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(\rdat1_o~42_combout ),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\rdat1_o~43_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~43 .lut_mask = 16'h0444;
defparam \rdat1_o~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N14
cycloneive_lcell_comb \rdat1_o~44 (
// Equation(s):
// \rdat1_o~44_combout  = (ifid_ifinstr_o_25 & (Mux4)) # (!ifid_ifinstr_o_25 & ((Mux41)))

	.dataa(Mux4),
	.datab(ifid_ifinstr_o_25),
	.datac(gnd),
	.datad(Mux41),
	.cin(gnd),
	.combout(\rdat1_o~44_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~44 .lut_mask = 16'hBB88;
defparam \rdat1_o~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N20
cycloneive_lcell_comb \rdat1_o~45 (
// Equation(s):
// \rdat1_o~45_combout  = (!huiffreeze & (\rdat1_o~44_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(\rdat1_o~44_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~45_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~45 .lut_mask = 16'h1050;
defparam \rdat1_o~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N30
cycloneive_lcell_comb \rdat1_o~46 (
// Equation(s):
// \rdat1_o~46_combout  = (ifid_ifinstr_o_25 & ((Mux6))) # (!ifid_ifinstr_o_25 & (Mux64))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_25),
	.datac(Mux64),
	.datad(Mux6),
	.cin(gnd),
	.combout(\rdat1_o~46_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~46 .lut_mask = 16'hFC30;
defparam \rdat1_o~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N28
cycloneive_lcell_comb \rdat1_o~47 (
// Equation(s):
// \rdat1_o~47_combout  = (!huiffreeze & (\rdat1_o~46_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat1_o~46_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~47_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~47 .lut_mask = 16'h1030;
defparam \rdat1_o~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N2
cycloneive_lcell_comb \rdat1_o~48 (
// Equation(s):
// \rdat1_o~48_combout  = (ifid_ifinstr_o_25 & ((Mux7))) # (!ifid_ifinstr_o_25 & (Mux71))

	.dataa(Mux71),
	.datab(gnd),
	.datac(ifid_ifinstr_o_25),
	.datad(Mux7),
	.cin(gnd),
	.combout(\rdat1_o~48_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~48 .lut_mask = 16'hFA0A;
defparam \rdat1_o~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N0
cycloneive_lcell_comb \rdat1_o~49 (
// Equation(s):
// \rdat1_o~49_combout  = (!huiffreeze & (\rdat1_o~48_combout  & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(\rdat1_o~48_combout ),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\rdat1_o~49_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~49 .lut_mask = 16'h0444;
defparam \rdat1_o~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N14
cycloneive_lcell_comb \rdat1_o~50 (
// Equation(s):
// \rdat1_o~50_combout  = (ifid_ifinstr_o_25 & (Mux9)) # (!ifid_ifinstr_o_25 & ((Mux91)))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_25),
	.datac(Mux9),
	.datad(Mux91),
	.cin(gnd),
	.combout(\rdat1_o~50_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~50 .lut_mask = 16'hF3C0;
defparam \rdat1_o~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N8
cycloneive_lcell_comb \rdat1_o~51 (
// Equation(s):
// \rdat1_o~51_combout  = (!huiffreeze & (\rdat1_o~50_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(\rdat1_o~50_combout ),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~51_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~51 .lut_mask = 16'h0444;
defparam \rdat1_o~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N16
cycloneive_lcell_comb \rdat1_o~52 (
// Equation(s):
// \rdat1_o~52_combout  = (ifid_ifinstr_o_25 & ((Mux8))) # (!ifid_ifinstr_o_25 & (Mux81))

	.dataa(Mux81),
	.datab(ifid_ifinstr_o_25),
	.datac(gnd),
	.datad(Mux8),
	.cin(gnd),
	.combout(\rdat1_o~52_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~52 .lut_mask = 16'hEE22;
defparam \rdat1_o~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N30
cycloneive_lcell_comb \rdat1_o~53 (
// Equation(s):
// \rdat1_o~53_combout  = (!huiffreeze & (\rdat1_o~52_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(\rdat1_o~52_combout ),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~53_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~53 .lut_mask = 16'h0444;
defparam \rdat1_o~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N0
cycloneive_lcell_comb \rdat1_o~54 (
// Equation(s):
// \rdat1_o~54_combout  = (ifid_ifinstr_o_25 & ((Mux10))) # (!ifid_ifinstr_o_25 & (Mux101))

	.dataa(Mux101),
	.datab(ifid_ifinstr_o_25),
	.datac(gnd),
	.datad(Mux10),
	.cin(gnd),
	.combout(\rdat1_o~54_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~54 .lut_mask = 16'hEE22;
defparam \rdat1_o~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N12
cycloneive_lcell_comb \rdat1_o~55 (
// Equation(s):
// \rdat1_o~55_combout  = (!huiffreeze & (\rdat1_o~54_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat1_o~54_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~55_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~55 .lut_mask = 16'h1030;
defparam \rdat1_o~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N30
cycloneive_lcell_comb \rdat1_o~56 (
// Equation(s):
// \rdat1_o~56_combout  = (ifid_ifinstr_o_25 & (Mux111)) # (!ifid_ifinstr_o_25 & ((Mux112)))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_25),
	.datac(Mux111),
	.datad(Mux112),
	.cin(gnd),
	.combout(\rdat1_o~56_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~56 .lut_mask = 16'hF3C0;
defparam \rdat1_o~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N30
cycloneive_lcell_comb \rdat1_o~57 (
// Equation(s):
// \rdat1_o~57_combout  = (!huiffreeze & (\rdat1_o~56_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat1_o~56_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~57_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~57 .lut_mask = 16'h1030;
defparam \rdat1_o~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N2
cycloneive_lcell_comb \rdat1_o~58 (
// Equation(s):
// \rdat1_o~58_combout  = (ifid_ifinstr_o_25 & (Mux13)) # (!ifid_ifinstr_o_25 & ((Mux131)))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_25),
	.datac(Mux13),
	.datad(Mux131),
	.cin(gnd),
	.combout(\rdat1_o~58_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~58 .lut_mask = 16'hF3C0;
defparam \rdat1_o~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N16
cycloneive_lcell_comb \rdat1_o~59 (
// Equation(s):
// \rdat1_o~59_combout  = (!huiffreeze & (\rdat1_o~58_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(\rdat1_o~58_combout ),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~59_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~59 .lut_mask = 16'h0444;
defparam \rdat1_o~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N4
cycloneive_lcell_comb \rdat1_o~60 (
// Equation(s):
// \rdat1_o~60_combout  = (ifid_ifinstr_o_25 & (Mux12)) # (!ifid_ifinstr_o_25 & ((Mux121)))

	.dataa(Mux12),
	.datab(ifid_ifinstr_o_25),
	.datac(gnd),
	.datad(Mux121),
	.cin(gnd),
	.combout(\rdat1_o~60_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~60 .lut_mask = 16'hBB88;
defparam \rdat1_o~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N14
cycloneive_lcell_comb \rdat1_o~61 (
// Equation(s):
// \rdat1_o~61_combout  = (!huiffreeze & (\rdat1_o~60_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(\rdat1_o~60_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat1_o~61_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~61 .lut_mask = 16'h1050;
defparam \rdat1_o~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N4
cycloneive_lcell_comb \rdat1_o~62 (
// Equation(s):
// \rdat1_o~62_combout  = (ifid_ifinstr_o_25 & (Mux14)) # (!ifid_ifinstr_o_25 & ((Mux141)))

	.dataa(Mux14),
	.datab(ifid_ifinstr_o_25),
	.datac(Mux141),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdat1_o~62_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~62 .lut_mask = 16'hB8B8;
defparam \rdat1_o~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N2
cycloneive_lcell_comb \rdat1_o~63 (
// Equation(s):
// \rdat1_o~63_combout  = (!huiffreeze & (\rdat1_o~62_combout  & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(\rdat1_o~62_combout ),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\rdat1_o~63_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_o~63 .lut_mask = 16'h0444;
defparam \rdat1_o~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N26
cycloneive_lcell_comb \imm_o~10 (
// Equation(s):
// \imm_o~10_combout  = (ifid_ifinstr_o_15 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(ifid_ifinstr_o_15),
	.datab(always1),
	.datac(huifflush),
	.datad(huiffreeze),
	.cin(gnd),
	.combout(\imm_o~10_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~10 .lut_mask = 16'h002A;
defparam \imm_o~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N28
cycloneive_lcell_comb \idex_if.imm_o[15]~feeder (
// Equation(s):
// \idex_if.imm_o[15]~feeder_combout  = \imm_o~10_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\imm_o~10_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\idex_if.imm_o[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \idex_if.imm_o[15]~feeder .lut_mask = 16'hF0F0;
defparam \idex_if.imm_o[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N8
cycloneive_lcell_comb \rdat2_o~10 (
// Equation(s):
// \rdat2_o~10_combout  = (ifid_ifinstr_o_20 & ((Mux321))) # (!ifid_ifinstr_o_20 & (Mux322))

	.dataa(ifid_ifinstr_o_20),
	.datab(gnd),
	.datac(Mux322),
	.datad(Mux321),
	.cin(gnd),
	.combout(\rdat2_o~10_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~10 .lut_mask = 16'hFA50;
defparam \rdat2_o~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N28
cycloneive_lcell_comb \rdat2_o~11 (
// Equation(s):
// \rdat2_o~11_combout  = (!huiffreeze & (\rdat2_o~10_combout  & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(\rdat2_o~10_combout ),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\rdat2_o~11_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~11 .lut_mask = 16'h0444;
defparam \rdat2_o~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N16
cycloneive_lcell_comb \rdat2_o~12 (
// Equation(s):
// \rdat2_o~12_combout  = (ifid_ifinstr_o_20 & ((Mux47))) # (!ifid_ifinstr_o_20 & (Mux471))

	.dataa(ifid_ifinstr_o_20),
	.datab(gnd),
	.datac(Mux471),
	.datad(Mux47),
	.cin(gnd),
	.combout(\rdat2_o~12_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~12 .lut_mask = 16'hFA50;
defparam \rdat2_o~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N12
cycloneive_lcell_comb \rdat2_o~13 (
// Equation(s):
// \rdat2_o~13_combout  = (\rdat2_o~12_combout  & (!huiffreeze & ((!always13) # (!huifflush))))

	.dataa(\rdat2_o~12_combout ),
	.datab(huiffreeze),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\rdat2_o~13_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~13 .lut_mask = 16'h0222;
defparam \rdat2_o~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N8
cycloneive_lcell_comb \rdat2_o~14 (
// Equation(s):
// \rdat2_o~14_combout  = (ifid_ifinstr_o_20 & ((Mux46))) # (!ifid_ifinstr_o_20 & (Mux461))

	.dataa(ifid_ifinstr_o_20),
	.datab(gnd),
	.datac(Mux461),
	.datad(Mux46),
	.cin(gnd),
	.combout(\rdat2_o~14_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~14 .lut_mask = 16'hFA50;
defparam \rdat2_o~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N20
cycloneive_lcell_comb \rdat2_o~15 (
// Equation(s):
// \rdat2_o~15_combout  = (!huiffreeze & (\rdat2_o~14_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat2_o~14_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~15_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~15 .lut_mask = 16'h1030;
defparam \rdat2_o~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N22
cycloneive_lcell_comb \rdat2_o~16 (
// Equation(s):
// \rdat2_o~16_combout  = (ifid_ifinstr_o_20 & ((Mux45))) # (!ifid_ifinstr_o_20 & (Mux451))

	.dataa(Mux451),
	.datab(gnd),
	.datac(ifid_ifinstr_o_20),
	.datad(Mux45),
	.cin(gnd),
	.combout(\rdat2_o~16_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~16 .lut_mask = 16'hFA0A;
defparam \rdat2_o~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N24
cycloneive_lcell_comb \rdat2_o~17 (
// Equation(s):
// \rdat2_o~17_combout  = (!huiffreeze & (\rdat2_o~16_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat2_o~16_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~17_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~17 .lut_mask = 16'h1030;
defparam \rdat2_o~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N14
cycloneive_lcell_comb \rdat2_o~18 (
// Equation(s):
// \rdat2_o~18_combout  = (ifid_ifinstr_o_20 & ((Mux44))) # (!ifid_ifinstr_o_20 & (Mux441))

	.dataa(gnd),
	.datab(Mux441),
	.datac(Mux44),
	.datad(ifid_ifinstr_o_20),
	.cin(gnd),
	.combout(\rdat2_o~18_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~18 .lut_mask = 16'hF0CC;
defparam \rdat2_o~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N0
cycloneive_lcell_comb \rdat2_o~19 (
// Equation(s):
// \rdat2_o~19_combout  = (\rdat2_o~18_combout  & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(\rdat2_o~18_combout ),
	.datab(huiffreeze),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~19_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~19 .lut_mask = 16'h0222;
defparam \rdat2_o~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N0
cycloneive_lcell_comb \rdat2_o~20 (
// Equation(s):
// \rdat2_o~20_combout  = (ifid_ifinstr_o_20 & ((Mux43))) # (!ifid_ifinstr_o_20 & (Mux431))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_20),
	.datac(Mux431),
	.datad(Mux43),
	.cin(gnd),
	.combout(\rdat2_o~20_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~20 .lut_mask = 16'hFC30;
defparam \rdat2_o~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N20
cycloneive_lcell_comb \rdat2_o~21 (
// Equation(s):
// \rdat2_o~21_combout  = (\rdat2_o~20_combout  & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(\rdat2_o~20_combout ),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~21_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~21 .lut_mask = 16'h040C;
defparam \rdat2_o~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N14
cycloneive_lcell_comb \rdat2_o~22 (
// Equation(s):
// \rdat2_o~22_combout  = (ifid_ifinstr_o_20 & (Mux42)) # (!ifid_ifinstr_o_20 & ((Mux421)))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_20),
	.datac(Mux42),
	.datad(Mux421),
	.cin(gnd),
	.combout(\rdat2_o~22_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~22 .lut_mask = 16'hF3C0;
defparam \rdat2_o~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N2
cycloneive_lcell_comb \rdat2_o~23 (
// Equation(s):
// \rdat2_o~23_combout  = (!huiffreeze & (\rdat2_o~22_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(huifflush),
	.datad(\rdat2_o~22_combout ),
	.cin(gnd),
	.combout(\rdat2_o~23_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~23 .lut_mask = 16'h1500;
defparam \rdat2_o~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N26
cycloneive_lcell_comb \rdat2_o~24 (
// Equation(s):
// \rdat2_o~24_combout  = (ifid_ifinstr_o_20 & (Mux411)) # (!ifid_ifinstr_o_20 & ((Mux412)))

	.dataa(Mux411),
	.datab(Mux412),
	.datac(ifid_ifinstr_o_20),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdat2_o~24_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~24 .lut_mask = 16'hACAC;
defparam \rdat2_o~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N24
cycloneive_lcell_comb \rdat2_o~25 (
// Equation(s):
// \rdat2_o~25_combout  = (\rdat2_o~24_combout  & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(\rdat2_o~24_combout ),
	.datab(always1),
	.datac(huifflush),
	.datad(huiffreeze),
	.cin(gnd),
	.combout(\rdat2_o~25_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~25 .lut_mask = 16'h002A;
defparam \rdat2_o~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N14
cycloneive_lcell_comb \rdat2_o~26 (
// Equation(s):
// \rdat2_o~26_combout  = (ifid_ifinstr_o_20 & ((Mux40))) # (!ifid_ifinstr_o_20 & (Mux401))

	.dataa(gnd),
	.datab(Mux401),
	.datac(ifid_ifinstr_o_20),
	.datad(Mux40),
	.cin(gnd),
	.combout(\rdat2_o~26_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~26 .lut_mask = 16'hFC0C;
defparam \rdat2_o~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N10
cycloneive_lcell_comb \rdat2_o~27 (
// Equation(s):
// \rdat2_o~27_combout  = (!huiffreeze & (\rdat2_o~26_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat2_o~26_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~27_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~27 .lut_mask = 16'h1030;
defparam \rdat2_o~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N8
cycloneive_lcell_comb \rdat2_o~28 (
// Equation(s):
// \rdat2_o~28_combout  = (ifid_ifinstr_o_20 & (Mux39)) # (!ifid_ifinstr_o_20 & ((Mux391)))

	.dataa(Mux39),
	.datab(gnd),
	.datac(ifid_ifinstr_o_20),
	.datad(Mux391),
	.cin(gnd),
	.combout(\rdat2_o~28_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~28 .lut_mask = 16'hAFA0;
defparam \rdat2_o~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N30
cycloneive_lcell_comb \rdat2_o~29 (
// Equation(s):
// \rdat2_o~29_combout  = (!huiffreeze & (\rdat2_o~28_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat2_o~28_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~29_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~29 .lut_mask = 16'h1030;
defparam \rdat2_o~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N14
cycloneive_lcell_comb \rdat2_o~30 (
// Equation(s):
// \rdat2_o~30_combout  = (ifid_ifinstr_o_20 & (Mux38)) # (!ifid_ifinstr_o_20 & ((Mux381)))

	.dataa(ifid_ifinstr_o_20),
	.datab(gnd),
	.datac(Mux38),
	.datad(Mux381),
	.cin(gnd),
	.combout(\rdat2_o~30_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~30 .lut_mask = 16'hF5A0;
defparam \rdat2_o~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N16
cycloneive_lcell_comb \rdat2_o~31 (
// Equation(s):
// \rdat2_o~31_combout  = (!huiffreeze & (\rdat2_o~30_combout  & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(\rdat2_o~30_combout ),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\rdat2_o~31_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~31 .lut_mask = 16'h0444;
defparam \rdat2_o~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N18
cycloneive_lcell_comb \rdat2_o~32 (
// Equation(s):
// \rdat2_o~32_combout  = (ifid_ifinstr_o_20 & ((Mux37))) # (!ifid_ifinstr_o_20 & (Mux371))

	.dataa(ifid_ifinstr_o_20),
	.datab(gnd),
	.datac(Mux371),
	.datad(Mux37),
	.cin(gnd),
	.combout(\rdat2_o~32_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~32 .lut_mask = 16'hFA50;
defparam \rdat2_o~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N12
cycloneive_lcell_comb \rdat2_o~33 (
// Equation(s):
// \rdat2_o~33_combout  = (!huiffreeze & (\rdat2_o~32_combout  & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(\rdat2_o~32_combout ),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\rdat2_o~33_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~33 .lut_mask = 16'h0444;
defparam \rdat2_o~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N12
cycloneive_lcell_comb \rdat2_o~34 (
// Equation(s):
// \rdat2_o~34_combout  = (ifid_ifinstr_o_20 & ((Mux58))) # (!ifid_ifinstr_o_20 & (Mux581))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_20),
	.datac(Mux581),
	.datad(Mux58),
	.cin(gnd),
	.combout(\rdat2_o~34_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~34 .lut_mask = 16'hFC30;
defparam \rdat2_o~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N0
cycloneive_lcell_comb \rdat2_o~35 (
// Equation(s):
// \rdat2_o~35_combout  = (!huiffreeze & (\rdat2_o~34_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat2_o~34_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~35_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~35 .lut_mask = 16'h1030;
defparam \rdat2_o~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N22
cycloneive_lcell_comb \imm_o~11 (
// Equation(s):
// \imm_o~11_combout  = (ifid_ifinstr_o_5 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(ifid_ifinstr_o_5),
	.datab(huiffreeze),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\imm_o~11_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~11 .lut_mask = 16'h0222;
defparam \imm_o~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N8
cycloneive_lcell_comb \rdat2_o~36 (
// Equation(s):
// \rdat2_o~36_combout  = (ifid_ifinstr_o_20 & ((Mux57))) # (!ifid_ifinstr_o_20 & (Mux571))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_20),
	.datac(Mux571),
	.datad(Mux57),
	.cin(gnd),
	.combout(\rdat2_o~36_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~36 .lut_mask = 16'hFC30;
defparam \rdat2_o~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N14
cycloneive_lcell_comb \rdat2_o~37 (
// Equation(s):
// \rdat2_o~37_combout  = (!huiffreeze & (\rdat2_o~36_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat2_o~36_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~37_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~37 .lut_mask = 16'h1030;
defparam \rdat2_o~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N8
cycloneive_lcell_comb \rdat2_o~38 (
// Equation(s):
// \rdat2_o~38_combout  = (ifid_ifinstr_o_20 & ((Mux56))) # (!ifid_ifinstr_o_20 & (Mux561))

	.dataa(ifid_ifinstr_o_20),
	.datab(gnd),
	.datac(Mux561),
	.datad(Mux56),
	.cin(gnd),
	.combout(\rdat2_o~38_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~38 .lut_mask = 16'hFA50;
defparam \rdat2_o~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N4
cycloneive_lcell_comb \rdat2_o~39 (
// Equation(s):
// \rdat2_o~39_combout  = (!huiffreeze & (\rdat2_o~38_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat2_o~38_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~39_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~39 .lut_mask = 16'h1030;
defparam \rdat2_o~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N26
cycloneive_lcell_comb \rdat2_o~40 (
// Equation(s):
// \rdat2_o~40_combout  = (ifid_ifinstr_o_20 & ((Mux55))) # (!ifid_ifinstr_o_20 & (Mux551))

	.dataa(gnd),
	.datab(Mux551),
	.datac(ifid_ifinstr_o_20),
	.datad(Mux55),
	.cin(gnd),
	.combout(\rdat2_o~40_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~40 .lut_mask = 16'hFC0C;
defparam \rdat2_o~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N2
cycloneive_lcell_comb \rdat2_o~41 (
// Equation(s):
// \rdat2_o~41_combout  = (!huiffreeze & (\rdat2_o~40_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat2_o~40_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~41_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~41 .lut_mask = 16'h1030;
defparam \rdat2_o~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N4
cycloneive_lcell_comb \rdat2_o~42 (
// Equation(s):
// \rdat2_o~42_combout  = (ifid_ifinstr_o_20 & (Mux36)) # (!ifid_ifinstr_o_20 & ((Mux361)))

	.dataa(ifid_ifinstr_o_20),
	.datab(gnd),
	.datac(Mux36),
	.datad(Mux361),
	.cin(gnd),
	.combout(\rdat2_o~42_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~42 .lut_mask = 16'hF5A0;
defparam \rdat2_o~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N22
cycloneive_lcell_comb \rdat2_o~43 (
// Equation(s):
// \rdat2_o~43_combout  = (!huiffreeze & (\rdat2_o~42_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat2_o~42_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~43_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~43 .lut_mask = 16'h1030;
defparam \rdat2_o~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N14
cycloneive_lcell_comb \rdat2_o~44 (
// Equation(s):
// \rdat2_o~44_combout  = (ifid_ifinstr_o_20 & ((Mux35))) # (!ifid_ifinstr_o_20 & (Mux351))

	.dataa(gnd),
	.datab(Mux351),
	.datac(ifid_ifinstr_o_20),
	.datad(Mux35),
	.cin(gnd),
	.combout(\rdat2_o~44_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~44 .lut_mask = 16'hFC0C;
defparam \rdat2_o~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N6
cycloneive_lcell_comb \rdat2_o~45 (
// Equation(s):
// \rdat2_o~45_combout  = (!huiffreeze & (\rdat2_o~44_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat2_o~44_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~45_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~45 .lut_mask = 16'h1030;
defparam \rdat2_o~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N16
cycloneive_lcell_comb \rdat2_o~46 (
// Equation(s):
// \rdat2_o~46_combout  = (ifid_ifinstr_o_20 & ((Mux34))) # (!ifid_ifinstr_o_20 & (Mux341))

	.dataa(Mux341),
	.datab(gnd),
	.datac(ifid_ifinstr_o_20),
	.datad(Mux34),
	.cin(gnd),
	.combout(\rdat2_o~46_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~46 .lut_mask = 16'hFA0A;
defparam \rdat2_o~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N20
cycloneive_lcell_comb \rdat2_o~47 (
// Equation(s):
// \rdat2_o~47_combout  = (!huiffreeze & (\rdat2_o~46_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(\rdat2_o~46_combout ),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~47_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~47 .lut_mask = 16'h0444;
defparam \rdat2_o~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N18
cycloneive_lcell_comb \rdat2_o~48 (
// Equation(s):
// \rdat2_o~48_combout  = (ifid_ifinstr_o_20 & (Mux33)) # (!ifid_ifinstr_o_20 & ((Mux331)))

	.dataa(gnd),
	.datab(ifid_ifinstr_o_20),
	.datac(Mux33),
	.datad(Mux331),
	.cin(gnd),
	.combout(\rdat2_o~48_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~48 .lut_mask = 16'hF3C0;
defparam \rdat2_o~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N22
cycloneive_lcell_comb \rdat2_o~49 (
// Equation(s):
// \rdat2_o~49_combout  = (!huiffreeze & (\rdat2_o~48_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(\rdat2_o~48_combout ),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~49_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~49 .lut_mask = 16'h0444;
defparam \rdat2_o~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N8
cycloneive_lcell_comb \rdat2_o~50 (
// Equation(s):
// \rdat2_o~50_combout  = (ifid_ifinstr_o_20 & ((Mux54))) # (!ifid_ifinstr_o_20 & (Mux541))

	.dataa(Mux541),
	.datab(ifid_ifinstr_o_20),
	.datac(Mux54),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdat2_o~50_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~50 .lut_mask = 16'hE2E2;
defparam \rdat2_o~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N16
cycloneive_lcell_comb \rdat2_o~51 (
// Equation(s):
// \rdat2_o~51_combout  = (!huiffreeze & (\rdat2_o~50_combout  & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(\rdat2_o~50_combout ),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\rdat2_o~51_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~51 .lut_mask = 16'h0444;
defparam \rdat2_o~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N16
cycloneive_lcell_comb \rdat2_o~52 (
// Equation(s):
// \rdat2_o~52_combout  = (ifid_ifinstr_o_20 & (Mux49)) # (!ifid_ifinstr_o_20 & ((Mux491)))

	.dataa(Mux49),
	.datab(ifid_ifinstr_o_20),
	.datac(gnd),
	.datad(Mux491),
	.cin(gnd),
	.combout(\rdat2_o~52_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~52 .lut_mask = 16'hBB88;
defparam \rdat2_o~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N10
cycloneive_lcell_comb \rdat2_o~53 (
// Equation(s):
// \rdat2_o~53_combout  = (\rdat2_o~52_combout  & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(\rdat2_o~52_combout ),
	.datac(huifflush),
	.datad(huiffreeze),
	.cin(gnd),
	.combout(\rdat2_o~53_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~53 .lut_mask = 16'h004C;
defparam \rdat2_o~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N4
cycloneive_lcell_comb \imm_o~12 (
// Equation(s):
// \imm_o~12_combout  = (ifid_ifinstr_o_14 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(ifid_ifinstr_o_14),
	.datac(huifflush),
	.datad(huiffreeze),
	.cin(gnd),
	.combout(\imm_o~12_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~12 .lut_mask = 16'h004C;
defparam \imm_o~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N24
cycloneive_lcell_comb \idex_if.imm_o[14]~feeder (
// Equation(s):
// \idex_if.imm_o[14]~feeder_combout  = \imm_o~12_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\imm_o~12_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\idex_if.imm_o[14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \idex_if.imm_o[14]~feeder .lut_mask = 16'hF0F0;
defparam \idex_if.imm_o[14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N22
cycloneive_lcell_comb \rdat2_o~54 (
// Equation(s):
// \rdat2_o~54_combout  = (ifid_ifinstr_o_20 & ((Mux48))) # (!ifid_ifinstr_o_20 & (Mux481))

	.dataa(ifid_ifinstr_o_20),
	.datab(Mux481),
	.datac(gnd),
	.datad(Mux48),
	.cin(gnd),
	.combout(\rdat2_o~54_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~54 .lut_mask = 16'hEE44;
defparam \rdat2_o~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N26
cycloneive_lcell_comb \rdat2_o~55 (
// Equation(s):
// \rdat2_o~55_combout  = (!huiffreeze & (\rdat2_o~54_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(huifflush),
	.datad(\rdat2_o~54_combout ),
	.cin(gnd),
	.combout(\rdat2_o~55_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~55 .lut_mask = 16'h1500;
defparam \rdat2_o~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N0
cycloneive_lcell_comb \rdat2_o~56 (
// Equation(s):
// \rdat2_o~56_combout  = (ifid_ifinstr_o_20 & ((Mux53))) # (!ifid_ifinstr_o_20 & (Mux531))

	.dataa(ifid_ifinstr_o_20),
	.datab(gnd),
	.datac(Mux531),
	.datad(Mux53),
	.cin(gnd),
	.combout(\rdat2_o~56_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~56 .lut_mask = 16'hFA50;
defparam \rdat2_o~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N12
cycloneive_lcell_comb \rdat2_o~57 (
// Equation(s):
// \rdat2_o~57_combout  = (!huiffreeze & (\rdat2_o~56_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(\rdat2_o~56_combout ),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~57_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~57 .lut_mask = 16'h0444;
defparam \rdat2_o~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N30
cycloneive_lcell_comb \rdat2_o~58 (
// Equation(s):
// \rdat2_o~58_combout  = (ifid_ifinstr_o_20 & ((Mux52))) # (!ifid_ifinstr_o_20 & (Mux521))

	.dataa(ifid_ifinstr_o_20),
	.datab(gnd),
	.datac(Mux521),
	.datad(Mux52),
	.cin(gnd),
	.combout(\rdat2_o~58_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~58 .lut_mask = 16'hFA50;
defparam \rdat2_o~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N0
cycloneive_lcell_comb \rdat2_o~59 (
// Equation(s):
// \rdat2_o~59_combout  = (!huiffreeze & (\rdat2_o~58_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat2_o~58_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~59_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~59 .lut_mask = 16'h1030;
defparam \rdat2_o~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N4
cycloneive_lcell_comb \imm_o~13 (
// Equation(s):
// \imm_o~13_combout  = (!huiffreeze & (ifid_ifinstr_o_11 & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(ifid_ifinstr_o_11),
	.datad(huifflush),
	.cin(gnd),
	.combout(\imm_o~13_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~13 .lut_mask = 16'h1030;
defparam \imm_o~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N14
cycloneive_lcell_comb \idex_if.imm_o[11]~feeder (
// Equation(s):
// \idex_if.imm_o[11]~feeder_combout  = \imm_o~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\imm_o~13_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\idex_if.imm_o[11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \idex_if.imm_o[11]~feeder .lut_mask = 16'hF0F0;
defparam \idex_if.imm_o[11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N4
cycloneive_lcell_comb \rdat2_o~60 (
// Equation(s):
// \rdat2_o~60_combout  = (ifid_ifinstr_o_20 & (Mux511)) # (!ifid_ifinstr_o_20 & ((Mux512)))

	.dataa(ifid_ifinstr_o_20),
	.datab(Mux511),
	.datac(gnd),
	.datad(Mux512),
	.cin(gnd),
	.combout(\rdat2_o~60_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~60 .lut_mask = 16'hDD88;
defparam \rdat2_o~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N22
cycloneive_lcell_comb \rdat2_o~61 (
// Equation(s):
// \rdat2_o~61_combout  = (!huiffreeze & (\rdat2_o~60_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat2_o~60_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~61_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~61 .lut_mask = 16'h1030;
defparam \rdat2_o~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N30
cycloneive_lcell_comb \imm_o~14 (
// Equation(s):
// \imm_o~14_combout  = (ifid_ifinstr_o_12 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(ifid_ifinstr_o_12),
	.datab(always1),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\imm_o~14_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~14 .lut_mask = 16'h020A;
defparam \imm_o~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N26
cycloneive_lcell_comb \rdat2_o~62 (
// Equation(s):
// \rdat2_o~62_combout  = (ifid_ifinstr_o_20 & ((Mux50))) # (!ifid_ifinstr_o_20 & (Mux501))

	.dataa(Mux501),
	.datab(gnd),
	.datac(ifid_ifinstr_o_20),
	.datad(Mux50),
	.cin(gnd),
	.combout(\rdat2_o~62_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~62 .lut_mask = 16'hFA0A;
defparam \rdat2_o~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N24
cycloneive_lcell_comb \rdat2_o~63 (
// Equation(s):
// \rdat2_o~63_combout  = (!huiffreeze & (\rdat2_o~62_combout  & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(\rdat2_o~62_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\rdat2_o~63_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_o~63 .lut_mask = 16'h1030;
defparam \rdat2_o~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N8
cycloneive_lcell_comb \imm_o~15 (
// Equation(s):
// \imm_o~15_combout  = (ifid_ifinstr_o_13 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(ifid_ifinstr_o_13),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\imm_o~15_combout ),
	.cout());
// synopsys translate_off
defparam \imm_o~15 .lut_mask = 16'h040C;
defparam \imm_o~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N28
cycloneive_lcell_comb \aluop_o~12 (
// Equation(s):
// \aluop_o~12_combout  = (\aluop_o~11_combout  & (!ifid_ifinstr_o_4 & (!ifid_ifinstr_o_26 & !ifid_ifinstr_o_29)))

	.dataa(\aluop_o~11_combout ),
	.datab(ifid_ifinstr_o_4),
	.datac(ifid_ifinstr_o_26),
	.datad(ifid_ifinstr_o_29),
	.cin(gnd),
	.combout(\aluop_o~12_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~12 .lut_mask = 16'h0002;
defparam \aluop_o~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N2
cycloneive_lcell_comb \aluop_o~13 (
// Equation(s):
// \aluop_o~13_combout  = (\aluop_o~12_combout ) # ((ifid_ifinstr_o_28 & ((ifid_ifinstr_o_26) # (!ifid_ifinstr_o_29))))

	.dataa(ifid_ifinstr_o_26),
	.datab(\aluop_o~12_combout ),
	.datac(ifid_ifinstr_o_28),
	.datad(ifid_ifinstr_o_29),
	.cin(gnd),
	.combout(\aluop_o~13_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~13 .lut_mask = 16'hECFC;
defparam \aluop_o~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N18
cycloneive_lcell_comb \aluop_o~14 (
// Equation(s):
// \aluop_o~14_combout  = (Equal0 & (\aluop_o~13_combout  & (!ifid_ifinstr_o_27 & !\always0~0_combout )))

	.dataa(Equal0),
	.datab(\aluop_o~13_combout ),
	.datac(ifid_ifinstr_o_27),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\aluop_o~14_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~14 .lut_mask = 16'h0008;
defparam \aluop_o~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N8
cycloneive_lcell_comb \aluop_o~16 (
// Equation(s):
// \aluop_o~16_combout  = (\aluop_o~15_combout  & (((ifid_ifinstr_o_3 & ifid_ifinstr_o_1)) # (!Equal3)))

	.dataa(\aluop_o~15_combout ),
	.datab(Equal3),
	.datac(ifid_ifinstr_o_3),
	.datad(ifid_ifinstr_o_1),
	.cin(gnd),
	.combout(\aluop_o~16_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~16 .lut_mask = 16'hA222;
defparam \aluop_o~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N22
cycloneive_lcell_comb \aluop_o~17 (
// Equation(s):
// \aluop_o~17_combout  = (Equal14 & (\aluop_o~16_combout  & Equal21))

	.dataa(gnd),
	.datab(Equal14),
	.datac(\aluop_o~16_combout ),
	.datad(Equal21),
	.cin(gnd),
	.combout(\aluop_o~17_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~17 .lut_mask = 16'hC000;
defparam \aluop_o~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y27_N30
cycloneive_lcell_comb \aluop_o~18 (
// Equation(s):
// \aluop_o~18_combout  = (\aluop_o~17_combout ) # ((ifid_ifinstr_o_29 & Equal01))

	.dataa(ifid_ifinstr_o_29),
	.datab(gnd),
	.datac(Equal01),
	.datad(\aluop_o~17_combout ),
	.cin(gnd),
	.combout(\aluop_o~18_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~18 .lut_mask = 16'hFFA0;
defparam \aluop_o~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N14
cycloneive_lcell_comb \aluop_o~19 (
// Equation(s):
// \aluop_o~19_combout  = (!huiffreeze & (\aluop_o~18_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(huifflush),
	.datad(\aluop_o~18_combout ),
	.cin(gnd),
	.combout(\aluop_o~19_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~19 .lut_mask = 16'h1500;
defparam \aluop_o~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N24
cycloneive_lcell_comb \aluop_o~20 (
// Equation(s):
// \aluop_o~20_combout  = (!ifid_ifinstr_o_28 & (ifid_ifinstr_o_27 & ifid_ifinstr_o_31))

	.dataa(ifid_ifinstr_o_28),
	.datab(ifid_ifinstr_o_27),
	.datac(gnd),
	.datad(ifid_ifinstr_o_31),
	.cin(gnd),
	.combout(\aluop_o~20_combout ),
	.cout());
// synopsys translate_off
defparam \aluop_o~20 .lut_mask = 16'h4400;
defparam \aluop_o~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N16
cycloneive_lcell_comb \instr_o~0 (
// Equation(s):
// \instr_o~0_combout  = (!huiffreeze & (ifid_ifinstr_o_26 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(ifid_ifinstr_o_26),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~0 .lut_mask = 16'h0444;
defparam \instr_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N26
cycloneive_lcell_comb \dWEN_o~0 (
// Equation(s):
// \dWEN_o~0_combout  = (ifid_ifinstr_o_29 & (\aluop_o~20_combout  & (!ifid_ifinstr_o_30 & \instr_o~0_combout )))

	.dataa(ifid_ifinstr_o_29),
	.datab(\aluop_o~20_combout ),
	.datac(ifid_ifinstr_o_30),
	.datad(\instr_o~0_combout ),
	.cin(gnd),
	.combout(\dWEN_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \dWEN_o~0 .lut_mask = 16'h0800;
defparam \dWEN_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N8
cycloneive_lcell_comb \dREN_o~0 (
// Equation(s):
// \dREN_o~0_combout  = (!ifid_ifinstr_o_29 & (\aluop_o~20_combout  & (!ifid_ifinstr_o_30 & \instr_o~0_combout )))

	.dataa(ifid_ifinstr_o_29),
	.datab(\aluop_o~20_combout ),
	.datac(ifid_ifinstr_o_30),
	.datad(\instr_o~0_combout ),
	.cin(gnd),
	.combout(\dREN_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \dREN_o~0 .lut_mask = 16'h0400;
defparam \dREN_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N12
cycloneive_lcell_comb \next_pc_o~0 (
// Equation(s):
// \next_pc_o~0_combout  = (ifid_ifnext_pc_o_1 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(ifid_ifnext_pc_o_1),
	.datab(huiffreeze),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~0 .lut_mask = 16'h0222;
defparam \next_pc_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N8
cycloneive_lcell_comb \jumpSel_o~2 (
// Equation(s):
// \jumpSel_o~2_combout  = (Equal21 & (((Equal5 & Equal3)))) # (!Equal21 & (\bne_o~0_combout ))

	.dataa(\bne_o~0_combout ),
	.datab(Equal5),
	.datac(Equal3),
	.datad(Equal21),
	.cin(gnd),
	.combout(\jumpSel_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \jumpSel_o~2 .lut_mask = 16'hC0AA;
defparam \jumpSel_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N16
cycloneive_lcell_comb \jumpSel_o~3 (
// Equation(s):
// \jumpSel_o~3_combout  = (!huiffreeze & (\jumpSel_o~2_combout  & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(\jumpSel_o~2_combout ),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\jumpSel_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \jumpSel_o~3 .lut_mask = 16'h0444;
defparam \jumpSel_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N10
cycloneive_lcell_comb \bne_o~0 (
// Equation(s):
// \bne_o~0_combout  = (Equal0 & (!ifid_ifinstr_o_27 & (ifid_ifinstr_o_28 & !ifid_ifinstr_o_29)))

	.dataa(Equal0),
	.datab(ifid_ifinstr_o_27),
	.datac(ifid_ifinstr_o_28),
	.datad(ifid_ifinstr_o_29),
	.cin(gnd),
	.combout(\bne_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \bne_o~0 .lut_mask = 16'h0020;
defparam \bne_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N30
cycloneive_lcell_comb \jumpSel_o~5 (
// Equation(s):
// \jumpSel_o~5_combout  = (\bne_o~0_combout ) # ((!ifid_ifinstr_o_29 & Equal01))

	.dataa(ifid_ifinstr_o_29),
	.datab(gnd),
	.datac(Equal01),
	.datad(\bne_o~0_combout ),
	.cin(gnd),
	.combout(\jumpSel_o~5_combout ),
	.cout());
// synopsys translate_off
defparam \jumpSel_o~5 .lut_mask = 16'hFF50;
defparam \jumpSel_o~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N26
cycloneive_lcell_comb \jumpSel_o~4 (
// Equation(s):
// \jumpSel_o~4_combout  = (!huiffreeze & (\jumpSel_o~5_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(\jumpSel_o~5_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\jumpSel_o~4_combout ),
	.cout());
// synopsys translate_off
defparam \jumpSel_o~4 .lut_mask = 16'h1050;
defparam \jumpSel_o~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N0
cycloneive_lcell_comb \instr_o~1 (
// Equation(s):
// \instr_o~1_combout  = (ifid_ifinstr_o_31 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(ifid_ifinstr_o_31),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~1 .lut_mask = 16'h040C;
defparam \instr_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N22
cycloneive_lcell_comb \instr_o~2 (
// Equation(s):
// \instr_o~2_combout  = (ifid_ifinstr_o_30 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(ifid_ifinstr_o_30),
	.datab(huiffreeze),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~2 .lut_mask = 16'h0222;
defparam \instr_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N18
cycloneive_lcell_comb \instr_o~3 (
// Equation(s):
// \instr_o~3_combout  = (!huiffreeze & (ifid_ifinstr_o_27 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(ifid_ifinstr_o_27),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~3 .lut_mask = 16'h0444;
defparam \instr_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N14
cycloneive_lcell_comb \instr_o~4 (
// Equation(s):
// \instr_o~4_combout  = (!huiffreeze & (ifid_ifinstr_o_28 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(ifid_ifinstr_o_28),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~4_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~4 .lut_mask = 16'h1050;
defparam \instr_o~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N0
cycloneive_lcell_comb \bne_o~1 (
// Equation(s):
// \bne_o~1_combout  = (\bne_o~0_combout  & \instr_o~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\bne_o~0_combout ),
	.datad(\instr_o~0_combout ),
	.cin(gnd),
	.combout(\bne_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \bne_o~1 .lut_mask = 16'hF000;
defparam \bne_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N18
cycloneive_lcell_comb \PCSel_o~0 (
// Equation(s):
// \PCSel_o~0_combout  = (ifid_ifinstr_o_29 & (((\bne_o~0_combout )))) # (!ifid_ifinstr_o_29 & ((Equal01 & (!ifid_ifinstr_o_26)) # (!Equal01 & ((\bne_o~0_combout )))))

	.dataa(ifid_ifinstr_o_29),
	.datab(ifid_ifinstr_o_26),
	.datac(Equal01),
	.datad(\bne_o~0_combout ),
	.cin(gnd),
	.combout(\PCSel_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \PCSel_o~0 .lut_mask = 16'hBF10;
defparam \PCSel_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N20
cycloneive_lcell_comb \PCSel_o~1 (
// Equation(s):
// \PCSel_o~1_combout  = (!huiffreeze & (\PCSel_o~0_combout  & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(\PCSel_o~0_combout ),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\PCSel_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \PCSel_o~1 .lut_mask = 16'h0444;
defparam \PCSel_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N24
cycloneive_lcell_comb \next_pc_o~1 (
// Equation(s):
// \next_pc_o~1_combout  = (ifid_ifnext_pc_o_0 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(ifid_ifnext_pc_o_0),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~1 .lut_mask = 16'h040C;
defparam \next_pc_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N26
cycloneive_lcell_comb \next_pc_o~2 (
// Equation(s):
// \next_pc_o~2_combout  = (!huiffreeze & (ifid_ifnext_pc_o_3 & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(ifid_ifnext_pc_o_3),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\next_pc_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~2 .lut_mask = 16'h0444;
defparam \next_pc_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N12
cycloneive_lcell_comb \next_pc_o~3 (
// Equation(s):
// \next_pc_o~3_combout  = (ifid_ifnext_pc_o_2 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(ifid_ifnext_pc_o_2),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~3 .lut_mask = 16'h040C;
defparam \next_pc_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N22
cycloneive_lcell_comb \next_pc_o~4 (
// Equation(s):
// \next_pc_o~4_combout  = (ifid_ifnext_pc_o_5 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(ifid_ifnext_pc_o_5),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~4_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~4 .lut_mask = 16'h040C;
defparam \next_pc_o~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N16
cycloneive_lcell_comb \next_pc_o~5 (
// Equation(s):
// \next_pc_o~5_combout  = (!huiffreeze & (ifid_ifnext_pc_o_4 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(huifflush),
	.datad(ifid_ifnext_pc_o_4),
	.cin(gnd),
	.combout(\next_pc_o~5_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~5 .lut_mask = 16'h1500;
defparam \next_pc_o~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N12
cycloneive_lcell_comb \next_pc_o~6 (
// Equation(s):
// \next_pc_o~6_combout  = (!huiffreeze & (ifid_ifnext_pc_o_7 & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(ifid_ifnext_pc_o_7),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\next_pc_o~6_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~6 .lut_mask = 16'h0444;
defparam \next_pc_o~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N2
cycloneive_lcell_comb \next_pc_o~7 (
// Equation(s):
// \next_pc_o~7_combout  = (ifid_ifnext_pc_o_6 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(ifid_ifnext_pc_o_6),
	.datab(huiffreeze),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~7_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~7 .lut_mask = 16'h0222;
defparam \next_pc_o~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N28
cycloneive_lcell_comb \next_pc_o~8 (
// Equation(s):
// \next_pc_o~8_combout  = (!huiffreeze & (ifid_ifnext_pc_o_9 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(ifid_ifnext_pc_o_9),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~8_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~8 .lut_mask = 16'h1050;
defparam \next_pc_o~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N14
cycloneive_lcell_comb \next_pc_o~9 (
// Equation(s):
// \next_pc_o~9_combout  = (ifid_ifnext_pc_o_8 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(ifid_ifnext_pc_o_8),
	.datab(always1),
	.datac(huifflush),
	.datad(huiffreeze),
	.cin(gnd),
	.combout(\next_pc_o~9_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~9 .lut_mask = 16'h002A;
defparam \next_pc_o~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N10
cycloneive_lcell_comb \next_pc_o~10 (
// Equation(s):
// \next_pc_o~10_combout  = (ifid_ifnext_pc_o_11 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(ifid_ifnext_pc_o_11),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~10_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~10 .lut_mask = 16'h040C;
defparam \next_pc_o~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N12
cycloneive_lcell_comb \next_pc_o~11 (
// Equation(s):
// \next_pc_o~11_combout  = (ifid_ifnext_pc_o_10 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(ifid_ifnext_pc_o_10),
	.datab(always1),
	.datac(huifflush),
	.datad(huiffreeze),
	.cin(gnd),
	.combout(\next_pc_o~11_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~11 .lut_mask = 16'h002A;
defparam \next_pc_o~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N28
cycloneive_lcell_comb \next_pc_o~12 (
// Equation(s):
// \next_pc_o~12_combout  = (!huiffreeze & (ifid_ifnext_pc_o_13 & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(ifid_ifnext_pc_o_13),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~12_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~12 .lut_mask = 16'h1030;
defparam \next_pc_o~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N28
cycloneive_lcell_comb \next_pc_o~13 (
// Equation(s):
// \next_pc_o~13_combout  = (!huiffreeze & (ifid_ifnext_pc_o_12 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(ifid_ifnext_pc_o_12),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~13_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~13 .lut_mask = 16'h1050;
defparam \next_pc_o~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N20
cycloneive_lcell_comb \next_pc_o~14 (
// Equation(s):
// \next_pc_o~14_combout  = (!huiffreeze & (ifid_ifnext_pc_o_15 & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(ifid_ifnext_pc_o_15),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~14_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~14 .lut_mask = 16'h1030;
defparam \next_pc_o~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N6
cycloneive_lcell_comb \next_pc_o~15 (
// Equation(s):
// \next_pc_o~15_combout  = (!huiffreeze & (ifid_ifnext_pc_o_14 & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(ifid_ifnext_pc_o_14),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~15_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~15 .lut_mask = 16'h1030;
defparam \next_pc_o~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N30
cycloneive_lcell_comb \next_pc_o~16 (
// Equation(s):
// \next_pc_o~16_combout  = (ifid_ifnext_pc_o_17 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(ifid_ifnext_pc_o_17),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~16_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~16 .lut_mask = 16'h040C;
defparam \next_pc_o~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N16
cycloneive_lcell_comb \next_pc_o~17 (
// Equation(s):
// \next_pc_o~17_combout  = (!huiffreeze & (ifid_ifnext_pc_o_16 & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(ifid_ifnext_pc_o_16),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~17_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~17 .lut_mask = 16'h1030;
defparam \next_pc_o~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N4
cycloneive_lcell_comb \next_pc_o~18 (
// Equation(s):
// \next_pc_o~18_combout  = (ifid_ifnext_pc_o_19 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(ifid_ifnext_pc_o_19),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~18_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~18 .lut_mask = 16'h040C;
defparam \next_pc_o~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N10
cycloneive_lcell_comb \next_pc_o~19 (
// Equation(s):
// \next_pc_o~19_combout  = (!huiffreeze & (ifid_ifnext_pc_o_18 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(ifid_ifnext_pc_o_18),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~19_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~19 .lut_mask = 16'h1050;
defparam \next_pc_o~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N10
cycloneive_lcell_comb \next_pc_o~20 (
// Equation(s):
// \next_pc_o~20_combout  = (ifid_ifnext_pc_o_21 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(ifid_ifnext_pc_o_21),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~20_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~20 .lut_mask = 16'h040C;
defparam \next_pc_o~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N28
cycloneive_lcell_comb \next_pc_o~21 (
// Equation(s):
// \next_pc_o~21_combout  = (!huiffreeze & (ifid_ifnext_pc_o_20 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(ifid_ifnext_pc_o_20),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~21_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~21 .lut_mask = 16'h1050;
defparam \next_pc_o~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N2
cycloneive_lcell_comb \next_pc_o~22 (
// Equation(s):
// \next_pc_o~22_combout  = (!huiffreeze & (ifid_ifnext_pc_o_23 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(ifid_ifnext_pc_o_23),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~22_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~22 .lut_mask = 16'h1050;
defparam \next_pc_o~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N26
cycloneive_lcell_comb \next_pc_o~23 (
// Equation(s):
// \next_pc_o~23_combout  = (ifid_ifnext_pc_o_22 & (!huiffreeze & ((!always13) # (!huifflush))))

	.dataa(ifid_ifnext_pc_o_22),
	.datab(huiffreeze),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\next_pc_o~23_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~23 .lut_mask = 16'h0222;
defparam \next_pc_o~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N0
cycloneive_lcell_comb \next_pc_o~24 (
// Equation(s):
// \next_pc_o~24_combout  = (!huiffreeze & (ifid_ifnext_pc_o_25 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(ifid_ifnext_pc_o_25),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~24_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~24 .lut_mask = 16'h1050;
defparam \next_pc_o~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N28
cycloneive_lcell_comb \next_pc_o~25 (
// Equation(s):
// \next_pc_o~25_combout  = (!huiffreeze & (ifid_ifnext_pc_o_24 & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(huifflush),
	.datad(ifid_ifnext_pc_o_24),
	.cin(gnd),
	.combout(\next_pc_o~25_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~25 .lut_mask = 16'h1300;
defparam \next_pc_o~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N6
cycloneive_lcell_comb \next_pc_o~26 (
// Equation(s):
// \next_pc_o~26_combout  = (!huiffreeze & (ifid_ifnext_pc_o_27 & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(huifflush),
	.datad(ifid_ifnext_pc_o_27),
	.cin(gnd),
	.combout(\next_pc_o~26_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~26 .lut_mask = 16'h1300;
defparam \next_pc_o~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N6
cycloneive_lcell_comb \next_pc_o~27 (
// Equation(s):
// \next_pc_o~27_combout  = (!huiffreeze & (ifid_ifnext_pc_o_26 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(ifid_ifnext_pc_o_26),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~27_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~27 .lut_mask = 16'h1050;
defparam \next_pc_o~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N10
cycloneive_lcell_comb \next_pc_o~28 (
// Equation(s):
// \next_pc_o~28_combout  = (ifid_ifnext_pc_o_29 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(ifid_ifnext_pc_o_29),
	.datab(huiffreeze),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~28_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~28 .lut_mask = 16'h0222;
defparam \next_pc_o~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N22
cycloneive_lcell_comb \next_pc_o~29 (
// Equation(s):
// \next_pc_o~29_combout  = (!huiffreeze & (ifid_ifnext_pc_o_28 & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(huiffreeze),
	.datac(ifid_ifnext_pc_o_28),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~29_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~29 .lut_mask = 16'h1030;
defparam \next_pc_o~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N20
cycloneive_lcell_comb \next_pc_o~30 (
// Equation(s):
// \next_pc_o~30_combout  = (ifid_ifnext_pc_o_31 & (!huiffreeze & ((!huifflush) # (!always13))))

	.dataa(ifid_ifnext_pc_o_31),
	.datab(always1),
	.datac(huiffreeze),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~30_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~30 .lut_mask = 16'h020A;
defparam \next_pc_o~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N26
cycloneive_lcell_comb \next_pc_o~31 (
// Equation(s):
// \next_pc_o~31_combout  = (!huiffreeze & (ifid_ifnext_pc_o_30 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(ifid_ifnext_pc_o_30),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~31_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~31 .lut_mask = 16'h1050;
defparam \next_pc_o~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N2
cycloneive_lcell_comb \lui_o~2 (
// Equation(s):
// \lui_o~2_combout  = (ifid_ifinstr_o_29 & (ifid_ifinstr_o_28 & ifid_ifinstr_o_27))

	.dataa(ifid_ifinstr_o_29),
	.datab(gnd),
	.datac(ifid_ifinstr_o_28),
	.datad(ifid_ifinstr_o_27),
	.cin(gnd),
	.combout(\lui_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \lui_o~2 .lut_mask = 16'hA000;
defparam \lui_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N12
cycloneive_lcell_comb \halt_o~0 (
// Equation(s):
// \halt_o~0_combout  = (ifid_ifinstr_o_31 & (\lui_o~2_combout  & (ifid_ifinstr_o_30 & \instr_o~0_combout )))

	.dataa(ifid_ifinstr_o_31),
	.datab(\lui_o~2_combout ),
	.datac(ifid_ifinstr_o_30),
	.datad(\instr_o~0_combout ),
	.cin(gnd),
	.combout(\halt_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \halt_o~0 .lut_mask = 16'h8000;
defparam \halt_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N16
cycloneive_lcell_comb \RegDest_o~0 (
// Equation(s):
// \RegDest_o~0_combout  = (ifid_ifinstr_o_29) # (!Equal01)

	.dataa(gnd),
	.datab(ifid_ifinstr_o_29),
	.datac(gnd),
	.datad(Equal01),
	.cin(gnd),
	.combout(\RegDest_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \RegDest_o~0 .lut_mask = 16'hCCFF;
defparam \RegDest_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N6
cycloneive_lcell_comb \RegDest_o~1 (
// Equation(s):
// \RegDest_o~1_combout  = (!huiffreeze & (!\RegDest_o~0_combout  & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(\RegDest_o~0_combout ),
	.datad(huifflush),
	.cin(gnd),
	.combout(\RegDest_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \RegDest_o~1 .lut_mask = 16'h0105;
defparam \RegDest_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N16
cycloneive_lcell_comb \idex_if.rd_o[1]~feeder (
// Equation(s):
// \idex_if.rd_o[1]~feeder_combout  = \imm_o~14_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\imm_o~14_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\idex_if.rd_o[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \idex_if.rd_o[1]~feeder .lut_mask = 16'hF0F0;
defparam \idex_if.rd_o[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N28
cycloneive_lcell_comb \RegDest_o~2 (
// Equation(s):
// \RegDest_o~2_combout  = (\RegDest_o~0_combout  & (((\aluop_o~16_combout  & !Equal14)) # (!Equal21)))

	.dataa(\RegDest_o~0_combout ),
	.datab(Equal21),
	.datac(\aluop_o~16_combout ),
	.datad(Equal14),
	.cin(gnd),
	.combout(\RegDest_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \RegDest_o~2 .lut_mask = 16'h22A2;
defparam \RegDest_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N10
cycloneive_lcell_comb \RegDest_o~3 (
// Equation(s):
// \RegDest_o~3_combout  = (!huiffreeze & (\RegDest_o~2_combout  & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(\RegDest_o~2_combout ),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\RegDest_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \RegDest_o~3 .lut_mask = 16'h0444;
defparam \RegDest_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N18
cycloneive_lcell_comb \idex_if.rd_o[2]~feeder (
// Equation(s):
// \idex_if.rd_o[2]~feeder_combout  = \imm_o~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\imm_o~15_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\idex_if.rd_o[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \idex_if.rd_o[2]~feeder .lut_mask = 16'hF0F0;
defparam \idex_if.rd_o[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N10
cycloneive_lcell_comb \regWEN_o~0 (
// Equation(s):
// \regWEN_o~0_combout  = (!huiffreeze & (cuifregWEN1 & ((!huifflush) # (!always13))))

	.dataa(huiffreeze),
	.datab(always1),
	.datac(cuifregWEN1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\regWEN_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \regWEN_o~0 .lut_mask = 16'h1050;
defparam \regWEN_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N24
cycloneive_lcell_comb \jal_o~0 (
// Equation(s):
// \jal_o~0_combout  = (!huiffreeze & (Equal1 & ((!always13) # (!huifflush))))

	.dataa(huiffreeze),
	.datab(Equal1),
	.datac(huifflush),
	.datad(always1),
	.cin(gnd),
	.combout(\jal_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \jal_o~0 .lut_mask = 16'h0444;
defparam \jal_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N10
cycloneive_lcell_comb \lui_o~3 (
// Equation(s):
// \lui_o~3_combout  = (!ifid_ifinstr_o_31 & (\lui_o~2_combout  & (!ifid_ifinstr_o_30 & \instr_o~0_combout )))

	.dataa(ifid_ifinstr_o_31),
	.datab(\lui_o~2_combout ),
	.datac(ifid_ifinstr_o_30),
	.datad(\instr_o~0_combout ),
	.cin(gnd),
	.combout(\lui_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \lui_o~3 .lut_mask = 16'h0400;
defparam \lui_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module if_id (
	nextpc_2,
	nextpc_3,
	nextpc_4,
	nextpc_5,
	nextpc_6,
	nextpc_7,
	nextpc_8,
	nextpc_9,
	nextpc_10,
	nextpc_11,
	nextpc_12,
	nextpc_13,
	nextpc_14,
	nextpc_15,
	nextpc_16,
	nextpc_17,
	nextpc_18,
	nextpc_19,
	nextpc_20,
	nextpc_21,
	nextpc_22,
	nextpc_23,
	nextpc_24,
	nextpc_25,
	nextpc_26,
	nextpc_27,
	nextpc_28,
	nextpc_29,
	nextpc_30,
	nextpc_31,
	ramiframload_0,
	pc_1,
	pc_0,
	ramiframload_1,
	always1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	always11,
	ifid_ifinstr_o_17,
	ifid_ifinstr_o_16,
	ifid_ifinstr_o_19,
	ifid_ifinstr_o_18,
	ifid_ifinstr_o_20,
	ifid_ifinstr_o_22,
	ifid_ifinstr_o_21,
	ifid_ifinstr_o_24,
	ifid_ifinstr_o_23,
	ifid_ifinstr_o_25,
	huiffreeze,
	huifflush,
	ifid_ifinstr_o_26,
	ifid_ifinstr_o_31,
	ifid_ifinstr_o_27,
	ifid_ifinstr_o_28,
	ifid_ifinstr_o_30,
	ifid_ifinstr_o_5,
	ifid_ifinstr_o_4,
	ifid_ifinstr_o_29,
	ifid_ifinstr_o_1,
	ifid_ifinstr_o_3,
	ifid_ifinstr_o_2,
	ifid_ifinstr_o_0,
	ifid_ifinstr_o_7,
	ifid_ifinstr_o_6,
	ifid_ifinstr_o_8,
	ifid_ifinstr_o_9,
	ifid_ifinstr_o_10,
	ifid_ifinstr_o_15,
	ifid_ifinstr_o_14,
	ifid_ifinstr_o_11,
	ifid_ifinstr_o_12,
	ifid_ifinstr_o_13,
	ifid_ifnext_pc_o_1,
	ifid_ifnext_pc_o_0,
	ifid_ifnext_pc_o_3,
	ifid_ifnext_pc_o_2,
	ifid_ifnext_pc_o_5,
	ifid_ifnext_pc_o_4,
	ifid_ifnext_pc_o_7,
	ifid_ifnext_pc_o_6,
	ifid_ifnext_pc_o_9,
	ifid_ifnext_pc_o_8,
	ifid_ifnext_pc_o_11,
	ifid_ifnext_pc_o_10,
	ifid_ifnext_pc_o_13,
	ifid_ifnext_pc_o_12,
	ifid_ifnext_pc_o_15,
	ifid_ifnext_pc_o_14,
	ifid_ifnext_pc_o_17,
	ifid_ifnext_pc_o_16,
	ifid_ifnext_pc_o_19,
	ifid_ifnext_pc_o_18,
	ifid_ifnext_pc_o_21,
	ifid_ifnext_pc_o_20,
	ifid_ifnext_pc_o_23,
	ifid_ifnext_pc_o_22,
	ifid_ifnext_pc_o_25,
	ifid_ifnext_pc_o_24,
	ifid_ifnext_pc_o_27,
	ifid_ifnext_pc_o_26,
	ifid_ifnext_pc_o_29,
	ifid_ifnext_pc_o_28,
	ifid_ifnext_pc_o_31,
	ifid_ifnext_pc_o_30,
	CPUCLK,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	nextpc_2;
input 	nextpc_3;
input 	nextpc_4;
input 	nextpc_5;
input 	nextpc_6;
input 	nextpc_7;
input 	nextpc_8;
input 	nextpc_9;
input 	nextpc_10;
input 	nextpc_11;
input 	nextpc_12;
input 	nextpc_13;
input 	nextpc_14;
input 	nextpc_15;
input 	nextpc_16;
input 	nextpc_17;
input 	nextpc_18;
input 	nextpc_19;
input 	nextpc_20;
input 	nextpc_21;
input 	nextpc_22;
input 	nextpc_23;
input 	nextpc_24;
input 	nextpc_25;
input 	nextpc_26;
input 	nextpc_27;
input 	nextpc_28;
input 	nextpc_29;
input 	nextpc_30;
input 	nextpc_31;
input 	ramiframload_0;
input 	pc_1;
input 	pc_0;
input 	ramiframload_1;
input 	always1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
input 	always11;
output 	ifid_ifinstr_o_17;
output 	ifid_ifinstr_o_16;
output 	ifid_ifinstr_o_19;
output 	ifid_ifinstr_o_18;
output 	ifid_ifinstr_o_20;
output 	ifid_ifinstr_o_22;
output 	ifid_ifinstr_o_21;
output 	ifid_ifinstr_o_24;
output 	ifid_ifinstr_o_23;
output 	ifid_ifinstr_o_25;
input 	huiffreeze;
input 	huifflush;
output 	ifid_ifinstr_o_26;
output 	ifid_ifinstr_o_31;
output 	ifid_ifinstr_o_27;
output 	ifid_ifinstr_o_28;
output 	ifid_ifinstr_o_30;
output 	ifid_ifinstr_o_5;
output 	ifid_ifinstr_o_4;
output 	ifid_ifinstr_o_29;
output 	ifid_ifinstr_o_1;
output 	ifid_ifinstr_o_3;
output 	ifid_ifinstr_o_2;
output 	ifid_ifinstr_o_0;
output 	ifid_ifinstr_o_7;
output 	ifid_ifinstr_o_6;
output 	ifid_ifinstr_o_8;
output 	ifid_ifinstr_o_9;
output 	ifid_ifinstr_o_10;
output 	ifid_ifinstr_o_15;
output 	ifid_ifinstr_o_14;
output 	ifid_ifinstr_o_11;
output 	ifid_ifinstr_o_12;
output 	ifid_ifinstr_o_13;
output 	ifid_ifnext_pc_o_1;
output 	ifid_ifnext_pc_o_0;
output 	ifid_ifnext_pc_o_3;
output 	ifid_ifnext_pc_o_2;
output 	ifid_ifnext_pc_o_5;
output 	ifid_ifnext_pc_o_4;
output 	ifid_ifnext_pc_o_7;
output 	ifid_ifnext_pc_o_6;
output 	ifid_ifnext_pc_o_9;
output 	ifid_ifnext_pc_o_8;
output 	ifid_ifnext_pc_o_11;
output 	ifid_ifnext_pc_o_10;
output 	ifid_ifnext_pc_o_13;
output 	ifid_ifnext_pc_o_12;
output 	ifid_ifnext_pc_o_15;
output 	ifid_ifnext_pc_o_14;
output 	ifid_ifnext_pc_o_17;
output 	ifid_ifnext_pc_o_16;
output 	ifid_ifnext_pc_o_19;
output 	ifid_ifnext_pc_o_18;
output 	ifid_ifnext_pc_o_21;
output 	ifid_ifnext_pc_o_20;
output 	ifid_ifnext_pc_o_23;
output 	ifid_ifnext_pc_o_22;
output 	ifid_ifnext_pc_o_25;
output 	ifid_ifnext_pc_o_24;
output 	ifid_ifnext_pc_o_27;
output 	ifid_ifnext_pc_o_26;
output 	ifid_ifnext_pc_o_29;
output 	ifid_ifnext_pc_o_28;
output 	ifid_ifnext_pc_o_31;
output 	ifid_ifnext_pc_o_30;
input 	CPUCLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \instr_o~0_combout ;
wire \ifid_if.instr_o[25]~0_combout ;
wire \instr_o~1_combout ;
wire \instr_o~2_combout ;
wire \instr_o~3_combout ;
wire \instr_o~4_combout ;
wire \instr_o~5_combout ;
wire \instr_o~6_combout ;
wire \instr_o~7_combout ;
wire \instr_o~8_combout ;
wire \instr_o~9_combout ;
wire \instr_o~10_combout ;
wire \instr_o~11_combout ;
wire \instr_o~12_combout ;
wire \instr_o~13_combout ;
wire \instr_o~14_combout ;
wire \instr_o~15_combout ;
wire \instr_o~16_combout ;
wire \instr_o~17_combout ;
wire \instr_o~18_combout ;
wire \instr_o~19_combout ;
wire \instr_o~20_combout ;
wire \instr_o~21_combout ;
wire \instr_o~22_combout ;
wire \instr_o~23_combout ;
wire \instr_o~24_combout ;
wire \instr_o~25_combout ;
wire \instr_o~26_combout ;
wire \instr_o~27_combout ;
wire \instr_o~28_combout ;
wire \instr_o~29_combout ;
wire \instr_o~30_combout ;
wire \instr_o~31_combout ;
wire \next_pc_o~0_combout ;
wire \next_pc_o~1_combout ;
wire \next_pc_o~2_combout ;
wire \next_pc_o~3_combout ;
wire \next_pc_o~4_combout ;
wire \next_pc_o~5_combout ;
wire \next_pc_o~6_combout ;
wire \next_pc_o~7_combout ;
wire \next_pc_o~8_combout ;
wire \next_pc_o~9_combout ;
wire \next_pc_o~10_combout ;
wire \next_pc_o~11_combout ;
wire \next_pc_o~12_combout ;
wire \next_pc_o~13_combout ;
wire \next_pc_o~14_combout ;
wire \next_pc_o~15_combout ;
wire \next_pc_o~16_combout ;
wire \next_pc_o~17_combout ;
wire \next_pc_o~18_combout ;
wire \next_pc_o~19_combout ;
wire \next_pc_o~20_combout ;
wire \next_pc_o~21_combout ;
wire \next_pc_o~22_combout ;
wire \next_pc_o~23_combout ;
wire \next_pc_o~24_combout ;
wire \next_pc_o~25_combout ;
wire \next_pc_o~26_combout ;
wire \next_pc_o~27_combout ;
wire \next_pc_o~28_combout ;
wire \next_pc_o~29_combout ;
wire \next_pc_o~30_combout ;
wire \next_pc_o~31_combout ;


// Location: FF_X62_Y31_N25
dffeas \ifid_if.instr_o[17] (
	.clk(CPUCLK),
	.d(\instr_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_17),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[17] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N17
dffeas \ifid_if.instr_o[16] (
	.clk(CPUCLK),
	.d(\instr_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_16),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[16] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N7
dffeas \ifid_if.instr_o[19] (
	.clk(CPUCLK),
	.d(\instr_o~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_19),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[19] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y27_N7
dffeas \ifid_if.instr_o[18] (
	.clk(CPUCLK),
	.d(\instr_o~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_18),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[18] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N21
dffeas \ifid_if.instr_o[20] (
	.clk(CPUCLK),
	.d(\instr_o~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_20),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[20] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N23
dffeas \ifid_if.instr_o[22] (
	.clk(CPUCLK),
	.d(\instr_o~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_22),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[22] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N19
dffeas \ifid_if.instr_o[21] (
	.clk(CPUCLK),
	.d(\instr_o~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_21),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[21] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N5
dffeas \ifid_if.instr_o[24] (
	.clk(CPUCLK),
	.d(\instr_o~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_24),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[24] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N11
dffeas \ifid_if.instr_o[23] (
	.clk(CPUCLK),
	.d(\instr_o~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_23),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[23] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N25
dffeas \ifid_if.instr_o[25] (
	.clk(CPUCLK),
	.d(\instr_o~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_25),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[25] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N25
dffeas \ifid_if.instr_o[26] (
	.clk(CPUCLK),
	.d(\instr_o~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_26),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[26] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N1
dffeas \ifid_if.instr_o[31] (
	.clk(CPUCLK),
	.d(\instr_o~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_31),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[31] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N31
dffeas \ifid_if.instr_o[27] (
	.clk(CPUCLK),
	.d(\instr_o~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_27),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[27] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N31
dffeas \ifid_if.instr_o[28] (
	.clk(CPUCLK),
	.d(\instr_o~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_28),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[28] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y27_N3
dffeas \ifid_if.instr_o[30] (
	.clk(CPUCLK),
	.d(\instr_o~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_30),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[30] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y28_N21
dffeas \ifid_if.instr_o[5] (
	.clk(CPUCLK),
	.d(\instr_o~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_5),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[5] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N5
dffeas \ifid_if.instr_o[4] (
	.clk(CPUCLK),
	.d(\instr_o~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[4] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N19
dffeas \ifid_if.instr_o[29] (
	.clk(CPUCLK),
	.d(\instr_o~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_29),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[29] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N13
dffeas \ifid_if.instr_o[1] (
	.clk(CPUCLK),
	.d(\instr_o~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[1] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y27_N5
dffeas \ifid_if.instr_o[3] (
	.clk(CPUCLK),
	.d(\instr_o~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[3] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N19
dffeas \ifid_if.instr_o[2] (
	.clk(CPUCLK),
	.d(\instr_o~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[2] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N17
dffeas \ifid_if.instr_o[0] (
	.clk(CPUCLK),
	.d(\instr_o~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[0] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N19
dffeas \ifid_if.instr_o[7] (
	.clk(CPUCLK),
	.d(\instr_o~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_7),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[7] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N25
dffeas \ifid_if.instr_o[6] (
	.clk(CPUCLK),
	.d(\instr_o~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_6),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[6] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N5
dffeas \ifid_if.instr_o[8] (
	.clk(CPUCLK),
	.d(\instr_o~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_8),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[8] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N31
dffeas \ifid_if.instr_o[9] (
	.clk(CPUCLK),
	.d(\instr_o~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_9),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[9] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N15
dffeas \ifid_if.instr_o[10] (
	.clk(CPUCLK),
	.d(\instr_o~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_10),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[10] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N13
dffeas \ifid_if.instr_o[15] (
	.clk(CPUCLK),
	.d(\instr_o~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_15),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[15] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N21
dffeas \ifid_if.instr_o[14] (
	.clk(CPUCLK),
	.d(\instr_o~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_14),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[14] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N15
dffeas \ifid_if.instr_o[11] (
	.clk(CPUCLK),
	.d(\instr_o~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_11),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[11] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N5
dffeas \ifid_if.instr_o[12] (
	.clk(CPUCLK),
	.d(\instr_o~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_12),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[12] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N9
dffeas \ifid_if.instr_o[13] (
	.clk(CPUCLK),
	.d(\instr_o~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifinstr_o_13),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.instr_o[13] .is_wysiwyg = "true";
defparam \ifid_if.instr_o[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y29_N31
dffeas \ifid_if.next_pc_o[1] (
	.clk(CPUCLK),
	.d(\next_pc_o~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[1] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y29_N1
dffeas \ifid_if.next_pc_o[0] (
	.clk(CPUCLK),
	.d(\next_pc_o~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[0] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N9
dffeas \ifid_if.next_pc_o[3] (
	.clk(CPUCLK),
	.d(\next_pc_o~2_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[3] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N7
dffeas \ifid_if.next_pc_o[2] (
	.clk(CPUCLK),
	.d(\next_pc_o~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[2] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N23
dffeas \ifid_if.next_pc_o[5] (
	.clk(CPUCLK),
	.d(\next_pc_o~4_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_5),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[5] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N23
dffeas \ifid_if.next_pc_o[4] (
	.clk(CPUCLK),
	.d(\next_pc_o~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[4] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N21
dffeas \ifid_if.next_pc_o[7] (
	.clk(CPUCLK),
	.d(\next_pc_o~6_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_7),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[7] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N21
dffeas \ifid_if.next_pc_o[6] (
	.clk(CPUCLK),
	.d(\next_pc_o~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_6),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[6] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y29_N23
dffeas \ifid_if.next_pc_o[9] (
	.clk(CPUCLK),
	.d(\next_pc_o~8_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_9),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[9] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y31_N23
dffeas \ifid_if.next_pc_o[8] (
	.clk(CPUCLK),
	.d(\next_pc_o~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_8),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[8] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N5
dffeas \ifid_if.next_pc_o[11] (
	.clk(CPUCLK),
	.d(\next_pc_o~10_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_11),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[11] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N23
dffeas \ifid_if.next_pc_o[10] (
	.clk(CPUCLK),
	.d(\next_pc_o~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_10),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[10] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N27
dffeas \ifid_if.next_pc_o[13] (
	.clk(CPUCLK),
	.d(\next_pc_o~12_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_13),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[13] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N27
dffeas \ifid_if.next_pc_o[12] (
	.clk(CPUCLK),
	.d(\next_pc_o~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_12),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[12] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y29_N29
dffeas \ifid_if.next_pc_o[15] (
	.clk(CPUCLK),
	.d(\next_pc_o~14_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_15),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[15] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N3
dffeas \ifid_if.next_pc_o[14] (
	.clk(CPUCLK),
	.d(\next_pc_o~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_14),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[14] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N21
dffeas \ifid_if.next_pc_o[17] (
	.clk(CPUCLK),
	.d(\next_pc_o~16_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_17),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[17] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y29_N15
dffeas \ifid_if.next_pc_o[16] (
	.clk(CPUCLK),
	.d(\next_pc_o~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_16),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[16] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N25
dffeas \ifid_if.next_pc_o[19] (
	.clk(CPUCLK),
	.d(\next_pc_o~18_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_19),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[19] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N31
dffeas \ifid_if.next_pc_o[18] (
	.clk(CPUCLK),
	.d(\next_pc_o~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_18),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[18] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N7
dffeas \ifid_if.next_pc_o[21] (
	.clk(CPUCLK),
	.d(\next_pc_o~20_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_21),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[21] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N5
dffeas \ifid_if.next_pc_o[20] (
	.clk(CPUCLK),
	.d(\next_pc_o~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_20),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[20] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N15
dffeas \ifid_if.next_pc_o[23] (
	.clk(CPUCLK),
	.d(\next_pc_o~22_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_23),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[23] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N31
dffeas \ifid_if.next_pc_o[22] (
	.clk(CPUCLK),
	.d(\next_pc_o~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_22),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[22] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N9
dffeas \ifid_if.next_pc_o[25] (
	.clk(CPUCLK),
	.d(\next_pc_o~24_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_25),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[25] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N9
dffeas \ifid_if.next_pc_o[24] (
	.clk(CPUCLK),
	.d(\next_pc_o~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_24),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[24] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N23
dffeas \ifid_if.next_pc_o[27] (
	.clk(CPUCLK),
	.d(\next_pc_o~26_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_27),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[27] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N31
dffeas \ifid_if.next_pc_o[26] (
	.clk(CPUCLK),
	.d(\next_pc_o~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_26),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[26] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N3
dffeas \ifid_if.next_pc_o[29] (
	.clk(CPUCLK),
	.d(\next_pc_o~28_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_29),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[29] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y28_N31
dffeas \ifid_if.next_pc_o[28] (
	.clk(CPUCLK),
	.d(\next_pc_o~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_28),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[28] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N13
dffeas \ifid_if.next_pc_o[31] (
	.clk(CPUCLK),
	.d(\next_pc_o~30_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_31),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[31] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N23
dffeas \ifid_if.next_pc_o[30] (
	.clk(CPUCLK),
	.d(\next_pc_o~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ifid_if.instr_o[25]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ifid_ifnext_pc_o_30),
	.prn(vcc));
// synopsys translate_off
defparam \ifid_if.next_pc_o[30] .is_wysiwyg = "true";
defparam \ifid_if.next_pc_o[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N24
cycloneive_lcell_comb \instr_o~0 (
// Equation(s):
// \instr_o~0_combout  = (ramiframload_17 & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(ramiframload_17),
	.datac(always11),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~0 .lut_mask = 16'h0CCC;
defparam \instr_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N30
cycloneive_lcell_comb \ifid_if.instr_o[25]~0 (
// Equation(s):
// \ifid_if.instr_o[25]~0_combout  = (always13 & ((huifflush) # (!huiffreeze)))

	.dataa(always11),
	.datab(huiffreeze),
	.datac(gnd),
	.datad(huifflush),
	.cin(gnd),
	.combout(\ifid_if.instr_o[25]~0_combout ),
	.cout());
// synopsys translate_off
defparam \ifid_if.instr_o[25]~0 .lut_mask = 16'hAA22;
defparam \ifid_if.instr_o[25]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N16
cycloneive_lcell_comb \instr_o~1 (
// Equation(s):
// \instr_o~1_combout  = (ramiframload_16 & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(huifflush),
	.datad(ramiframload_16),
	.cin(gnd),
	.combout(\instr_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~1 .lut_mask = 16'h3F00;
defparam \instr_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N6
cycloneive_lcell_comb \instr_o~2 (
// Equation(s):
// \instr_o~2_combout  = (ramiframload_19 & ((!huifflush) # (!always13)))

	.dataa(always11),
	.datab(ramiframload_19),
	.datac(gnd),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~2 .lut_mask = 16'h44CC;
defparam \instr_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N6
cycloneive_lcell_comb \instr_o~3 (
// Equation(s):
// \instr_o~3_combout  = (ramiframload_18 & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(huifflush),
	.datad(ramiframload_18),
	.cin(gnd),
	.combout(\instr_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~3 .lut_mask = 16'h3F00;
defparam \instr_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N20
cycloneive_lcell_comb \instr_o~4 (
// Equation(s):
// \instr_o~4_combout  = (ramiframload_20 & ((!huifflush) # (!always13)))

	.dataa(ramiframload_20),
	.datab(always11),
	.datac(huifflush),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr_o~4_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~4 .lut_mask = 16'h2A2A;
defparam \instr_o~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N22
cycloneive_lcell_comb \instr_o~5 (
// Equation(s):
// \instr_o~5_combout  = (ramiframload_22 & ((!huifflush) # (!always13)))

	.dataa(ramiframload_22),
	.datab(always11),
	.datac(gnd),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~5_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~5 .lut_mask = 16'h22AA;
defparam \instr_o~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N18
cycloneive_lcell_comb \instr_o~6 (
// Equation(s):
// \instr_o~6_combout  = (ramiframload_21 & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(huifflush),
	.datad(ramiframload_21),
	.cin(gnd),
	.combout(\instr_o~6_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~6 .lut_mask = 16'h3F00;
defparam \instr_o~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N4
cycloneive_lcell_comb \instr_o~7 (
// Equation(s):
// \instr_o~7_combout  = (ramiframload_24 & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(ramiframload_24),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~7_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~7 .lut_mask = 16'h30F0;
defparam \instr_o~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N10
cycloneive_lcell_comb \instr_o~8 (
// Equation(s):
// \instr_o~8_combout  = (ramiframload_23 & ((!huifflush) # (!always13)))

	.dataa(ramiframload_23),
	.datab(always11),
	.datac(gnd),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~8_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~8 .lut_mask = 16'h22AA;
defparam \instr_o~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N24
cycloneive_lcell_comb \instr_o~9 (
// Equation(s):
// \instr_o~9_combout  = (ramiframload_25 & ((!huifflush) # (!always13)))

	.dataa(ramiframload_25),
	.datab(always11),
	.datac(huifflush),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr_o~9_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~9 .lut_mask = 16'h2A2A;
defparam \instr_o~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N24
cycloneive_lcell_comb \instr_o~10 (
// Equation(s):
// \instr_o~10_combout  = (ramiframload_26 & ((!huifflush) # (!always13)))

	.dataa(always11),
	.datab(gnd),
	.datac(ramiframload_26),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~10_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~10 .lut_mask = 16'h50F0;
defparam \instr_o~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N0
cycloneive_lcell_comb \instr_o~11 (
// Equation(s):
// \instr_o~11_combout  = (ramiframload_31 & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(huifflush),
	.datad(ramiframload_31),
	.cin(gnd),
	.combout(\instr_o~11_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~11 .lut_mask = 16'h3F00;
defparam \instr_o~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N30
cycloneive_lcell_comb \instr_o~12 (
// Equation(s):
// \instr_o~12_combout  = (ramiframload_27 & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(huifflush),
	.datad(ramiframload_27),
	.cin(gnd),
	.combout(\instr_o~12_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~12 .lut_mask = 16'h3F00;
defparam \instr_o~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N30
cycloneive_lcell_comb \instr_o~13 (
// Equation(s):
// \instr_o~13_combout  = (ramiframload_28 & ((!huifflush) # (!always13)))

	.dataa(ramiframload_28),
	.datab(always11),
	.datac(gnd),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~13_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~13 .lut_mask = 16'h22AA;
defparam \instr_o~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N2
cycloneive_lcell_comb \instr_o~14 (
// Equation(s):
// \instr_o~14_combout  = (ramiframload_30 & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(huifflush),
	.datad(ramiframload_30),
	.cin(gnd),
	.combout(\instr_o~14_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~14 .lut_mask = 16'h3F00;
defparam \instr_o~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N20
cycloneive_lcell_comb \instr_o~15 (
// Equation(s):
// \instr_o~15_combout  = (ramiframload_5 & ((!huifflush) # (!always13)))

	.dataa(ramiframload_5),
	.datab(gnd),
	.datac(always11),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~15_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~15 .lut_mask = 16'h0AAA;
defparam \instr_o~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N4
cycloneive_lcell_comb \instr_o~16 (
// Equation(s):
// \instr_o~16_combout  = (ramiframload_4 & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(ramiframload_4),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~16_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~16 .lut_mask = 16'h30F0;
defparam \instr_o~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N18
cycloneive_lcell_comb \instr_o~17 (
// Equation(s):
// \instr_o~17_combout  = (ramiframload_29 & ((!huifflush) # (!always13)))

	.dataa(ramiframload_29),
	.datab(always11),
	.datac(gnd),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~17_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~17 .lut_mask = 16'h22AA;
defparam \instr_o~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N12
cycloneive_lcell_comb \instr_o~18 (
// Equation(s):
// \instr_o~18_combout  = (always11 & (ramiframload_1 & ((!huifflush) # (!always13))))

	.dataa(always1),
	.datab(always11),
	.datac(ramiframload_1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~18_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~18 .lut_mask = 16'h20A0;
defparam \instr_o~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N4
cycloneive_lcell_comb \instr_o~19 (
// Equation(s):
// \instr_o~19_combout  = (ramiframload_3 & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(huifflush),
	.datad(ramiframload_3),
	.cin(gnd),
	.combout(\instr_o~19_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~19 .lut_mask = 16'h3F00;
defparam \instr_o~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N18
cycloneive_lcell_comb \instr_o~20 (
// Equation(s):
// \instr_o~20_combout  = (ramiframload_2 & ((!huifflush) # (!always13)))

	.dataa(ramiframload_2),
	.datab(always11),
	.datac(gnd),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~20_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~20 .lut_mask = 16'h22AA;
defparam \instr_o~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N16
cycloneive_lcell_comb \instr_o~21 (
// Equation(s):
// \instr_o~21_combout  = (ramiframload_0 & (((!huifflush)) # (!always13))) # (!ramiframload_0 & (!always11 & ((!huifflush) # (!always13))))

	.dataa(ramiframload_0),
	.datab(always11),
	.datac(always1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~21_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~21 .lut_mask = 16'h23AF;
defparam \instr_o~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N18
cycloneive_lcell_comb \instr_o~22 (
// Equation(s):
// \instr_o~22_combout  = (ramiframload_7 & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(ramiframload_7),
	.datac(always11),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~22_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~22 .lut_mask = 16'h0CCC;
defparam \instr_o~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N24
cycloneive_lcell_comb \instr_o~23 (
// Equation(s):
// \instr_o~23_combout  = (ramiframload_6 & ((!always13) # (!huifflush)))

	.dataa(ramiframload_6),
	.datab(gnd),
	.datac(huifflush),
	.datad(always11),
	.cin(gnd),
	.combout(\instr_o~23_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~23 .lut_mask = 16'h0AAA;
defparam \instr_o~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N4
cycloneive_lcell_comb \instr_o~24 (
// Equation(s):
// \instr_o~24_combout  = (ramiframload_8 & ((!huifflush) # (!always13)))

	.dataa(ramiframload_8),
	.datab(always11),
	.datac(gnd),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~24_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~24 .lut_mask = 16'h22AA;
defparam \instr_o~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N30
cycloneive_lcell_comb \instr_o~25 (
// Equation(s):
// \instr_o~25_combout  = (ramiframload_9 & ((!huifflush) # (!always13)))

	.dataa(ramiframload_9),
	.datab(always11),
	.datac(huifflush),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr_o~25_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~25 .lut_mask = 16'h2A2A;
defparam \instr_o~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N14
cycloneive_lcell_comb \instr_o~26 (
// Equation(s):
// \instr_o~26_combout  = (ramiframload_10 & ((!huifflush) # (!always13)))

	.dataa(ramiframload_10),
	.datab(always11),
	.datac(huifflush),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr_o~26_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~26 .lut_mask = 16'h2A2A;
defparam \instr_o~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N12
cycloneive_lcell_comb \instr_o~27 (
// Equation(s):
// \instr_o~27_combout  = (ramiframload_15 & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(ramiframload_15),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~27_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~27 .lut_mask = 16'h30F0;
defparam \instr_o~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N20
cycloneive_lcell_comb \instr_o~28 (
// Equation(s):
// \instr_o~28_combout  = (ramiframload_14 & ((!always13) # (!huifflush)))

	.dataa(gnd),
	.datab(ramiframload_14),
	.datac(huifflush),
	.datad(always11),
	.cin(gnd),
	.combout(\instr_o~28_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~28 .lut_mask = 16'h0CCC;
defparam \instr_o~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N14
cycloneive_lcell_comb \instr_o~29 (
// Equation(s):
// \instr_o~29_combout  = (ramiframload_111 & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(ramiframload_11),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~29_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~29 .lut_mask = 16'h30F0;
defparam \instr_o~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N4
cycloneive_lcell_comb \instr_o~30 (
// Equation(s):
// \instr_o~30_combout  = (ramiframload_12 & ((!huifflush) # (!always13)))

	.dataa(always11),
	.datab(ramiframload_12),
	.datac(huifflush),
	.datad(gnd),
	.cin(gnd),
	.combout(\instr_o~30_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~30 .lut_mask = 16'h4C4C;
defparam \instr_o~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N8
cycloneive_lcell_comb \instr_o~31 (
// Equation(s):
// \instr_o~31_combout  = (ramiframload_13 & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(ramiframload_13),
	.datad(huifflush),
	.cin(gnd),
	.combout(\instr_o~31_combout ),
	.cout());
// synopsys translate_off
defparam \instr_o~31 .lut_mask = 16'h30F0;
defparam \instr_o~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N30
cycloneive_lcell_comb \next_pc_o~0 (
// Equation(s):
// \next_pc_o~0_combout  = (pc_1 & ((!huifflush) # (!always13)))

	.dataa(always11),
	.datab(gnd),
	.datac(pc_1),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~0_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~0 .lut_mask = 16'h50F0;
defparam \next_pc_o~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N0
cycloneive_lcell_comb \next_pc_o~1 (
// Equation(s):
// \next_pc_o~1_combout  = (pc_0 & ((!huifflush) # (!always13)))

	.dataa(always11),
	.datab(pc_0),
	.datac(gnd),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~1_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~1 .lut_mask = 16'h44CC;
defparam \next_pc_o~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N8
cycloneive_lcell_comb \next_pc_o~2 (
// Equation(s):
// \next_pc_o~2_combout  = (\nextpc[3]~2_combout  & ((!huifflush) # (!always13)))

	.dataa(nextpc_3),
	.datab(always11),
	.datac(huifflush),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pc_o~2_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~2 .lut_mask = 16'h2A2A;
defparam \next_pc_o~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N6
cycloneive_lcell_comb \next_pc_o~3 (
// Equation(s):
// \next_pc_o~3_combout  = (\nextpc[2]~0_combout  & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(nextpc_2),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~3_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~3 .lut_mask = 16'h30F0;
defparam \next_pc_o~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N22
cycloneive_lcell_comb \next_pc_o~4 (
// Equation(s):
// \next_pc_o~4_combout  = (\nextpc[5]~6_combout  & ((!huifflush) # (!always13)))

	.dataa(nextpc_5),
	.datab(always11),
	.datac(huifflush),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pc_o~4_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~4 .lut_mask = 16'h2A2A;
defparam \next_pc_o~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N22
cycloneive_lcell_comb \next_pc_o~5 (
// Equation(s):
// \next_pc_o~5_combout  = (\nextpc[4]~4_combout  & ((!huifflush) # (!always13)))

	.dataa(nextpc_4),
	.datab(gnd),
	.datac(always11),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~5_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~5 .lut_mask = 16'h0AAA;
defparam \next_pc_o~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N20
cycloneive_lcell_comb \next_pc_o~6 (
// Equation(s):
// \next_pc_o~6_combout  = (\nextpc[7]~10_combout  & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(nextpc_7),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~6_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~6 .lut_mask = 16'h30F0;
defparam \next_pc_o~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N20
cycloneive_lcell_comb \next_pc_o~7 (
// Equation(s):
// \next_pc_o~7_combout  = (\nextpc[6]~8_combout  & ((!huifflush) # (!always13)))

	.dataa(nextpc_6),
	.datab(always11),
	.datac(huifflush),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pc_o~7_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~7 .lut_mask = 16'h2A2A;
defparam \next_pc_o~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N22
cycloneive_lcell_comb \next_pc_o~8 (
// Equation(s):
// \next_pc_o~8_combout  = (\nextpc[9]~14_combout  & ((!huifflush) # (!always13)))

	.dataa(always11),
	.datab(gnd),
	.datac(nextpc_9),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~8_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~8 .lut_mask = 16'h50F0;
defparam \next_pc_o~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N22
cycloneive_lcell_comb \next_pc_o~9 (
// Equation(s):
// \next_pc_o~9_combout  = (\nextpc[8]~12_combout  & ((!always13) # (!huifflush)))

	.dataa(nextpc_8),
	.datab(huifflush),
	.datac(always11),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pc_o~9_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~9 .lut_mask = 16'h2A2A;
defparam \next_pc_o~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N4
cycloneive_lcell_comb \next_pc_o~10 (
// Equation(s):
// \next_pc_o~10_combout  = (\nextpc[11]~18_combout  & ((!huifflush) # (!always13)))

	.dataa(nextpc_11),
	.datab(always11),
	.datac(gnd),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~10_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~10 .lut_mask = 16'h22AA;
defparam \next_pc_o~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N22
cycloneive_lcell_comb \next_pc_o~11 (
// Equation(s):
// \next_pc_o~11_combout  = (\nextpc[10]~16_combout  & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(huifflush),
	.datad(nextpc_10),
	.cin(gnd),
	.combout(\next_pc_o~11_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~11 .lut_mask = 16'h3F00;
defparam \next_pc_o~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N26
cycloneive_lcell_comb \next_pc_o~12 (
// Equation(s):
// \next_pc_o~12_combout  = (\nextpc[13]~22_combout  & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(nextpc_13),
	.datac(always11),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~12_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~12 .lut_mask = 16'h0CCC;
defparam \next_pc_o~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N26
cycloneive_lcell_comb \next_pc_o~13 (
// Equation(s):
// \next_pc_o~13_combout  = (\nextpc[12]~20_combout  & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(nextpc_12),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~13_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~13 .lut_mask = 16'h30F0;
defparam \next_pc_o~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N28
cycloneive_lcell_comb \next_pc_o~14 (
// Equation(s):
// \next_pc_o~14_combout  = (\nextpc[15]~26_combout  & ((!huifflush) # (!always13)))

	.dataa(always11),
	.datab(nextpc_15),
	.datac(gnd),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~14_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~14 .lut_mask = 16'h44CC;
defparam \next_pc_o~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N2
cycloneive_lcell_comb \next_pc_o~15 (
// Equation(s):
// \next_pc_o~15_combout  = (\nextpc[14]~24_combout  & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(nextpc_14),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~15_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~15 .lut_mask = 16'h30F0;
defparam \next_pc_o~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N20
cycloneive_lcell_comb \next_pc_o~16 (
// Equation(s):
// \next_pc_o~16_combout  = (\nextpc[17]~30_combout  & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(nextpc_17),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~16_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~16 .lut_mask = 16'h30F0;
defparam \next_pc_o~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N14
cycloneive_lcell_comb \next_pc_o~17 (
// Equation(s):
// \next_pc_o~17_combout  = (\nextpc[16]~28_combout  & ((!huifflush) # (!always13)))

	.dataa(always11),
	.datab(gnd),
	.datac(nextpc_16),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~17_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~17 .lut_mask = 16'h50F0;
defparam \next_pc_o~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N24
cycloneive_lcell_comb \next_pc_o~18 (
// Equation(s):
// \next_pc_o~18_combout  = (\nextpc[19]~34_combout  & ((!huifflush) # (!always13)))

	.dataa(nextpc_19),
	.datab(always11),
	.datac(huifflush),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pc_o~18_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~18 .lut_mask = 16'h2A2A;
defparam \next_pc_o~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N30
cycloneive_lcell_comb \next_pc_o~19 (
// Equation(s):
// \next_pc_o~19_combout  = (\nextpc[18]~32_combout  & ((!huifflush) # (!always13)))

	.dataa(always11),
	.datab(nextpc_18),
	.datac(gnd),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~19_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~19 .lut_mask = 16'h44CC;
defparam \next_pc_o~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N6
cycloneive_lcell_comb \next_pc_o~20 (
// Equation(s):
// \next_pc_o~20_combout  = (\nextpc[21]~38_combout  & ((!huifflush) # (!always13)))

	.dataa(nextpc_21),
	.datab(always11),
	.datac(huifflush),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pc_o~20_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~20 .lut_mask = 16'h2A2A;
defparam \next_pc_o~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N4
cycloneive_lcell_comb \next_pc_o~21 (
// Equation(s):
// \next_pc_o~21_combout  = (\nextpc[20]~36_combout  & ((!huifflush) # (!always13)))

	.dataa(always11),
	.datab(gnd),
	.datac(nextpc_20),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~21_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~21 .lut_mask = 16'h50F0;
defparam \next_pc_o~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N14
cycloneive_lcell_comb \next_pc_o~22 (
// Equation(s):
// \next_pc_o~22_combout  = (\nextpc[23]~42_combout  & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(nextpc_23),
	.datac(always11),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~22_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~22 .lut_mask = 16'h0CCC;
defparam \next_pc_o~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N30
cycloneive_lcell_comb \next_pc_o~23 (
// Equation(s):
// \next_pc_o~23_combout  = (\nextpc[22]~40_combout  & ((!always13) # (!huifflush)))

	.dataa(nextpc_22),
	.datab(huifflush),
	.datac(always11),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pc_o~23_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~23 .lut_mask = 16'h2A2A;
defparam \next_pc_o~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N8
cycloneive_lcell_comb \next_pc_o~24 (
// Equation(s):
// \next_pc_o~24_combout  = (\nextpc[25]~46_combout  & ((!huifflush) # (!always13)))

	.dataa(always11),
	.datab(gnd),
	.datac(nextpc_25),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~24_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~24 .lut_mask = 16'h50F0;
defparam \next_pc_o~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N8
cycloneive_lcell_comb \next_pc_o~25 (
// Equation(s):
// \next_pc_o~25_combout  = (\nextpc[24]~44_combout  & ((!huifflush) # (!always13)))

	.dataa(always11),
	.datab(huifflush),
	.datac(nextpc_24),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pc_o~25_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~25 .lut_mask = 16'h7070;
defparam \next_pc_o~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N22
cycloneive_lcell_comb \next_pc_o~26 (
// Equation(s):
// \next_pc_o~26_combout  = (\nextpc[27]~50_combout  & ((!huifflush) # (!always13)))

	.dataa(always11),
	.datab(huifflush),
	.datac(nextpc_27),
	.datad(gnd),
	.cin(gnd),
	.combout(\next_pc_o~26_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~26 .lut_mask = 16'h7070;
defparam \next_pc_o~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N30
cycloneive_lcell_comb \next_pc_o~27 (
// Equation(s):
// \next_pc_o~27_combout  = (\nextpc[26]~48_combout  & ((!huifflush) # (!always13)))

	.dataa(always11),
	.datab(gnd),
	.datac(nextpc_26),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~27_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~27 .lut_mask = 16'h50F0;
defparam \next_pc_o~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N2
cycloneive_lcell_comb \next_pc_o~28 (
// Equation(s):
// \next_pc_o~28_combout  = (\nextpc[29]~54_combout  & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(always11),
	.datac(nextpc_29),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~28_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~28 .lut_mask = 16'h30F0;
defparam \next_pc_o~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N30
cycloneive_lcell_comb \next_pc_o~29 (
// Equation(s):
// \next_pc_o~29_combout  = (\nextpc[28]~52_combout  & ((!huifflush) # (!always13)))

	.dataa(gnd),
	.datab(nextpc_28),
	.datac(always11),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~29_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~29 .lut_mask = 16'h0CCC;
defparam \next_pc_o~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N12
cycloneive_lcell_comb \next_pc_o~30 (
// Equation(s):
// \next_pc_o~30_combout  = (\nextpc[31]~58_combout  & ((!huifflush) # (!always13)))

	.dataa(nextpc_31),
	.datab(gnd),
	.datac(always11),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~30_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~30 .lut_mask = 16'h0AAA;
defparam \next_pc_o~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N22
cycloneive_lcell_comb \next_pc_o~31 (
// Equation(s):
// \next_pc_o~31_combout  = (\nextpc[30]~56_combout  & ((!huifflush) # (!always13)))

	.dataa(always11),
	.datab(gnd),
	.datac(nextpc_30),
	.datad(huifflush),
	.cin(gnd),
	.combout(\next_pc_o~31_combout ),
	.cout());
// synopsys translate_off
defparam \next_pc_o~31 .lut_mask = 16'h50F0;
defparam \next_pc_o~31 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module mem_wb (
	exmem_ifout_o_1,
	exmem_ifout_o_0,
	exmem_ifout_o_3,
	exmem_ifout_o_2,
	exmem_ifout_o_5,
	exmem_ifout_o_4,
	exmem_ifout_o_7,
	exmem_ifout_o_6,
	exmem_ifout_o_9,
	exmem_ifout_o_8,
	exmem_ifout_o_11,
	exmem_ifout_o_10,
	exmem_ifout_o_13,
	exmem_ifout_o_12,
	exmem_ifout_o_15,
	exmem_ifout_o_14,
	exmem_ifout_o_17,
	exmem_ifout_o_16,
	exmem_ifout_o_19,
	exmem_ifout_o_18,
	exmem_ifout_o_21,
	exmem_ifout_o_20,
	exmem_ifout_o_23,
	exmem_ifout_o_22,
	exmem_ifout_o_25,
	exmem_ifout_o_24,
	exmem_ifout_o_27,
	exmem_ifout_o_26,
	exmem_ifout_o_29,
	exmem_ifout_o_28,
	exmem_ifout_o_31,
	exmem_ifout_o_30,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	exmem_ifRegDest_o_1,
	exmem_ifrt_o_1,
	exmem_ifrd_o_1,
	exmem_ifRegDest_o_0,
	exmem_ifrt_o_0,
	exmem_ifrd_o_0,
	exmem_ifrt_o_3,
	exmem_ifrd_o_3,
	exmem_ifrt_o_2,
	exmem_ifrd_o_2,
	exmem_ifregWEN_o,
	exmem_ifrt_o_4,
	exmem_ifrd_o_4,
	memwb_ifRegDest_o_1,
	memwb_ifrt_o_1,
	memwb_ifrd_o_1,
	memwb_ifRegDest_o_0,
	memwb_ifrt_o_0,
	memwb_ifrd_o_0,
	memwb_ifrt_o_3,
	memwb_ifrd_o_3,
	memwb_ifrt_o_2,
	memwb_ifrd_o_2,
	memwb_ifregWEN_o,
	memwb_ifrt_o_4,
	memwb_ifrd_o_4,
	memwb_ifdmemload_o_1,
	memwb_ifout_o_1,
	memwb_ifmemToReg_o,
	memwb_ifjal_o,
	memwb_ifnext_pc_o_1,
	memwb_iflui_o,
	exmem_ifjal_o,
	exmem_iflui_o,
	exmem_ifnext_pc_o_1,
	exmem_ifmemToReg_o,
	exmem_ifnext_pc_o_0,
	memwb_ifdmemload_o_0,
	memwb_ifout_o_0,
	memwb_ifnext_pc_o_0,
	memwb_ifdmemload_o_2,
	memwb_ifout_o_2,
	memwb_ifnext_pc_o_2,
	exmem_ifnext_pc_o_2,
	memwb_ifdmemload_o_4,
	memwb_ifout_o_4,
	memwb_ifnext_pc_o_4,
	exmem_ifnext_pc_o_4,
	memwb_ifdmemload_o_3,
	memwb_ifout_o_3,
	memwb_ifnext_pc_o_3,
	exmem_ifnext_pc_o_3,
	memwb_ifdmemload_o_8,
	memwb_ifout_o_8,
	memwb_ifnext_pc_o_8,
	exmem_ifnext_pc_o_8,
	memwb_ifdmemload_o_7,
	memwb_ifout_o_7,
	memwb_ifnext_pc_o_7,
	exmem_ifnext_pc_o_7,
	memwb_ifdmemload_o_6,
	memwb_ifout_o_6,
	memwb_ifnext_pc_o_6,
	exmem_ifnext_pc_o_6,
	memwb_ifdmemload_o_5,
	memwb_ifout_o_5,
	memwb_ifnext_pc_o_5,
	exmem_ifnext_pc_o_5,
	memwb_ifdmemload_o_16,
	memwb_ifnext_pc_o_16,
	memwb_ifout_o_16,
	memwb_ifimm_o_0,
	exmem_ifimm_o_0,
	exmem_ifnext_pc_o_16,
	memwb_ifdmemload_o_15,
	memwb_ifout_o_15,
	memwb_ifnext_pc_o_15,
	exmem_ifnext_pc_o_15,
	memwb_ifdmemload_o_14,
	memwb_ifout_o_14,
	memwb_ifnext_pc_o_14,
	exmem_ifnext_pc_o_14,
	memwb_ifdmemload_o_13,
	memwb_ifout_o_13,
	memwb_ifnext_pc_o_13,
	exmem_ifnext_pc_o_13,
	memwb_ifdmemload_o_12,
	memwb_ifout_o_12,
	memwb_ifnext_pc_o_12,
	exmem_ifnext_pc_o_12,
	memwb_ifdmemload_o_11,
	memwb_ifout_o_11,
	memwb_ifnext_pc_o_11,
	exmem_ifnext_pc_o_11,
	memwb_ifdmemload_o_10,
	memwb_ifout_o_10,
	memwb_ifnext_pc_o_10,
	exmem_ifnext_pc_o_10,
	memwb_ifdmemload_o_9,
	memwb_ifout_o_9,
	memwb_ifnext_pc_o_9,
	exmem_ifnext_pc_o_9,
	memwb_ifnext_pc_o_31,
	memwb_ifdmemload_o_31,
	memwb_ifout_o_31,
	memwb_ifimm_o_15,
	exmem_ifnext_pc_o_31,
	exmem_ifimm_o_15,
	memwb_ifnext_pc_o_29,
	memwb_ifdmemload_o_29,
	memwb_ifout_o_29,
	memwb_ifimm_o_13,
	exmem_ifnext_pc_o_29,
	exmem_ifimm_o_13,
	memwb_ifdmemload_o_30,
	memwb_ifnext_pc_o_30,
	memwb_ifout_o_30,
	memwb_ifimm_o_14,
	exmem_ifimm_o_14,
	exmem_ifnext_pc_o_30,
	memwb_ifdmemload_o_28,
	memwb_ifnext_pc_o_28,
	memwb_ifout_o_28,
	memwb_ifimm_o_12,
	exmem_ifimm_o_12,
	exmem_ifnext_pc_o_28,
	memwb_ifdmemload_o_26,
	memwb_ifnext_pc_o_26,
	memwb_ifout_o_26,
	memwb_ifimm_o_10,
	exmem_ifimm_o_10,
	exmem_ifnext_pc_o_26,
	memwb_ifnext_pc_o_27,
	memwb_ifdmemload_o_27,
	memwb_ifout_o_27,
	memwb_ifimm_o_11,
	exmem_ifnext_pc_o_27,
	exmem_ifimm_o_11,
	memwb_ifnext_pc_o_25,
	memwb_ifdmemload_o_25,
	memwb_ifout_o_25,
	memwb_ifimm_o_9,
	exmem_ifnext_pc_o_25,
	exmem_ifimm_o_9,
	memwb_ifdmemload_o_24,
	memwb_ifnext_pc_o_24,
	memwb_ifout_o_24,
	memwb_ifimm_o_8,
	exmem_ifimm_o_8,
	exmem_ifnext_pc_o_24,
	memwb_ifdmemload_o_22,
	memwb_ifnext_pc_o_22,
	memwb_ifout_o_22,
	memwb_ifimm_o_6,
	exmem_ifimm_o_6,
	exmem_ifnext_pc_o_22,
	memwb_ifnext_pc_o_23,
	memwb_ifdmemload_o_23,
	memwb_ifout_o_23,
	memwb_ifimm_o_7,
	exmem_ifnext_pc_o_23,
	exmem_ifimm_o_7,
	memwb_ifnext_pc_o_21,
	memwb_ifdmemload_o_21,
	memwb_ifout_o_21,
	memwb_ifimm_o_5,
	exmem_ifnext_pc_o_21,
	exmem_ifimm_o_5,
	memwb_ifdmemload_o_20,
	memwb_ifnext_pc_o_20,
	memwb_ifout_o_20,
	memwb_ifimm_o_4,
	exmem_ifimm_o_4,
	exmem_ifnext_pc_o_20,
	memwb_ifdmemload_o_18,
	memwb_ifnext_pc_o_18,
	memwb_ifout_o_18,
	memwb_ifimm_o_2,
	exmem_ifimm_o_2,
	exmem_ifnext_pc_o_18,
	memwb_ifnext_pc_o_19,
	memwb_ifdmemload_o_19,
	memwb_ifout_o_19,
	memwb_ifimm_o_3,
	exmem_ifnext_pc_o_19,
	exmem_ifimm_o_3,
	memwb_ifnext_pc_o_17,
	memwb_ifdmemload_o_17,
	memwb_ifout_o_17,
	memwb_ifimm_o_1,
	exmem_ifnext_pc_o_17,
	exmem_ifimm_o_1,
	exmem_ifimm_o_01,
	CPUCLK,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	exmem_ifout_o_1;
input 	exmem_ifout_o_0;
input 	exmem_ifout_o_3;
input 	exmem_ifout_o_2;
input 	exmem_ifout_o_5;
input 	exmem_ifout_o_4;
input 	exmem_ifout_o_7;
input 	exmem_ifout_o_6;
input 	exmem_ifout_o_9;
input 	exmem_ifout_o_8;
input 	exmem_ifout_o_11;
input 	exmem_ifout_o_10;
input 	exmem_ifout_o_13;
input 	exmem_ifout_o_12;
input 	exmem_ifout_o_15;
input 	exmem_ifout_o_14;
input 	exmem_ifout_o_17;
input 	exmem_ifout_o_16;
input 	exmem_ifout_o_19;
input 	exmem_ifout_o_18;
input 	exmem_ifout_o_21;
input 	exmem_ifout_o_20;
input 	exmem_ifout_o_23;
input 	exmem_ifout_o_22;
input 	exmem_ifout_o_25;
input 	exmem_ifout_o_24;
input 	exmem_ifout_o_27;
input 	exmem_ifout_o_26;
input 	exmem_ifout_o_29;
input 	exmem_ifout_o_28;
input 	exmem_ifout_o_31;
input 	exmem_ifout_o_30;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
input 	exmem_ifRegDest_o_1;
input 	exmem_ifrt_o_1;
input 	exmem_ifrd_o_1;
input 	exmem_ifRegDest_o_0;
input 	exmem_ifrt_o_0;
input 	exmem_ifrd_o_0;
input 	exmem_ifrt_o_3;
input 	exmem_ifrd_o_3;
input 	exmem_ifrt_o_2;
input 	exmem_ifrd_o_2;
input 	exmem_ifregWEN_o;
input 	exmem_ifrt_o_4;
input 	exmem_ifrd_o_4;
output 	memwb_ifRegDest_o_1;
output 	memwb_ifrt_o_1;
output 	memwb_ifrd_o_1;
output 	memwb_ifRegDest_o_0;
output 	memwb_ifrt_o_0;
output 	memwb_ifrd_o_0;
output 	memwb_ifrt_o_3;
output 	memwb_ifrd_o_3;
output 	memwb_ifrt_o_2;
output 	memwb_ifrd_o_2;
output 	memwb_ifregWEN_o;
output 	memwb_ifrt_o_4;
output 	memwb_ifrd_o_4;
output 	memwb_ifdmemload_o_1;
output 	memwb_ifout_o_1;
output 	memwb_ifmemToReg_o;
output 	memwb_ifjal_o;
output 	memwb_ifnext_pc_o_1;
output 	memwb_iflui_o;
input 	exmem_ifjal_o;
input 	exmem_iflui_o;
input 	exmem_ifnext_pc_o_1;
input 	exmem_ifmemToReg_o;
input 	exmem_ifnext_pc_o_0;
output 	memwb_ifdmemload_o_0;
output 	memwb_ifout_o_0;
output 	memwb_ifnext_pc_o_0;
output 	memwb_ifdmemload_o_2;
output 	memwb_ifout_o_2;
output 	memwb_ifnext_pc_o_2;
input 	exmem_ifnext_pc_o_2;
output 	memwb_ifdmemload_o_4;
output 	memwb_ifout_o_4;
output 	memwb_ifnext_pc_o_4;
input 	exmem_ifnext_pc_o_4;
output 	memwb_ifdmemload_o_3;
output 	memwb_ifout_o_3;
output 	memwb_ifnext_pc_o_3;
input 	exmem_ifnext_pc_o_3;
output 	memwb_ifdmemload_o_8;
output 	memwb_ifout_o_8;
output 	memwb_ifnext_pc_o_8;
input 	exmem_ifnext_pc_o_8;
output 	memwb_ifdmemload_o_7;
output 	memwb_ifout_o_7;
output 	memwb_ifnext_pc_o_7;
input 	exmem_ifnext_pc_o_7;
output 	memwb_ifdmemload_o_6;
output 	memwb_ifout_o_6;
output 	memwb_ifnext_pc_o_6;
input 	exmem_ifnext_pc_o_6;
output 	memwb_ifdmemload_o_5;
output 	memwb_ifout_o_5;
output 	memwb_ifnext_pc_o_5;
input 	exmem_ifnext_pc_o_5;
output 	memwb_ifdmemload_o_16;
output 	memwb_ifnext_pc_o_16;
output 	memwb_ifout_o_16;
output 	memwb_ifimm_o_0;
input 	exmem_ifimm_o_0;
input 	exmem_ifnext_pc_o_16;
output 	memwb_ifdmemload_o_15;
output 	memwb_ifout_o_15;
output 	memwb_ifnext_pc_o_15;
input 	exmem_ifnext_pc_o_15;
output 	memwb_ifdmemload_o_14;
output 	memwb_ifout_o_14;
output 	memwb_ifnext_pc_o_14;
input 	exmem_ifnext_pc_o_14;
output 	memwb_ifdmemload_o_13;
output 	memwb_ifout_o_13;
output 	memwb_ifnext_pc_o_13;
input 	exmem_ifnext_pc_o_13;
output 	memwb_ifdmemload_o_12;
output 	memwb_ifout_o_12;
output 	memwb_ifnext_pc_o_12;
input 	exmem_ifnext_pc_o_12;
output 	memwb_ifdmemload_o_11;
output 	memwb_ifout_o_11;
output 	memwb_ifnext_pc_o_11;
input 	exmem_ifnext_pc_o_11;
output 	memwb_ifdmemload_o_10;
output 	memwb_ifout_o_10;
output 	memwb_ifnext_pc_o_10;
input 	exmem_ifnext_pc_o_10;
output 	memwb_ifdmemload_o_9;
output 	memwb_ifout_o_9;
output 	memwb_ifnext_pc_o_9;
input 	exmem_ifnext_pc_o_9;
output 	memwb_ifnext_pc_o_31;
output 	memwb_ifdmemload_o_31;
output 	memwb_ifout_o_31;
output 	memwb_ifimm_o_15;
input 	exmem_ifnext_pc_o_31;
input 	exmem_ifimm_o_15;
output 	memwb_ifnext_pc_o_29;
output 	memwb_ifdmemload_o_29;
output 	memwb_ifout_o_29;
output 	memwb_ifimm_o_13;
input 	exmem_ifnext_pc_o_29;
input 	exmem_ifimm_o_13;
output 	memwb_ifdmemload_o_30;
output 	memwb_ifnext_pc_o_30;
output 	memwb_ifout_o_30;
output 	memwb_ifimm_o_14;
input 	exmem_ifimm_o_14;
input 	exmem_ifnext_pc_o_30;
output 	memwb_ifdmemload_o_28;
output 	memwb_ifnext_pc_o_28;
output 	memwb_ifout_o_28;
output 	memwb_ifimm_o_12;
input 	exmem_ifimm_o_12;
input 	exmem_ifnext_pc_o_28;
output 	memwb_ifdmemload_o_26;
output 	memwb_ifnext_pc_o_26;
output 	memwb_ifout_o_26;
output 	memwb_ifimm_o_10;
input 	exmem_ifimm_o_10;
input 	exmem_ifnext_pc_o_26;
output 	memwb_ifnext_pc_o_27;
output 	memwb_ifdmemload_o_27;
output 	memwb_ifout_o_27;
output 	memwb_ifimm_o_11;
input 	exmem_ifnext_pc_o_27;
input 	exmem_ifimm_o_11;
output 	memwb_ifnext_pc_o_25;
output 	memwb_ifdmemload_o_25;
output 	memwb_ifout_o_25;
output 	memwb_ifimm_o_9;
input 	exmem_ifnext_pc_o_25;
input 	exmem_ifimm_o_9;
output 	memwb_ifdmemload_o_24;
output 	memwb_ifnext_pc_o_24;
output 	memwb_ifout_o_24;
output 	memwb_ifimm_o_8;
input 	exmem_ifimm_o_8;
input 	exmem_ifnext_pc_o_24;
output 	memwb_ifdmemload_o_22;
output 	memwb_ifnext_pc_o_22;
output 	memwb_ifout_o_22;
output 	memwb_ifimm_o_6;
input 	exmem_ifimm_o_6;
input 	exmem_ifnext_pc_o_22;
output 	memwb_ifnext_pc_o_23;
output 	memwb_ifdmemload_o_23;
output 	memwb_ifout_o_23;
output 	memwb_ifimm_o_7;
input 	exmem_ifnext_pc_o_23;
input 	exmem_ifimm_o_7;
output 	memwb_ifnext_pc_o_21;
output 	memwb_ifdmemload_o_21;
output 	memwb_ifout_o_21;
output 	memwb_ifimm_o_5;
input 	exmem_ifnext_pc_o_21;
input 	exmem_ifimm_o_5;
output 	memwb_ifdmemload_o_20;
output 	memwb_ifnext_pc_o_20;
output 	memwb_ifout_o_20;
output 	memwb_ifimm_o_4;
input 	exmem_ifimm_o_4;
input 	exmem_ifnext_pc_o_20;
output 	memwb_ifdmemload_o_18;
output 	memwb_ifnext_pc_o_18;
output 	memwb_ifout_o_18;
output 	memwb_ifimm_o_2;
input 	exmem_ifimm_o_2;
input 	exmem_ifnext_pc_o_18;
output 	memwb_ifnext_pc_o_19;
output 	memwb_ifdmemload_o_19;
output 	memwb_ifout_o_19;
output 	memwb_ifimm_o_3;
input 	exmem_ifnext_pc_o_19;
input 	exmem_ifimm_o_3;
output 	memwb_ifnext_pc_o_17;
output 	memwb_ifdmemload_o_17;
output 	memwb_ifout_o_17;
output 	memwb_ifimm_o_1;
input 	exmem_ifnext_pc_o_17;
input 	exmem_ifimm_o_1;
input 	exmem_ifimm_o_01;
input 	CPUCLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \memwb_if.RegDest_o[1]~feeder_combout ;
wire \memwb_if.rt_o[1]~feeder_combout ;
wire \memwb_if.RegDest_o[0]~feeder_combout ;
wire \memwb_if.rt_o[0]~feeder_combout ;
wire \memwb_if.rt_o[3]~feeder_combout ;
wire \memwb_if.rt_o[2]~feeder_combout ;
wire \memwb_if.rt_o[4]~feeder_combout ;
wire \memwb_if.memToReg_o~feeder_combout ;
wire \memwb_if.jal_o~feeder_combout ;
wire \memwb_if.lui_o~feeder_combout ;
wire \memwb_if.dmemload_o[0]~feeder_combout ;
wire \memwb_if.dmemload_o[2]~feeder_combout ;
wire \memwb_if.dmemload_o[4]~feeder_combout ;
wire \memwb_if.next_pc_o[4]~feeder_combout ;
wire \memwb_if.dmemload_o[3]~feeder_combout ;
wire \memwb_if.dmemload_o[7]~feeder_combout ;
wire \memwb_if.next_pc_o[7]~feeder_combout ;
wire \memwb_if.dmemload_o[6]~feeder_combout ;
wire \memwb_if.dmemload_o[5]~feeder_combout ;
wire \memwb_if.next_pc_o[5]~feeder_combout ;
wire \memwb_if.dmemload_o[16]~feeder_combout ;
wire \memwb_if.next_pc_o[16]~feeder_combout ;
wire \memwb_if.dmemload_o[15]~feeder_combout ;
wire \memwb_if.dmemload_o[14]~feeder_combout ;
wire \memwb_if.dmemload_o[13]~feeder_combout ;
wire \memwb_if.dmemload_o[10]~feeder_combout ;
wire \memwb_if.dmemload_o[9]~feeder_combout ;
wire \memwb_if.dmemload_o[31]~feeder_combout ;
wire \memwb_if.dmemload_o[29]~feeder_combout ;
wire \memwb_if.imm_o[13]~feeder_combout ;
wire \memwb_if.next_pc_o[30]~feeder_combout ;
wire \memwb_if.imm_o[14]~feeder_combout ;
wire \memwb_if.dmemload_o[27]~feeder_combout ;
wire \memwb_if.imm_o[11]~feeder_combout ;
wire \memwb_if.dmemload_o[25]~feeder_combout ;
wire \memwb_if.next_pc_o[24]~feeder_combout ;
wire \memwb_if.imm_o[8]~feeder_combout ;
wire \memwb_if.dmemload_o[23]~feeder_combout ;
wire \memwb_if.imm_o[7]~feeder_combout ;
wire \memwb_if.dmemload_o[21]~feeder_combout ;
wire \memwb_if.imm_o[5]~feeder_combout ;
wire \memwb_if.next_pc_o[20]~feeder_combout ;
wire \memwb_if.imm_o[4]~feeder_combout ;
wire \memwb_if.next_pc_o[18]~feeder_combout ;
wire \memwb_if.imm_o[2]~feeder_combout ;
wire \memwb_if.dmemload_o[19]~feeder_combout ;
wire \memwb_if.next_pc_o[17]~feeder_combout ;
wire \memwb_if.dmemload_o[17]~feeder_combout ;


// Location: FF_X53_Y35_N29
dffeas \memwb_if.RegDest_o[1] (
	.clk(CPUCLK),
	.d(\memwb_if.RegDest_o[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifRegDest_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.RegDest_o[1] .is_wysiwyg = "true";
defparam \memwb_if.RegDest_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N19
dffeas \memwb_if.rt_o[1] (
	.clk(CPUCLK),
	.d(\memwb_if.rt_o[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifrt_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.rt_o[1] .is_wysiwyg = "true";
defparam \memwb_if.rt_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N17
dffeas \memwb_if.rd_o[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifrd_o_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifrd_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.rd_o[1] .is_wysiwyg = "true";
defparam \memwb_if.rd_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N23
dffeas \memwb_if.RegDest_o[0] (
	.clk(CPUCLK),
	.d(\memwb_if.RegDest_o[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifRegDest_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.RegDest_o[0] .is_wysiwyg = "true";
defparam \memwb_if.RegDest_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N25
dffeas \memwb_if.rt_o[0] (
	.clk(CPUCLK),
	.d(\memwb_if.rt_o[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifrt_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.rt_o[0] .is_wysiwyg = "true";
defparam \memwb_if.rt_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N15
dffeas \memwb_if.rd_o[0] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifrd_o_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifrd_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.rd_o[0] .is_wysiwyg = "true";
defparam \memwb_if.rd_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N1
dffeas \memwb_if.rt_o[3] (
	.clk(CPUCLK),
	.d(\memwb_if.rt_o[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifrt_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.rt_o[3] .is_wysiwyg = "true";
defparam \memwb_if.rt_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N11
dffeas \memwb_if.rd_o[3] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifrd_o_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifrd_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.rd_o[3] .is_wysiwyg = "true";
defparam \memwb_if.rd_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N13
dffeas \memwb_if.rt_o[2] (
	.clk(CPUCLK),
	.d(\memwb_if.rt_o[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifrt_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.rt_o[2] .is_wysiwyg = "true";
defparam \memwb_if.rt_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N7
dffeas \memwb_if.rd_o[2] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifrd_o_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifrd_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.rd_o[2] .is_wysiwyg = "true";
defparam \memwb_if.rd_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N7
dffeas \memwb_if.regWEN_o (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifregWEN_o),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifregWEN_o),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.regWEN_o .is_wysiwyg = "true";
defparam \memwb_if.regWEN_o .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N5
dffeas \memwb_if.rt_o[4] (
	.clk(CPUCLK),
	.d(\memwb_if.rt_o[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifrt_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.rt_o[4] .is_wysiwyg = "true";
defparam \memwb_if.rt_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N3
dffeas \memwb_if.rd_o[4] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifrd_o_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifrd_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.rd_o[4] .is_wysiwyg = "true";
defparam \memwb_if.rd_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N9
dffeas \memwb_if.dmemload_o[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[1] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N19
dffeas \memwb_if.out_o[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[1] .is_wysiwyg = "true";
defparam \memwb_if.out_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N21
dffeas \memwb_if.memToReg_o (
	.clk(CPUCLK),
	.d(\memwb_if.memToReg_o~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifmemToReg_o),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.memToReg_o .is_wysiwyg = "true";
defparam \memwb_if.memToReg_o .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N23
dffeas \memwb_if.jal_o (
	.clk(CPUCLK),
	.d(\memwb_if.jal_o~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifjal_o),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.jal_o .is_wysiwyg = "true";
defparam \memwb_if.jal_o .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N29
dffeas \memwb_if.next_pc_o[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[1] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N9
dffeas \memwb_if.lui_o (
	.clk(CPUCLK),
	.d(\memwb_if.lui_o~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_iflui_o),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.lui_o .is_wysiwyg = "true";
defparam \memwb_if.lui_o .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N29
dffeas \memwb_if.dmemload_o[0] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[0] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N19
dffeas \memwb_if.out_o[0] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[0] .is_wysiwyg = "true";
defparam \memwb_if.out_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N21
dffeas \memwb_if.next_pc_o[0] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[0] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N3
dffeas \memwb_if.dmemload_o[2] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[2] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N13
dffeas \memwb_if.out_o[2] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[2] .is_wysiwyg = "true";
defparam \memwb_if.out_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N31
dffeas \memwb_if.next_pc_o[2] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[2] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N23
dffeas \memwb_if.dmemload_o[4] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[4] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N9
dffeas \memwb_if.out_o[4] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[4] .is_wysiwyg = "true";
defparam \memwb_if.out_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N17
dffeas \memwb_if.next_pc_o[4] (
	.clk(CPUCLK),
	.d(\memwb_if.next_pc_o[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[4] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N31
dffeas \memwb_if.dmemload_o[3] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[3] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N17
dffeas \memwb_if.out_o[3] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[3] .is_wysiwyg = "true";
defparam \memwb_if.out_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N27
dffeas \memwb_if.next_pc_o[3] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[3] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N23
dffeas \memwb_if.dmemload_o[8] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_8),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[8] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N3
dffeas \memwb_if.out_o[8] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_8),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[8] .is_wysiwyg = "true";
defparam \memwb_if.out_o[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N7
dffeas \memwb_if.next_pc_o[8] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_8),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[8] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N5
dffeas \memwb_if.dmemload_o[7] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_7),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[7] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N15
dffeas \memwb_if.out_o[7] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_7),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[7] .is_wysiwyg = "true";
defparam \memwb_if.out_o[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N3
dffeas \memwb_if.next_pc_o[7] (
	.clk(CPUCLK),
	.d(\memwb_if.next_pc_o[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_7),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[7] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N21
dffeas \memwb_if.dmemload_o[6] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_6),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[6] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N7
dffeas \memwb_if.out_o[6] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_6),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[6] .is_wysiwyg = "true";
defparam \memwb_if.out_o[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N5
dffeas \memwb_if.next_pc_o[6] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_6),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[6] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N7
dffeas \memwb_if.dmemload_o[5] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_5),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[5] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N25
dffeas \memwb_if.out_o[5] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_5),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[5] .is_wysiwyg = "true";
defparam \memwb_if.out_o[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N17
dffeas \memwb_if.next_pc_o[5] (
	.clk(CPUCLK),
	.d(\memwb_if.next_pc_o[5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_5),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[5] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N1
dffeas \memwb_if.dmemload_o[16] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_16),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[16] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N31
dffeas \memwb_if.next_pc_o[16] (
	.clk(CPUCLK),
	.d(\memwb_if.next_pc_o[16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_16),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[16] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N27
dffeas \memwb_if.out_o[16] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_16),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[16] .is_wysiwyg = "true";
defparam \memwb_if.out_o[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N5
dffeas \memwb_if.imm_o[0] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifimm_o_0),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifimm_o_0),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.imm_o[0] .is_wysiwyg = "true";
defparam \memwb_if.imm_o[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N11
dffeas \memwb_if.dmemload_o[15] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_15),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[15] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N9
dffeas \memwb_if.out_o[15] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_15),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[15] .is_wysiwyg = "true";
defparam \memwb_if.out_o[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N29
dffeas \memwb_if.next_pc_o[15] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_15),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[15] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N5
dffeas \memwb_if.dmemload_o[14] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_14),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[14] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N19
dffeas \memwb_if.out_o[14] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_14),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[14] .is_wysiwyg = "true";
defparam \memwb_if.out_o[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N1
dffeas \memwb_if.next_pc_o[14] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_14),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[14] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N7
dffeas \memwb_if.dmemload_o[13] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_13),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[13] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N11
dffeas \memwb_if.out_o[13] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_13),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[13] .is_wysiwyg = "true";
defparam \memwb_if.out_o[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N21
dffeas \memwb_if.next_pc_o[13] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_13),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[13] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N29
dffeas \memwb_if.dmemload_o[12] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_12),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[12] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N21
dffeas \memwb_if.out_o[12] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_12),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[12] .is_wysiwyg = "true";
defparam \memwb_if.out_o[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N9
dffeas \memwb_if.next_pc_o[12] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_12),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[12] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N7
dffeas \memwb_if.dmemload_o[11] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_11),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[11] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N11
dffeas \memwb_if.out_o[11] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_11),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[11] .is_wysiwyg = "true";
defparam \memwb_if.out_o[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y38_N29
dffeas \memwb_if.next_pc_o[11] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_11),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[11] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N19
dffeas \memwb_if.dmemload_o[10] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_10),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[10] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N13
dffeas \memwb_if.out_o[10] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_10),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[10] .is_wysiwyg = "true";
defparam \memwb_if.out_o[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y34_N27
dffeas \memwb_if.next_pc_o[10] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_10),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[10] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N19
dffeas \memwb_if.dmemload_o[9] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_9),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[9] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N23
dffeas \memwb_if.out_o[9] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_9),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[9] .is_wysiwyg = "true";
defparam \memwb_if.out_o[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N5
dffeas \memwb_if.next_pc_o[9] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_9),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[9] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N3
dffeas \memwb_if.next_pc_o[31] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_31),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[31] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N1
dffeas \memwb_if.dmemload_o[31] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_31),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[31] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N19
dffeas \memwb_if.out_o[31] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_31),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[31] .is_wysiwyg = "true";
defparam \memwb_if.out_o[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N11
dffeas \memwb_if.imm_o[15] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifimm_o_15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifimm_o_15),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.imm_o[15] .is_wysiwyg = "true";
defparam \memwb_if.imm_o[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N13
dffeas \memwb_if.next_pc_o[29] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_29),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[29] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N25
dffeas \memwb_if.dmemload_o[29] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_29),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[29] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N17
dffeas \memwb_if.out_o[29] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_29),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[29] .is_wysiwyg = "true";
defparam \memwb_if.out_o[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N7
dffeas \memwb_if.imm_o[13] (
	.clk(CPUCLK),
	.d(\memwb_if.imm_o[13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifimm_o_13),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.imm_o[13] .is_wysiwyg = "true";
defparam \memwb_if.imm_o[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N31
dffeas \memwb_if.dmemload_o[30] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_30),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[30] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N21
dffeas \memwb_if.next_pc_o[30] (
	.clk(CPUCLK),
	.d(\memwb_if.next_pc_o[30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_30),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[30] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N29
dffeas \memwb_if.out_o[30] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_30),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[30] .is_wysiwyg = "true";
defparam \memwb_if.out_o[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N19
dffeas \memwb_if.imm_o[14] (
	.clk(CPUCLK),
	.d(\memwb_if.imm_o[14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifimm_o_14),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.imm_o[14] .is_wysiwyg = "true";
defparam \memwb_if.imm_o[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N23
dffeas \memwb_if.dmemload_o[28] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_28),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[28] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N17
dffeas \memwb_if.next_pc_o[28] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_28),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[28] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N1
dffeas \memwb_if.out_o[28] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_28),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[28] .is_wysiwyg = "true";
defparam \memwb_if.out_o[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N19
dffeas \memwb_if.imm_o[12] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifimm_o_12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifimm_o_12),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.imm_o[12] .is_wysiwyg = "true";
defparam \memwb_if.imm_o[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N21
dffeas \memwb_if.dmemload_o[26] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_26),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[26] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N3
dffeas \memwb_if.next_pc_o[26] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_26),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[26] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y36_N25
dffeas \memwb_if.out_o[26] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_26),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[26] .is_wysiwyg = "true";
defparam \memwb_if.out_o[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N7
dffeas \memwb_if.imm_o[10] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifimm_o_10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifimm_o_10),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.imm_o[10] .is_wysiwyg = "true";
defparam \memwb_if.imm_o[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N17
dffeas \memwb_if.next_pc_o[27] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_27),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[27] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N19
dffeas \memwb_if.dmemload_o[27] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_27),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[27] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N21
dffeas \memwb_if.out_o[27] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_27),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[27] .is_wysiwyg = "true";
defparam \memwb_if.out_o[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N23
dffeas \memwb_if.imm_o[11] (
	.clk(CPUCLK),
	.d(\memwb_if.imm_o[11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifimm_o_11),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.imm_o[11] .is_wysiwyg = "true";
defparam \memwb_if.imm_o[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N25
dffeas \memwb_if.next_pc_o[25] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_25),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[25] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N3
dffeas \memwb_if.dmemload_o[25] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_25),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[25] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N1
dffeas \memwb_if.out_o[25] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_25),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[25] .is_wysiwyg = "true";
defparam \memwb_if.out_o[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N11
dffeas \memwb_if.imm_o[9] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifimm_o_9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifimm_o_9),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.imm_o[9] .is_wysiwyg = "true";
defparam \memwb_if.imm_o[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N29
dffeas \memwb_if.dmemload_o[24] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_24),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[24] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N23
dffeas \memwb_if.next_pc_o[24] (
	.clk(CPUCLK),
	.d(\memwb_if.next_pc_o[24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_24),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[24] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N21
dffeas \memwb_if.out_o[24] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_24),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[24] .is_wysiwyg = "true";
defparam \memwb_if.out_o[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N29
dffeas \memwb_if.imm_o[8] (
	.clk(CPUCLK),
	.d(\memwb_if.imm_o[8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifimm_o_8),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.imm_o[8] .is_wysiwyg = "true";
defparam \memwb_if.imm_o[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N21
dffeas \memwb_if.dmemload_o[22] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_22),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[22] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N19
dffeas \memwb_if.next_pc_o[22] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_22),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[22] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N5
dffeas \memwb_if.out_o[22] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_22),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[22] .is_wysiwyg = "true";
defparam \memwb_if.out_o[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N17
dffeas \memwb_if.imm_o[6] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifimm_o_6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifimm_o_6),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.imm_o[6] .is_wysiwyg = "true";
defparam \memwb_if.imm_o[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N27
dffeas \memwb_if.next_pc_o[23] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_23),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[23] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N13
dffeas \memwb_if.dmemload_o[23] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_23),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[23] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N11
dffeas \memwb_if.out_o[23] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_23),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[23] .is_wysiwyg = "true";
defparam \memwb_if.out_o[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N29
dffeas \memwb_if.imm_o[7] (
	.clk(CPUCLK),
	.d(\memwb_if.imm_o[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifimm_o_7),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.imm_o[7] .is_wysiwyg = "true";
defparam \memwb_if.imm_o[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N27
dffeas \memwb_if.next_pc_o[21] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_21),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[21] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N17
dffeas \memwb_if.dmemload_o[21] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_21),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[21] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N15
dffeas \memwb_if.out_o[21] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_21),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[21] .is_wysiwyg = "true";
defparam \memwb_if.out_o[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N13
dffeas \memwb_if.imm_o[5] (
	.clk(CPUCLK),
	.d(\memwb_if.imm_o[5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifimm_o_5),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.imm_o[5] .is_wysiwyg = "true";
defparam \memwb_if.imm_o[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N31
dffeas \memwb_if.dmemload_o[20] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_20),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[20] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N9
dffeas \memwb_if.next_pc_o[20] (
	.clk(CPUCLK),
	.d(\memwb_if.next_pc_o[20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_20),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[20] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N19
dffeas \memwb_if.out_o[20] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_20),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[20] .is_wysiwyg = "true";
defparam \memwb_if.out_o[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N25
dffeas \memwb_if.imm_o[4] (
	.clk(CPUCLK),
	.d(\memwb_if.imm_o[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifimm_o_4),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.imm_o[4] .is_wysiwyg = "true";
defparam \memwb_if.imm_o[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N7
dffeas \memwb_if.dmemload_o[18] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(ramiframload_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_18),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[18] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N21
dffeas \memwb_if.next_pc_o[18] (
	.clk(CPUCLK),
	.d(\memwb_if.next_pc_o[18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_18),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[18] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N27
dffeas \memwb_if.out_o[18] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_18),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[18] .is_wysiwyg = "true";
defparam \memwb_if.out_o[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N1
dffeas \memwb_if.imm_o[2] (
	.clk(CPUCLK),
	.d(\memwb_if.imm_o[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifimm_o_2),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.imm_o[2] .is_wysiwyg = "true";
defparam \memwb_if.imm_o[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N3
dffeas \memwb_if.next_pc_o[19] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifnext_pc_o_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_19),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[19] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N3
dffeas \memwb_if.dmemload_o[19] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_19),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[19] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y38_N13
dffeas \memwb_if.out_o[19] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_19),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[19] .is_wysiwyg = "true";
defparam \memwb_if.out_o[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y30_N21
dffeas \memwb_if.imm_o[3] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifimm_o_3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifimm_o_3),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.imm_o[3] .is_wysiwyg = "true";
defparam \memwb_if.imm_o[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N17
dffeas \memwb_if.next_pc_o[17] (
	.clk(CPUCLK),
	.d(\memwb_if.next_pc_o[17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifnext_pc_o_17),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.next_pc_o[17] .is_wysiwyg = "true";
defparam \memwb_if.next_pc_o[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N17
dffeas \memwb_if.dmemload_o[17] (
	.clk(CPUCLK),
	.d(\memwb_if.dmemload_o[17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifdmemload_o_17),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.dmemload_o[17] .is_wysiwyg = "true";
defparam \memwb_if.dmemload_o[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N31
dffeas \memwb_if.out_o[17] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifout_o_17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifout_o_17),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.out_o[17] .is_wysiwyg = "true";
defparam \memwb_if.out_o[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N17
dffeas \memwb_if.imm_o[1] (
	.clk(CPUCLK),
	.d(gnd),
	.asdata(exmem_ifimm_o_1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(exmem_ifimm_o_01),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(memwb_ifimm_o_1),
	.prn(vcc));
// synopsys translate_off
defparam \memwb_if.imm_o[1] .is_wysiwyg = "true";
defparam \memwb_if.imm_o[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N28
cycloneive_lcell_comb \memwb_if.RegDest_o[1]~feeder (
// Equation(s):
// \memwb_if.RegDest_o[1]~feeder_combout  = exmem_ifRegDest_o_1

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifRegDest_o_1),
	.cin(gnd),
	.combout(\memwb_if.RegDest_o[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.RegDest_o[1]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.RegDest_o[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N18
cycloneive_lcell_comb \memwb_if.rt_o[1]~feeder (
// Equation(s):
// \memwb_if.rt_o[1]~feeder_combout  = exmem_ifrt_o_1

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifrt_o_1),
	.cin(gnd),
	.combout(\memwb_if.rt_o[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.rt_o[1]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.rt_o[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N22
cycloneive_lcell_comb \memwb_if.RegDest_o[0]~feeder (
// Equation(s):
// \memwb_if.RegDest_o[0]~feeder_combout  = exmem_ifRegDest_o_0

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifRegDest_o_0),
	.cin(gnd),
	.combout(\memwb_if.RegDest_o[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.RegDest_o[0]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.RegDest_o[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N24
cycloneive_lcell_comb \memwb_if.rt_o[0]~feeder (
// Equation(s):
// \memwb_if.rt_o[0]~feeder_combout  = exmem_ifrt_o_0

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifrt_o_0),
	.cin(gnd),
	.combout(\memwb_if.rt_o[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.rt_o[0]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.rt_o[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N0
cycloneive_lcell_comb \memwb_if.rt_o[3]~feeder (
// Equation(s):
// \memwb_if.rt_o[3]~feeder_combout  = exmem_ifrt_o_3

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifrt_o_3),
	.cin(gnd),
	.combout(\memwb_if.rt_o[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.rt_o[3]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.rt_o[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N12
cycloneive_lcell_comb \memwb_if.rt_o[2]~feeder (
// Equation(s):
// \memwb_if.rt_o[2]~feeder_combout  = exmem_ifrt_o_2

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifrt_o_2),
	.cin(gnd),
	.combout(\memwb_if.rt_o[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.rt_o[2]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.rt_o[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N4
cycloneive_lcell_comb \memwb_if.rt_o[4]~feeder (
// Equation(s):
// \memwb_if.rt_o[4]~feeder_combout  = exmem_ifrt_o_4

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifrt_o_4),
	.cin(gnd),
	.combout(\memwb_if.rt_o[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.rt_o[4]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.rt_o[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N20
cycloneive_lcell_comb \memwb_if.memToReg_o~feeder (
// Equation(s):
// \memwb_if.memToReg_o~feeder_combout  = exmem_ifmemToReg_o

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifmemToReg_o),
	.cin(gnd),
	.combout(\memwb_if.memToReg_o~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.memToReg_o~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.memToReg_o~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N22
cycloneive_lcell_comb \memwb_if.jal_o~feeder (
// Equation(s):
// \memwb_if.jal_o~feeder_combout  = exmem_ifjal_o

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifjal_o),
	.cin(gnd),
	.combout(\memwb_if.jal_o~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.jal_o~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.jal_o~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N8
cycloneive_lcell_comb \memwb_if.lui_o~feeder (
// Equation(s):
// \memwb_if.lui_o~feeder_combout  = exmem_iflui_o

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_iflui_o),
	.cin(gnd),
	.combout(\memwb_if.lui_o~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.lui_o~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.lui_o~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N28
cycloneive_lcell_comb \memwb_if.dmemload_o[0]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[0]~feeder_combout  = ramiframload_01

	.dataa(ramiframload_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[0]~feeder .lut_mask = 16'hAAAA;
defparam \memwb_if.dmemload_o[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N2
cycloneive_lcell_comb \memwb_if.dmemload_o[2]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[2]~feeder_combout  = ramiframload_2

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_2),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[2]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.dmemload_o[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N22
cycloneive_lcell_comb \memwb_if.dmemload_o[4]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[4]~feeder_combout  = ramiframload_4

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_4),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[4]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.dmemload_o[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N16
cycloneive_lcell_comb \memwb_if.next_pc_o[4]~feeder (
// Equation(s):
// \memwb_if.next_pc_o[4]~feeder_combout  = exmem_ifnext_pc_o_4

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifnext_pc_o_4),
	.cin(gnd),
	.combout(\memwb_if.next_pc_o[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.next_pc_o[4]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.next_pc_o[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N30
cycloneive_lcell_comb \memwb_if.dmemload_o[3]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[3]~feeder_combout  = ramiframload_3

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_3),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[3]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.dmemload_o[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N4
cycloneive_lcell_comb \memwb_if.dmemload_o[7]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[7]~feeder_combout  = ramiframload_7

	.dataa(ramiframload_7),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[7]~feeder .lut_mask = 16'hAAAA;
defparam \memwb_if.dmemload_o[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N2
cycloneive_lcell_comb \memwb_if.next_pc_o[7]~feeder (
// Equation(s):
// \memwb_if.next_pc_o[7]~feeder_combout  = exmem_ifnext_pc_o_7

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifnext_pc_o_7),
	.cin(gnd),
	.combout(\memwb_if.next_pc_o[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.next_pc_o[7]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.next_pc_o[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N20
cycloneive_lcell_comb \memwb_if.dmemload_o[6]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[6]~feeder_combout  = ramiframload_6

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_6),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[6]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.dmemload_o[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N6
cycloneive_lcell_comb \memwb_if.dmemload_o[5]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[5]~feeder_combout  = ramiframload_5

	.dataa(ramiframload_5),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[5]~feeder .lut_mask = 16'hAAAA;
defparam \memwb_if.dmemload_o[5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N16
cycloneive_lcell_comb \memwb_if.next_pc_o[5]~feeder (
// Equation(s):
// \memwb_if.next_pc_o[5]~feeder_combout  = exmem_ifnext_pc_o_5

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifnext_pc_o_5),
	.cin(gnd),
	.combout(\memwb_if.next_pc_o[5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.next_pc_o[5]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.next_pc_o[5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N0
cycloneive_lcell_comb \memwb_if.dmemload_o[16]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[16]~feeder_combout  = ramiframload_16

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_16),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[16]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.dmemload_o[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N30
cycloneive_lcell_comb \memwb_if.next_pc_o[16]~feeder (
// Equation(s):
// \memwb_if.next_pc_o[16]~feeder_combout  = exmem_ifnext_pc_o_16

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifnext_pc_o_16),
	.cin(gnd),
	.combout(\memwb_if.next_pc_o[16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.next_pc_o[16]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.next_pc_o[16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N10
cycloneive_lcell_comb \memwb_if.dmemload_o[15]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[15]~feeder_combout  = ramiframload_15

	.dataa(gnd),
	.datab(gnd),
	.datac(ramiframload_15),
	.datad(gnd),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[15]~feeder .lut_mask = 16'hF0F0;
defparam \memwb_if.dmemload_o[15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N4
cycloneive_lcell_comb \memwb_if.dmemload_o[14]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[14]~feeder_combout  = ramiframload_14

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_14),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[14]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.dmemload_o[14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N6
cycloneive_lcell_comb \memwb_if.dmemload_o[13]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[13]~feeder_combout  = ramiframload_13

	.dataa(gnd),
	.datab(ramiframload_13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[13]~feeder .lut_mask = 16'hCCCC;
defparam \memwb_if.dmemload_o[13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N18
cycloneive_lcell_comb \memwb_if.dmemload_o[10]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[10]~feeder_combout  = ramiframload_10

	.dataa(gnd),
	.datab(gnd),
	.datac(ramiframload_10),
	.datad(gnd),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[10]~feeder .lut_mask = 16'hF0F0;
defparam \memwb_if.dmemload_o[10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N18
cycloneive_lcell_comb \memwb_if.dmemload_o[9]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[9]~feeder_combout  = ramiframload_9

	.dataa(ramiframload_9),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[9]~feeder .lut_mask = 16'hAAAA;
defparam \memwb_if.dmemload_o[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N0
cycloneive_lcell_comb \memwb_if.dmemload_o[31]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[31]~feeder_combout  = ramiframload_31

	.dataa(ramiframload_31),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[31]~feeder .lut_mask = 16'hAAAA;
defparam \memwb_if.dmemload_o[31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N24
cycloneive_lcell_comb \memwb_if.dmemload_o[29]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[29]~feeder_combout  = ramiframload_29

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_29),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[29]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.dmemload_o[29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N6
cycloneive_lcell_comb \memwb_if.imm_o[13]~feeder (
// Equation(s):
// \memwb_if.imm_o[13]~feeder_combout  = exmem_ifimm_o_13

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifimm_o_13),
	.cin(gnd),
	.combout(\memwb_if.imm_o[13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.imm_o[13]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.imm_o[13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N20
cycloneive_lcell_comb \memwb_if.next_pc_o[30]~feeder (
// Equation(s):
// \memwb_if.next_pc_o[30]~feeder_combout  = exmem_ifnext_pc_o_30

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifnext_pc_o_30),
	.cin(gnd),
	.combout(\memwb_if.next_pc_o[30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.next_pc_o[30]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.next_pc_o[30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N18
cycloneive_lcell_comb \memwb_if.imm_o[14]~feeder (
// Equation(s):
// \memwb_if.imm_o[14]~feeder_combout  = exmem_ifimm_o_14

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifimm_o_14),
	.cin(gnd),
	.combout(\memwb_if.imm_o[14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.imm_o[14]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.imm_o[14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N18
cycloneive_lcell_comb \memwb_if.dmemload_o[27]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[27]~feeder_combout  = ramiframload_27

	.dataa(gnd),
	.datab(gnd),
	.datac(ramiframload_27),
	.datad(gnd),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[27]~feeder .lut_mask = 16'hF0F0;
defparam \memwb_if.dmemload_o[27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N22
cycloneive_lcell_comb \memwb_if.imm_o[11]~feeder (
// Equation(s):
// \memwb_if.imm_o[11]~feeder_combout  = exmem_ifimm_o_11

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifimm_o_11),
	.cin(gnd),
	.combout(\memwb_if.imm_o[11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.imm_o[11]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.imm_o[11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N2
cycloneive_lcell_comb \memwb_if.dmemload_o[25]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[25]~feeder_combout  = ramiframload_25

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_25),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[25]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.dmemload_o[25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N22
cycloneive_lcell_comb \memwb_if.next_pc_o[24]~feeder (
// Equation(s):
// \memwb_if.next_pc_o[24]~feeder_combout  = exmem_ifnext_pc_o_24

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifnext_pc_o_24),
	.cin(gnd),
	.combout(\memwb_if.next_pc_o[24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.next_pc_o[24]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.next_pc_o[24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N28
cycloneive_lcell_comb \memwb_if.imm_o[8]~feeder (
// Equation(s):
// \memwb_if.imm_o[8]~feeder_combout  = exmem_ifimm_o_8

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifimm_o_8),
	.cin(gnd),
	.combout(\memwb_if.imm_o[8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.imm_o[8]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.imm_o[8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N12
cycloneive_lcell_comb \memwb_if.dmemload_o[23]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[23]~feeder_combout  = ramiframload_23

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_23),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[23]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.dmemload_o[23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N28
cycloneive_lcell_comb \memwb_if.imm_o[7]~feeder (
// Equation(s):
// \memwb_if.imm_o[7]~feeder_combout  = exmem_ifimm_o_7

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifimm_o_7),
	.cin(gnd),
	.combout(\memwb_if.imm_o[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.imm_o[7]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.imm_o[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N16
cycloneive_lcell_comb \memwb_if.dmemload_o[21]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[21]~feeder_combout  = ramiframload_21

	.dataa(gnd),
	.datab(gnd),
	.datac(ramiframload_21),
	.datad(gnd),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[21]~feeder .lut_mask = 16'hF0F0;
defparam \memwb_if.dmemload_o[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N12
cycloneive_lcell_comb \memwb_if.imm_o[5]~feeder (
// Equation(s):
// \memwb_if.imm_o[5]~feeder_combout  = exmem_ifimm_o_5

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifimm_o_5),
	.cin(gnd),
	.combout(\memwb_if.imm_o[5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.imm_o[5]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.imm_o[5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N8
cycloneive_lcell_comb \memwb_if.next_pc_o[20]~feeder (
// Equation(s):
// \memwb_if.next_pc_o[20]~feeder_combout  = exmem_ifnext_pc_o_20

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifnext_pc_o_20),
	.cin(gnd),
	.combout(\memwb_if.next_pc_o[20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.next_pc_o[20]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.next_pc_o[20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N24
cycloneive_lcell_comb \memwb_if.imm_o[4]~feeder (
// Equation(s):
// \memwb_if.imm_o[4]~feeder_combout  = exmem_ifimm_o_4

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifimm_o_4),
	.cin(gnd),
	.combout(\memwb_if.imm_o[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.imm_o[4]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.imm_o[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N20
cycloneive_lcell_comb \memwb_if.next_pc_o[18]~feeder (
// Equation(s):
// \memwb_if.next_pc_o[18]~feeder_combout  = exmem_ifnext_pc_o_18

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifnext_pc_o_18),
	.cin(gnd),
	.combout(\memwb_if.next_pc_o[18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.next_pc_o[18]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.next_pc_o[18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N0
cycloneive_lcell_comb \memwb_if.imm_o[2]~feeder (
// Equation(s):
// \memwb_if.imm_o[2]~feeder_combout  = exmem_ifimm_o_2

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifimm_o_2),
	.cin(gnd),
	.combout(\memwb_if.imm_o[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.imm_o[2]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.imm_o[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N2
cycloneive_lcell_comb \memwb_if.dmemload_o[19]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[19]~feeder_combout  = ramiframload_19

	.dataa(gnd),
	.datab(gnd),
	.datac(ramiframload_19),
	.datad(gnd),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[19]~feeder .lut_mask = 16'hF0F0;
defparam \memwb_if.dmemload_o[19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N16
cycloneive_lcell_comb \memwb_if.next_pc_o[17]~feeder (
// Equation(s):
// \memwb_if.next_pc_o[17]~feeder_combout  = exmem_ifnext_pc_o_17

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(exmem_ifnext_pc_o_17),
	.cin(gnd),
	.combout(\memwb_if.next_pc_o[17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.next_pc_o[17]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.next_pc_o[17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N16
cycloneive_lcell_comb \memwb_if.dmemload_o[17]~feeder (
// Equation(s):
// \memwb_if.dmemload_o[17]~feeder_combout  = ramiframload_17

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramiframload_17),
	.cin(gnd),
	.combout(\memwb_if.dmemload_o[17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \memwb_if.dmemload_o[17]~feeder .lut_mask = 16'hFF00;
defparam \memwb_if.dmemload_o[17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module register_file (
	rwWB,
	rwWB1,
	rwWB2,
	rwWB3,
	memwb_ifregWEN_o,
	rwWB4,
	wdat,
	wdat1,
	wdat2,
	wdat3,
	wdat4,
	wdat5,
	wdat6,
	wdat7,
	wdat8,
	wdat9,
	wdat10,
	wdat11,
	wdat12,
	wdat13,
	wdat14,
	wdat15,
	wdat16,
	wdat17,
	wdat18,
	wdat19,
	wdat20,
	wdat21,
	wdat22,
	wdat23,
	wdat24,
	wdat25,
	wdat26,
	wdat27,
	wdat28,
	wdat29,
	wdat30,
	wdat31,
	ifid_ifinstr_o_17,
	ifid_ifinstr_o_16,
	ifid_ifinstr_o_19,
	ifid_ifinstr_o_18,
	ifid_ifinstr_o_22,
	ifid_ifinstr_o_21,
	ifid_ifinstr_o_24,
	ifid_ifinstr_o_23,
	Mux62,
	Mux621,
	Mux30,
	Mux301,
	Mux63,
	Mux631,
	Mux31,
	Mux311,
	Mux29,
	Mux291,
	Mux27,
	Mux271,
	Mux28,
	Mux281,
	Mux61,
	Mux611,
	Mux23,
	Mux231,
	Mux24,
	Mux241,
	Mux25,
	Mux251,
	Mux26,
	Mux261,
	Mux60,
	Mux601,
	Mux15,
	Mux151,
	Mux16,
	Mux161,
	Mux17,
	Mux171,
	Mux18,
	Mux181,
	Mux19,
	Mux191,
	Mux20,
	Mux201,
	Mux21,
	Mux211,
	Mux22,
	Mux221,
	Mux59,
	Mux591,
	Mux0,
	Mux01,
	Mux2,
	Mux210,
	Mux1,
	Mux11,
	Mux3,
	Mux32,
	Mux5,
	Mux51,
	Mux4,
	Mux41,
	Mux6,
	Mux64,
	Mux7,
	Mux71,
	Mux9,
	Mux91,
	Mux8,
	Mux81,
	Mux10,
	Mux101,
	Mux111,
	Mux112,
	Mux13,
	Mux131,
	Mux12,
	Mux121,
	Mux14,
	Mux141,
	Mux321,
	Mux322,
	Mux47,
	Mux471,
	Mux46,
	Mux461,
	Mux45,
	Mux451,
	Mux44,
	Mux441,
	Mux43,
	Mux431,
	Mux42,
	Mux421,
	Mux411,
	Mux412,
	Mux40,
	Mux401,
	Mux39,
	Mux391,
	Mux38,
	Mux381,
	Mux37,
	Mux371,
	Mux58,
	Mux581,
	Mux57,
	Mux571,
	Mux56,
	Mux561,
	Mux55,
	Mux551,
	Mux36,
	Mux361,
	Mux35,
	Mux351,
	Mux34,
	Mux341,
	Mux33,
	Mux331,
	Mux54,
	Mux541,
	Mux49,
	Mux491,
	Mux48,
	Mux481,
	Mux53,
	Mux531,
	Mux52,
	Mux521,
	Mux511,
	Mux512,
	Mux50,
	Mux501,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	rwWB;
input 	rwWB1;
input 	rwWB2;
input 	rwWB3;
input 	memwb_ifregWEN_o;
input 	rwWB4;
input 	wdat;
input 	wdat1;
input 	wdat2;
input 	wdat3;
input 	wdat4;
input 	wdat5;
input 	wdat6;
input 	wdat7;
input 	wdat8;
input 	wdat9;
input 	wdat10;
input 	wdat11;
input 	wdat12;
input 	wdat13;
input 	wdat14;
input 	wdat15;
input 	wdat16;
input 	wdat17;
input 	wdat18;
input 	wdat19;
input 	wdat20;
input 	wdat21;
input 	wdat22;
input 	wdat23;
input 	wdat24;
input 	wdat25;
input 	wdat26;
input 	wdat27;
input 	wdat28;
input 	wdat29;
input 	wdat30;
input 	wdat31;
input 	ifid_ifinstr_o_17;
input 	ifid_ifinstr_o_16;
input 	ifid_ifinstr_o_19;
input 	ifid_ifinstr_o_18;
input 	ifid_ifinstr_o_22;
input 	ifid_ifinstr_o_21;
input 	ifid_ifinstr_o_24;
input 	ifid_ifinstr_o_23;
output 	Mux62;
output 	Mux621;
output 	Mux30;
output 	Mux301;
output 	Mux63;
output 	Mux631;
output 	Mux31;
output 	Mux311;
output 	Mux29;
output 	Mux291;
output 	Mux27;
output 	Mux271;
output 	Mux28;
output 	Mux281;
output 	Mux61;
output 	Mux611;
output 	Mux23;
output 	Mux231;
output 	Mux24;
output 	Mux241;
output 	Mux25;
output 	Mux251;
output 	Mux26;
output 	Mux261;
output 	Mux60;
output 	Mux601;
output 	Mux15;
output 	Mux151;
output 	Mux16;
output 	Mux161;
output 	Mux17;
output 	Mux171;
output 	Mux18;
output 	Mux181;
output 	Mux19;
output 	Mux191;
output 	Mux20;
output 	Mux201;
output 	Mux21;
output 	Mux211;
output 	Mux22;
output 	Mux221;
output 	Mux59;
output 	Mux591;
output 	Mux0;
output 	Mux01;
output 	Mux2;
output 	Mux210;
output 	Mux1;
output 	Mux11;
output 	Mux3;
output 	Mux32;
output 	Mux5;
output 	Mux51;
output 	Mux4;
output 	Mux41;
output 	Mux6;
output 	Mux64;
output 	Mux7;
output 	Mux71;
output 	Mux9;
output 	Mux91;
output 	Mux8;
output 	Mux81;
output 	Mux10;
output 	Mux101;
output 	Mux111;
output 	Mux112;
output 	Mux13;
output 	Mux131;
output 	Mux12;
output 	Mux121;
output 	Mux14;
output 	Mux141;
output 	Mux321;
output 	Mux322;
output 	Mux47;
output 	Mux471;
output 	Mux46;
output 	Mux461;
output 	Mux45;
output 	Mux451;
output 	Mux44;
output 	Mux441;
output 	Mux43;
output 	Mux431;
output 	Mux42;
output 	Mux421;
output 	Mux411;
output 	Mux412;
output 	Mux40;
output 	Mux401;
output 	Mux39;
output 	Mux391;
output 	Mux38;
output 	Mux381;
output 	Mux37;
output 	Mux371;
output 	Mux58;
output 	Mux581;
output 	Mux57;
output 	Mux571;
output 	Mux56;
output 	Mux561;
output 	Mux55;
output 	Mux551;
output 	Mux36;
output 	Mux361;
output 	Mux35;
output 	Mux351;
output 	Mux34;
output 	Mux341;
output 	Mux33;
output 	Mux331;
output 	Mux54;
output 	Mux541;
output 	Mux49;
output 	Mux491;
output 	Mux48;
output 	Mux481;
output 	Mux53;
output 	Mux531;
output 	Mux52;
output 	Mux521;
output 	Mux511;
output 	Mux512;
output 	Mux50;
output 	Mux501;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Mux62~14_combout ;
wire \Reg[3][4]~q ;
wire \Reg[1][4]~q ;
wire \Mux27~14_combout ;
wire \Reg[1][3]~q ;
wire \Mux28~14_combout ;
wire \Mux61~2_combout ;
wire \Mux61~12_combout ;
wire \Mux24~4_combout ;
wire \Mux24~12_combout ;
wire \Reg[3][6]~q ;
wire \Mux25~14_combout ;
wire \Mux60~2_combout ;
wire \Mux15~2_combout ;
wire \Reg[28][16]~q ;
wire \Reg[8][15]~q ;
wire \Mux16~12_combout ;
wire \Reg[30][14]~q ;
wire \Mux17~4_combout ;
wire \Mux18~12_combout ;
wire \Reg[22][11]~q ;
wire \Mux20~4_combout ;
wire \Reg[3][9]~q ;
wire \Mux22~14_combout ;
wire \Mux59~12_combout ;
wire \Mux59~14_combout ;
wire \Reg[24][31]~q ;
wire \Mux0~4_combout ;
wire \Reg[8][31]~q ;
wire \Reg[20][29]~q ;
wire \Mux1~12_combout ;
wire \Reg[3][30]~q ;
wire \Mux1~14_combout ;
wire \Mux3~12_combout ;
wire \Reg[30][26]~q ;
wire \Reg[4][26]~q ;
wire \Reg[28][27]~q ;
wire \Reg[3][24]~q ;
wire \Reg[3][23]~q ;
wire \Reg[26][21]~q ;
wire \Reg[4][21]~q ;
wire \Mux10~12_combout ;
wire \Reg[4][20]~q ;
wire \Reg[3][20]~q ;
wire \Reg[1][20]~q ;
wire \Mux11~14_combout ;
wire \Mux13~4_combout ;
wire \Reg[28][19]~q ;
wire \Mux14~12_combout ;
wire \Mux32~2_combout ;
wire \Mux32~12_combout ;
wire \Mux32~14_combout ;
wire \Mux47~12_combout ;
wire \Mux46~14_combout ;
wire \Mux45~12_combout ;
wire \Mux45~14_combout ;
wire \Mux43~12_combout ;
wire \Mux43~14_combout ;
wire \Mux42~14_combout ;
wire \Mux40~4_combout ;
wire \Mux40~14_combout ;
wire \Mux39~14_combout ;
wire \Mux37~12_combout ;
wire \Mux58~2_combout ;
wire \Mux35~4_combout ;
wire \Mux35~12_combout ;
wire \Mux35~14_combout ;
wire \Mux33~4_combout ;
wire \Mux33~12_combout ;
wire \Mux49~12_combout ;
wire \Mux48~12_combout ;
wire \Mux53~2_combout ;
wire \Mux52~2_combout ;
wire \Mux51~12_combout ;
wire \Mux51~14_combout ;
wire \Reg[28][16]~feeder_combout ;
wire \Reg[30][14]~feeder_combout ;
wire \Reg[22][11]~feeder_combout ;
wire \Reg[20][29]~feeder_combout ;
wire \Reg[30][26]~feeder_combout ;
wire \Reg[28][27]~feeder_combout ;
wire \Reg[3][24]~feeder_combout ;
wire \Reg[3][23]~feeder_combout ;
wire \Reg[26][21]~feeder_combout ;
wire \Reg[28][19]~feeder_combout ;
wire \Reg[21][1]~feeder_combout ;
wire \Decoder0~0_combout ;
wire \Decoder0~1_combout ;
wire \Reg[21][1]~q ;
wire \Reg[29][1]~feeder_combout ;
wire \Decoder0~4_combout ;
wire \Reg[29][1]~q ;
wire \Decoder0~2_combout ;
wire \Reg[25][1]~q ;
wire \Decoder0~3_combout ;
wire \Reg[17][1]~q ;
wire \Mux62~0_combout ;
wire \Mux62~1_combout ;
wire \Decoder0~5_combout ;
wire \Decoder0~6_combout ;
wire \Reg[26][1]~q ;
wire \Decoder0~7_combout ;
wire \Reg[22][1]~q ;
wire \Decoder0~8_combout ;
wire \Reg[18][1]~q ;
wire \Mux62~2_combout ;
wire \Mux62~3_combout ;
wire \Decoder0~11_combout ;
wire \Reg[20][1]~q ;
wire \Decoder0~12_combout ;
wire \Reg[16][1]~q ;
wire \Mux62~4_combout ;
wire \Decoder0~13_combout ;
wire \Reg[28][1]~q ;
wire \Reg[24][1]~feeder_combout ;
wire \Decoder0~10_combout ;
wire \Reg[24][1]~q ;
wire \Mux62~5_combout ;
wire \Mux62~6_combout ;
wire \Decoder0~14_combout ;
wire \Reg[23][1]~q ;
wire \Decoder0~16_combout ;
wire \Reg[19][1]~q ;
wire \Decoder0~15_combout ;
wire \Reg[27][1]~q ;
wire \Mux62~7_combout ;
wire \Decoder0~17_combout ;
wire \Reg[31][1]~q ;
wire \Mux62~8_combout ;
wire \Decoder0~36_combout ;
wire \Reg[15][1]~q ;
wire \Decoder0~18_combout ;
wire \Decoder0~33_combout ;
wire \Reg[14][1]~q ;
wire \Decoder0~35_combout ;
wire \Reg[12][1]~q ;
wire \Decoder0~20_combout ;
wire \Decoder0~34_combout ;
wire \Reg[13][1]~q ;
wire \Mux62~17_combout ;
wire \Mux62~18_combout ;
wire \Decoder0~21_combout ;
wire \Reg[5][1]~q ;
wire \Mux62~10_combout ;
wire \Reg[7][1]~feeder_combout ;
wire \Decoder0~23_combout ;
wire \Reg[7][1]~q ;
wire \Reg[6][1]~feeder_combout ;
wire \Decoder0~19_combout ;
wire \Reg[6][1]~q ;
wire \Mux62~11_combout ;
wire \Reg[2][1]~feeder_combout ;
wire \Decoder0~26_combout ;
wire \Decoder0~32_combout ;
wire \Reg[2][1]~q ;
wire \Mux62~15_combout ;
wire \Decoder0~24_combout ;
wire \Decoder0~25_combout ;
wire \Reg[9][1]~q ;
wire \Decoder0~29_combout ;
wire \Reg[11][1]~q ;
wire \Decoder0~28_combout ;
wire \Reg[8][1]~q ;
wire \Decoder0~27_combout ;
wire \Reg[10][1]~q ;
wire \Mux62~12_combout ;
wire \Mux62~13_combout ;
wire \Mux62~16_combout ;
wire \Mux30~0_combout ;
wire \Mux30~1_combout ;
wire \Mux30~2_combout ;
wire \Decoder0~9_combout ;
wire \Reg[30][1]~q ;
wire \Mux30~3_combout ;
wire \Mux30~4_combout ;
wire \Mux30~5_combout ;
wire \Mux30~6_combout ;
wire \Mux30~7_combout ;
wire \Mux30~8_combout ;
wire \Mux30~10_combout ;
wire \Mux30~11_combout ;
wire \Decoder0~22_combout ;
wire \Reg[4][1]~q ;
wire \Mux30~12_combout ;
wire \Mux30~13_combout ;
wire \Decoder0~31_combout ;
wire \Reg[1][1]~q ;
wire \Decoder0~30_combout ;
wire \Reg[3][1]~q ;
wire \Mux30~14_combout ;
wire \Mux30~15_combout ;
wire \Mux30~16_combout ;
wire \Mux30~17_combout ;
wire \Mux30~18_combout ;
wire \Reg[25][0]~feeder_combout ;
wire \Reg[25][0]~q ;
wire \Reg[29][0]~feeder_combout ;
wire \Reg[29][0]~q ;
wire \Reg[21][0]~feeder_combout ;
wire \Reg[21][0]~q ;
wire \Reg[17][0]~feeder_combout ;
wire \Reg[17][0]~q ;
wire \Mux63~0_combout ;
wire \Mux63~1_combout ;
wire \Reg[19][0]~q ;
wire \Reg[23][0]~q ;
wire \Mux63~7_combout ;
wire \Reg[27][0]~q ;
wire \Reg[31][0]~q ;
wire \Mux63~8_combout ;
wire \Reg[28][0]~feeder_combout ;
wire \Reg[28][0]~q ;
wire \Reg[24][0]~q ;
wire \Reg[16][0]~feeder_combout ;
wire \Reg[16][0]~q ;
wire \Mux63~4_combout ;
wire \Mux63~5_combout ;
wire \Reg[30][0]~feeder_combout ;
wire \Reg[30][0]~q ;
wire \Reg[18][0]~q ;
wire \Reg[26][0]~q ;
wire \Mux63~2_combout ;
wire \Reg[22][0]~feeder_combout ;
wire \Reg[22][0]~q ;
wire \Mux63~3_combout ;
wire \Mux63~6_combout ;
wire \Reg[15][0]~feeder_combout ;
wire \Reg[15][0]~q ;
wire \Reg[14][0]~feeder_combout ;
wire \Reg[14][0]~q ;
wire \Reg[13][0]~q ;
wire \Mux63~17_combout ;
wire \Mux63~18_combout ;
wire \Reg[1][0]~q ;
wire \Reg[3][0]~feeder_combout ;
wire \Reg[3][0]~q ;
wire \Mux63~14_combout ;
wire \Reg[2][0]~feeder_combout ;
wire \Reg[2][0]~q ;
wire \Mux63~15_combout ;
wire \Reg[4][0]~q ;
wire \Reg[5][0]~q ;
wire \Mux63~12_combout ;
wire \Reg[7][0]~q ;
wire \Reg[6][0]~q ;
wire \Mux63~13_combout ;
wire \Mux63~16_combout ;
wire \Reg[11][0]~q ;
wire \Reg[10][0]~q ;
wire \Reg[8][0]~q ;
wire \Mux63~10_combout ;
wire \Reg[9][0]~q ;
wire \Mux63~11_combout ;
wire \Mux31~0_combout ;
wire \Mux31~1_combout ;
wire \Mux31~7_combout ;
wire \Mux31~8_combout ;
wire \Reg[20][0]~feeder_combout ;
wire \Reg[20][0]~q ;
wire \Mux31~4_combout ;
wire \Mux31~5_combout ;
wire \Mux31~2_combout ;
wire \Mux31~3_combout ;
wire \Mux31~6_combout ;
wire \Reg[12][0]~q ;
wire \Mux31~17_combout ;
wire \Mux31~18_combout ;
wire \Mux31~14_combout ;
wire \Mux31~15_combout ;
wire \Mux31~12_combout ;
wire \Mux31~13_combout ;
wire \Mux31~16_combout ;
wire \Mux31~10_combout ;
wire \Mux31~11_combout ;
wire \Reg[21][2]~feeder_combout ;
wire \Reg[21][2]~q ;
wire \Reg[29][2]~feeder_combout ;
wire \Reg[29][2]~q ;
wire \Reg[17][2]~feeder_combout ;
wire \Reg[17][2]~q ;
wire \Mux29~0_combout ;
wire \Mux29~1_combout ;
wire \Reg[27][2]~q ;
wire \Reg[19][2]~q ;
wire \Mux29~7_combout ;
wire \Reg[31][2]~q ;
wire \Reg[23][2]~feeder_combout ;
wire \Reg[23][2]~q ;
wire \Mux29~8_combout ;
wire \Reg[26][2]~q ;
wire \Reg[18][2]~q ;
wire \Reg[22][2]~q ;
wire \Mux29~2_combout ;
wire \Mux29~3_combout ;
wire \Reg[24][2]~q ;
wire \Reg[28][2]~q ;
wire \Reg[16][2]~q ;
wire \Reg[20][2]~q ;
wire \Mux29~4_combout ;
wire \Mux29~5_combout ;
wire \Mux29~6_combout ;
wire \Reg[4][2]~q ;
wire \Reg[5][2]~q ;
wire \Mux29~10_combout ;
wire \Reg[6][2]~feeder_combout ;
wire \Reg[6][2]~q ;
wire \Reg[7][2]~q ;
wire \Mux29~11_combout ;
wire \Reg[12][2]~q ;
wire \Reg[13][2]~q ;
wire \Mux29~17_combout ;
wire \Reg[15][2]~q ;
wire \Reg[14][2]~q ;
wire \Mux29~18_combout ;
wire \Reg[2][2]~q ;
wire \Reg[3][2]~q ;
wire \Mux29~14_combout ;
wire \Mux29~15_combout ;
wire \Reg[9][2]~q ;
wire \Reg[11][2]~q ;
wire \Reg[10][2]~q ;
wire \Reg[8][2]~q ;
wire \Mux29~12_combout ;
wire \Mux29~13_combout ;
wire \Mux29~16_combout ;
wire \Reg[29][4]~feeder_combout ;
wire \Reg[29][4]~q ;
wire \Reg[17][4]~q ;
wire \Reg[25][4]~feeder_combout ;
wire \Reg[25][4]~q ;
wire \Mux27~0_combout ;
wire \Reg[21][4]~q ;
wire \Mux27~1_combout ;
wire \Reg[16][4]~q ;
wire \Reg[20][4]~feeder_combout ;
wire \Reg[20][4]~q ;
wire \Mux27~4_combout ;
wire \Reg[24][4]~q ;
wire \Reg[28][4]~q ;
wire \Mux27~5_combout ;
wire \Reg[22][4]~feeder_combout ;
wire \Reg[22][4]~q ;
wire \Mux27~2_combout ;
wire \Reg[30][4]~q ;
wire \Mux27~3_combout ;
wire \Mux27~6_combout ;
wire \Reg[23][4]~feeder_combout ;
wire \Reg[23][4]~q ;
wire \Reg[27][4]~q ;
wire \Reg[19][4]~q ;
wire \Mux27~7_combout ;
wire \Reg[31][4]~q ;
wire \Mux27~8_combout ;
wire \Reg[2][4]~q ;
wire \Mux27~15_combout ;
wire \Reg[10][4]~q ;
wire \Reg[8][4]~q ;
wire \Mux27~12_combout ;
wire \Reg[11][4]~q ;
wire \Reg[9][4]~q ;
wire \Mux27~13_combout ;
wire \Mux27~16_combout ;
wire \Reg[5][4]~q ;
wire \Reg[4][4]~q ;
wire \Mux27~10_combout ;
wire \Reg[6][4]~q ;
wire \Reg[7][4]~q ;
wire \Mux27~11_combout ;
wire \Reg[14][4]~q ;
wire \Reg[15][4]~q ;
wire \Reg[12][4]~q ;
wire \Reg[13][4]~q ;
wire \Mux27~17_combout ;
wire \Mux27~18_combout ;
wire \Reg[19][3]~q ;
wire \Reg[23][3]~q ;
wire \Mux28~7_combout ;
wire \Reg[31][3]~q ;
wire \Reg[27][3]~feeder_combout ;
wire \Reg[27][3]~q ;
wire \Mux28~8_combout ;
wire \Reg[25][3]~q ;
wire \Reg[29][3]~feeder_combout ;
wire \Reg[29][3]~q ;
wire \Reg[21][3]~q ;
wire \Reg[17][3]~q ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \Reg[30][3]~feeder_combout ;
wire \Reg[30][3]~q ;
wire \Reg[22][3]~q ;
wire \Reg[26][3]~feeder_combout ;
wire \Reg[26][3]~q ;
wire \Reg[18][3]~feeder_combout ;
wire \Reg[18][3]~q ;
wire \Mux28~2_combout ;
wire \Mux28~3_combout ;
wire \Reg[16][3]~q ;
wire \Reg[24][3]~feeder_combout ;
wire \Reg[24][3]~q ;
wire \Mux28~4_combout ;
wire \Reg[20][3]~q ;
wire \Reg[28][3]~q ;
wire \Mux28~5_combout ;
wire \Mux28~6_combout ;
wire \Reg[5][3]~q ;
wire \Reg[4][3]~q ;
wire \Mux28~12_combout ;
wire \Reg[7][3]~q ;
wire \Mux28~13_combout ;
wire \Reg[2][3]~q ;
wire \Mux28~15_combout ;
wire \Mux28~16_combout ;
wire \Reg[13][3]~q ;
wire \Reg[12][3]~q ;
wire \Mux28~17_combout ;
wire \Reg[14][3]~q ;
wire \Reg[15][3]~q ;
wire \Mux28~18_combout ;
wire \Reg[11][3]~q ;
wire \Reg[9][3]~q ;
wire \Reg[10][3]~q ;
wire \Mux28~10_combout ;
wire \Mux28~11_combout ;
wire \Mux61~4_combout ;
wire \Mux61~5_combout ;
wire \Reg[30][2]~q ;
wire \Mux61~3_combout ;
wire \Mux61~6_combout ;
wire \Mux61~7_combout ;
wire \Mux61~8_combout ;
wire \Mux61~0_combout ;
wire \Reg[25][2]~feeder_combout ;
wire \Reg[25][2]~q ;
wire \Mux61~1_combout ;
wire \Mux61~10_combout ;
wire \Mux61~11_combout ;
wire \Mux61~17_combout ;
wire \Mux61~18_combout ;
wire \Reg[1][2]~feeder_combout ;
wire \Reg[1][2]~q ;
wire \Mux61~14_combout ;
wire \Mux61~15_combout ;
wire \Mux61~13_combout ;
wire \Mux61~16_combout ;
wire \Reg[30][8]~q ;
wire \Reg[26][8]~q ;
wire \Reg[18][8]~feeder_combout ;
wire \Reg[18][8]~q ;
wire \Reg[22][8]~q ;
wire \Mux23~2_combout ;
wire \Mux23~3_combout ;
wire \Reg[24][8]~q ;
wire \Reg[16][8]~q ;
wire \Reg[20][8]~feeder_combout ;
wire \Reg[20][8]~q ;
wire \Mux23~4_combout ;
wire \Mux23~5_combout ;
wire \Mux23~6_combout ;
wire \Reg[23][8]~q ;
wire \Reg[31][8]~q ;
wire \Reg[27][8]~q ;
wire \Mux23~7_combout ;
wire \Mux23~8_combout ;
wire \Reg[21][8]~feeder_combout ;
wire \Reg[21][8]~q ;
wire \Reg[25][8]~feeder_combout ;
wire \Reg[25][8]~q ;
wire \Reg[17][8]~feeder_combout ;
wire \Reg[17][8]~q ;
wire \Mux23~0_combout ;
wire \Reg[29][8]~feeder_combout ;
wire \Reg[29][8]~q ;
wire \Mux23~1_combout ;
wire \Reg[7][8]~q ;
wire \Reg[6][8]~q ;
wire \Reg[5][8]~q ;
wire \Reg[4][8]~q ;
wire \Mux23~10_combout ;
wire \Mux23~11_combout ;
wire \Reg[12][8]~q ;
wire \Reg[13][8]~feeder_combout ;
wire \Reg[13][8]~q ;
wire \Mux23~17_combout ;
wire \Reg[15][8]~q ;
wire \Reg[14][8]~q ;
wire \Mux23~18_combout ;
wire \Reg[11][8]~q ;
wire \Reg[10][8]~q ;
wire \Reg[8][8]~q ;
wire \Mux23~12_combout ;
wire \Mux23~13_combout ;
wire \Reg[2][8]~q ;
wire \Reg[1][8]~q ;
wire \Reg[3][8]~q ;
wire \Mux23~14_combout ;
wire \Mux23~15_combout ;
wire \Mux23~16_combout ;
wire \Reg[31][7]~feeder_combout ;
wire \Reg[31][7]~q ;
wire \Reg[19][7]~q ;
wire \Reg[23][7]~q ;
wire \Mux24~7_combout ;
wire \Reg[27][7]~feeder_combout ;
wire \Reg[27][7]~q ;
wire \Mux24~8_combout ;
wire \Reg[25][7]~q ;
wire \Reg[17][7]~q ;
wire \Mux24~0_combout ;
wire \Reg[29][7]~feeder_combout ;
wire \Reg[29][7]~q ;
wire \Mux24~1_combout ;
wire \Reg[28][7]~q ;
wire \Reg[20][7]~q ;
wire \Mux24~5_combout ;
wire \Reg[18][7]~q ;
wire \Reg[26][7]~q ;
wire \Mux24~2_combout ;
wire \Reg[22][7]~q ;
wire \Mux24~3_combout ;
wire \Mux24~6_combout ;
wire \Reg[2][7]~q ;
wire \Reg[1][7]~q ;
wire \Reg[3][7]~q ;
wire \Mux24~14_combout ;
wire \Mux24~15_combout ;
wire \Reg[6][7]~q ;
wire \Reg[7][7]~q ;
wire \Mux24~13_combout ;
wire \Mux24~16_combout ;
wire \Reg[14][7]~q ;
wire \Reg[15][7]~q ;
wire \Reg[13][7]~q ;
wire \Mux24~17_combout ;
wire \Mux24~18_combout ;
wire \Reg[9][7]~feeder_combout ;
wire \Reg[9][7]~q ;
wire \Reg[11][7]~feeder_combout ;
wire \Reg[11][7]~q ;
wire \Reg[10][7]~q ;
wire \Mux24~10_combout ;
wire \Mux24~11_combout ;
wire \Reg[24][6]~feeder_combout ;
wire \Reg[24][6]~q ;
wire \Reg[28][6]~q ;
wire \Reg[20][6]~q ;
wire \Reg[16][6]~q ;
wire \Mux25~4_combout ;
wire \Mux25~5_combout ;
wire \Reg[26][6]~q ;
wire \Reg[18][6]~q ;
wire \Reg[22][6]~feeder_combout ;
wire \Reg[22][6]~q ;
wire \Mux25~2_combout ;
wire \Mux25~3_combout ;
wire \Mux25~6_combout ;
wire \Reg[21][6]~feeder_combout ;
wire \Reg[21][6]~q ;
wire \Reg[25][6]~feeder_combout ;
wire \Reg[25][6]~q ;
wire \Mux25~0_combout ;
wire \Reg[29][6]~feeder_combout ;
wire \Reg[29][6]~q ;
wire \Mux25~1_combout ;
wire \Reg[23][6]~q ;
wire \Reg[19][6]~q ;
wire \Reg[27][6]~q ;
wire \Mux25~7_combout ;
wire \Reg[31][6]~q ;
wire \Mux25~8_combout ;
wire \Reg[14][6]~q ;
wire \Reg[15][6]~q ;
wire \Reg[13][6]~q ;
wire \Reg[12][6]~q ;
wire \Mux25~17_combout ;
wire \Mux25~18_combout ;
wire \Reg[5][6]~q ;
wire \Reg[4][6]~q ;
wire \Mux25~10_combout ;
wire \Reg[6][6]~q ;
wire \Reg[7][6]~q ;
wire \Mux25~11_combout ;
wire \Reg[2][6]~q ;
wire \Mux25~15_combout ;
wire \Reg[9][6]~q ;
wire \Reg[11][6]~q ;
wire \Reg[8][6]~q ;
wire \Reg[10][6]~q ;
wire \Mux25~12_combout ;
wire \Mux25~13_combout ;
wire \Mux25~16_combout ;
wire \Reg[27][5]~feeder_combout ;
wire \Reg[27][5]~q ;
wire \Reg[31][5]~q ;
wire \Reg[23][5]~q ;
wire \Mux26~7_combout ;
wire \Mux26~8_combout ;
wire \Reg[21][5]~feeder_combout ;
wire \Reg[21][5]~q ;
wire \Reg[17][5]~q ;
wire \Mux26~0_combout ;
wire \Reg[29][5]~q ;
wire \Reg[25][5]~q ;
wire \Mux26~1_combout ;
wire \Reg[16][5]~q ;
wire \Reg[24][5]~q ;
wire \Mux26~4_combout ;
wire \Reg[28][5]~q ;
wire \Reg[20][5]~q ;
wire \Mux26~5_combout ;
wire \Reg[18][5]~q ;
wire \Reg[26][5]~feeder_combout ;
wire \Reg[26][5]~q ;
wire \Mux26~2_combout ;
wire \Reg[22][5]~q ;
wire \Reg[30][5]~feeder_combout ;
wire \Reg[30][5]~q ;
wire \Mux26~3_combout ;
wire \Mux26~6_combout ;
wire \Reg[7][5]~q ;
wire \Reg[4][5]~q ;
wire \Reg[5][5]~q ;
wire \Mux26~12_combout ;
wire \Mux26~13_combout ;
wire \Reg[2][5]~q ;
wire \Reg[1][5]~q ;
wire \Reg[3][5]~feeder_combout ;
wire \Reg[3][5]~q ;
wire \Mux26~14_combout ;
wire \Mux26~15_combout ;
wire \Mux26~16_combout ;
wire \Reg[10][5]~q ;
wire \Mux26~10_combout ;
wire \Reg[11][5]~q ;
wire \Reg[9][5]~feeder_combout ;
wire \Reg[9][5]~q ;
wire \Mux26~11_combout ;
wire \Reg[15][5]~q ;
wire \Reg[14][5]~q ;
wire \Reg[13][5]~feeder_combout ;
wire \Reg[13][5]~q ;
wire \Mux26~17_combout ;
wire \Mux26~18_combout ;
wire \Mux60~7_combout ;
wire \Mux60~8_combout ;
wire \Mux60~0_combout ;
wire \Mux60~1_combout ;
wire \Mux60~3_combout ;
wire \Mux60~4_combout ;
wire \Mux60~5_combout ;
wire \Mux60~6_combout ;
wire \Reg[6][3]~feeder_combout ;
wire \Reg[6][3]~q ;
wire \Mux60~10_combout ;
wire \Mux60~11_combout ;
wire \Mux60~17_combout ;
wire \Mux60~18_combout ;
wire \Reg[8][3]~q ;
wire \Mux60~12_combout ;
wire \Mux60~13_combout ;
wire \Reg[3][3]~q ;
wire \Mux60~14_combout ;
wire \Mux60~15_combout ;
wire \Mux60~16_combout ;
wire \Reg[31][16]~q ;
wire \Reg[27][16]~q ;
wire \Reg[19][16]~q ;
wire \Mux15~7_combout ;
wire \Reg[23][16]~q ;
wire \Mux15~8_combout ;
wire \Reg[17][16]~q ;
wire \Reg[25][16]~feeder_combout ;
wire \Reg[25][16]~q ;
wire \Mux15~0_combout ;
wire \Reg[29][16]~feeder_combout ;
wire \Reg[29][16]~q ;
wire \Reg[21][16]~q ;
wire \Mux15~1_combout ;
wire \Reg[24][16]~q ;
wire \Reg[16][16]~q ;
wire \Mux15~4_combout ;
wire \Mux15~5_combout ;
wire \Reg[30][16]~q ;
wire \Reg[26][16]~q ;
wire \Mux15~3_combout ;
wire \Mux15~6_combout ;
wire \Reg[15][16]~q ;
wire \Reg[14][16]~q ;
wire \Reg[13][16]~q ;
wire \Reg[12][16]~q ;
wire \Mux15~17_combout ;
wire \Mux15~18_combout ;
wire \Reg[7][16]~q ;
wire \Reg[6][16]~q ;
wire \Reg[5][16]~q ;
wire \Reg[4][16]~q ;
wire \Mux15~10_combout ;
wire \Mux15~11_combout ;
wire \Reg[1][16]~q ;
wire \Reg[3][16]~q ;
wire \Mux15~14_combout ;
wire \Reg[2][16]~feeder_combout ;
wire \Reg[2][16]~q ;
wire \Mux15~15_combout ;
wire \Reg[9][16]~q ;
wire \Reg[11][16]~q ;
wire \Reg[8][16]~q ;
wire \Reg[10][16]~q ;
wire \Mux15~12_combout ;
wire \Mux15~13_combout ;
wire \Mux15~16_combout ;
wire \Reg[25][15]~feeder_combout ;
wire \Reg[25][15]~q ;
wire \Reg[29][15]~q ;
wire \Reg[21][15]~q ;
wire \Reg[17][15]~q ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \Reg[31][15]~feeder_combout ;
wire \Reg[31][15]~q ;
wire \Reg[27][15]~q ;
wire \Reg[23][15]~q ;
wire \Reg[19][15]~q ;
wire \Mux16~7_combout ;
wire \Mux16~8_combout ;
wire \Reg[26][15]~q ;
wire \Mux16~2_combout ;
wire \Reg[30][15]~q ;
wire \Reg[22][15]~feeder_combout ;
wire \Reg[22][15]~q ;
wire \Mux16~3_combout ;
wire \Reg[20][15]~q ;
wire \Reg[28][15]~q ;
wire \Reg[16][15]~q ;
wire \Reg[24][15]~q ;
wire \Mux16~4_combout ;
wire \Mux16~5_combout ;
wire \Mux16~6_combout ;
wire \Reg[3][15]~q ;
wire \Reg[1][15]~q ;
wire \Mux16~14_combout ;
wire \Reg[2][15]~feeder_combout ;
wire \Reg[2][15]~q ;
wire \Mux16~15_combout ;
wire \Reg[6][15]~q ;
wire \Reg[7][15]~q ;
wire \Mux16~13_combout ;
wire \Mux16~16_combout ;
wire \Reg[12][15]~q ;
wire \Reg[13][15]~q ;
wire \Mux16~17_combout ;
wire \Reg[14][15]~q ;
wire \Reg[15][15]~q ;
wire \Mux16~18_combout ;
wire \Reg[9][15]~q ;
wire \Reg[11][15]~feeder_combout ;
wire \Reg[11][15]~q ;
wire \Reg[10][15]~q ;
wire \Mux16~10_combout ;
wire \Mux16~11_combout ;
wire \Reg[21][14]~feeder_combout ;
wire \Reg[21][14]~q ;
wire \Reg[29][14]~q ;
wire \Reg[17][14]~feeder_combout ;
wire \Reg[17][14]~q ;
wire \Reg[25][14]~feeder_combout ;
wire \Reg[25][14]~q ;
wire \Mux17~0_combout ;
wire \Mux17~1_combout ;
wire \Reg[28][14]~q ;
wire \Reg[24][14]~feeder_combout ;
wire \Reg[24][14]~q ;
wire \Mux17~5_combout ;
wire \Reg[26][14]~q ;
wire \Reg[18][14]~q ;
wire \Reg[22][14]~feeder_combout ;
wire \Reg[22][14]~q ;
wire \Mux17~2_combout ;
wire \Mux17~3_combout ;
wire \Mux17~6_combout ;
wire \Reg[31][14]~q ;
wire \Reg[23][14]~q ;
wire \Reg[19][14]~q ;
wire \Reg[27][14]~feeder_combout ;
wire \Reg[27][14]~q ;
wire \Mux17~7_combout ;
wire \Mux17~8_combout ;
wire \Reg[15][14]~q ;
wire \Reg[14][14]~q ;
wire \Reg[13][14]~q ;
wire \Reg[12][14]~q ;
wire \Mux17~17_combout ;
wire \Mux17~18_combout ;
wire \Reg[7][14]~q ;
wire \Reg[6][14]~q ;
wire \Reg[5][14]~q ;
wire \Reg[4][14]~q ;
wire \Mux17~10_combout ;
wire \Mux17~11_combout ;
wire \Reg[8][14]~q ;
wire \Reg[10][14]~q ;
wire \Mux17~12_combout ;
wire \Reg[11][14]~q ;
wire \Reg[9][14]~q ;
wire \Mux17~13_combout ;
wire \Reg[2][14]~feeder_combout ;
wire \Reg[2][14]~q ;
wire \Reg[3][14]~q ;
wire \Reg[1][14]~q ;
wire \Mux17~14_combout ;
wire \Mux17~15_combout ;
wire \Mux17~16_combout ;
wire \Reg[19][13]~q ;
wire \Reg[23][13]~q ;
wire \Mux18~7_combout ;
wire \Reg[27][13]~feeder_combout ;
wire \Reg[27][13]~q ;
wire \Reg[31][13]~q ;
wire \Mux18~8_combout ;
wire \Reg[21][13]~feeder_combout ;
wire \Reg[21][13]~q ;
wire \Reg[17][13]~q ;
wire \Mux18~0_combout ;
wire \Reg[29][13]~feeder_combout ;
wire \Reg[29][13]~q ;
wire \Reg[25][13]~feeder_combout ;
wire \Reg[25][13]~q ;
wire \Mux18~1_combout ;
wire \Reg[16][13]~feeder_combout ;
wire \Reg[16][13]~q ;
wire \Reg[24][13]~q ;
wire \Mux18~4_combout ;
wire \Reg[20][13]~feeder_combout ;
wire \Reg[20][13]~q ;
wire \Mux18~5_combout ;
wire \Reg[30][13]~feeder_combout ;
wire \Reg[30][13]~q ;
wire \Reg[26][13]~q ;
wire \Reg[18][13]~q ;
wire \Mux18~2_combout ;
wire \Mux18~3_combout ;
wire \Mux18~6_combout ;
wire \Reg[3][13]~q ;
wire \Reg[1][13]~q ;
wire \Mux18~14_combout ;
wire \Reg[2][13]~q ;
wire \Mux18~15_combout ;
wire \Reg[7][13]~q ;
wire \Reg[6][13]~q ;
wire \Mux18~13_combout ;
wire \Mux18~16_combout ;
wire \Reg[14][13]~q ;
wire \Reg[15][13]~feeder_combout ;
wire \Reg[15][13]~q ;
wire \Reg[13][13]~q ;
wire \Reg[12][13]~q ;
wire \Mux18~17_combout ;
wire \Mux18~18_combout ;
wire \Reg[10][13]~q ;
wire \Reg[8][13]~q ;
wire \Mux18~10_combout ;
wire \Reg[9][13]~q ;
wire \Reg[11][13]~q ;
wire \Mux18~11_combout ;
wire \Reg[25][12]~feeder_combout ;
wire \Reg[25][12]~q ;
wire \Reg[17][12]~q ;
wire \Mux19~0_combout ;
wire \Reg[29][12]~q ;
wire \Reg[21][12]~q ;
wire \Mux19~1_combout ;
wire \Reg[31][12]~q ;
wire \Reg[23][12]~q ;
wire \Reg[19][12]~q ;
wire \Reg[27][12]~feeder_combout ;
wire \Reg[27][12]~q ;
wire \Mux19~7_combout ;
wire \Mux19~8_combout ;
wire \Reg[22][12]~q ;
wire \Mux19~2_combout ;
wire \Reg[30][12]~q ;
wire \Reg[26][12]~feeder_combout ;
wire \Reg[26][12]~q ;
wire \Mux19~3_combout ;
wire \Reg[20][12]~q ;
wire \Reg[16][12]~q ;
wire \Mux19~4_combout ;
wire \Reg[28][12]~q ;
wire \Mux19~5_combout ;
wire \Mux19~6_combout ;
wire \Reg[15][12]~feeder_combout ;
wire \Reg[15][12]~q ;
wire \Reg[14][12]~q ;
wire \Reg[13][12]~q ;
wire \Reg[12][12]~q ;
wire \Mux19~17_combout ;
wire \Mux19~18_combout ;
wire \Reg[5][12]~q ;
wire \Reg[4][12]~q ;
wire \Mux19~10_combout ;
wire \Reg[6][12]~q ;
wire \Reg[7][12]~q ;
wire \Mux19~11_combout ;
wire \Reg[9][12]~q ;
wire \Reg[11][12]~q ;
wire \Reg[8][12]~q ;
wire \Reg[10][12]~q ;
wire \Mux19~12_combout ;
wire \Mux19~13_combout ;
wire \Reg[2][12]~q ;
wire \Reg[3][12]~q ;
wire \Reg[1][12]~q ;
wire \Mux19~14_combout ;
wire \Mux19~15_combout ;
wire \Mux19~16_combout ;
wire \Reg[20][11]~feeder_combout ;
wire \Reg[20][11]~q ;
wire \Reg[28][11]~q ;
wire \Mux20~5_combout ;
wire \Reg[18][11]~q ;
wire \Reg[26][11]~q ;
wire \Mux20~2_combout ;
wire \Reg[30][11]~feeder_combout ;
wire \Reg[30][11]~q ;
wire \Mux20~3_combout ;
wire \Mux20~6_combout ;
wire \Reg[29][11]~q ;
wire \Reg[17][11]~q ;
wire \Reg[21][11]~feeder_combout ;
wire \Reg[21][11]~q ;
wire \Mux20~0_combout ;
wire \Reg[25][11]~feeder_combout ;
wire \Reg[25][11]~q ;
wire \Mux20~1_combout ;
wire \Reg[31][11]~q ;
wire \Reg[23][11]~feeder_combout ;
wire \Reg[23][11]~q ;
wire \Reg[19][11]~feeder_combout ;
wire \Reg[19][11]~q ;
wire \Mux20~7_combout ;
wire \Reg[27][11]~q ;
wire \Mux20~8_combout ;
wire \Reg[13][11]~q ;
wire \Mux20~17_combout ;
wire \Reg[15][11]~feeder_combout ;
wire \Reg[15][11]~q ;
wire \Reg[14][11]~q ;
wire \Mux20~18_combout ;
wire \Reg[9][11]~feeder_combout ;
wire \Reg[9][11]~q ;
wire \Reg[11][11]~q ;
wire \Reg[10][11]~q ;
wire \Mux20~10_combout ;
wire \Mux20~11_combout ;
wire \Reg[4][11]~q ;
wire \Reg[5][11]~q ;
wire \Mux20~12_combout ;
wire \Reg[7][11]~q ;
wire \Reg[6][11]~q ;
wire \Mux20~13_combout ;
wire \Reg[2][11]~q ;
wire \Reg[1][11]~q ;
wire \Reg[3][11]~q ;
wire \Mux20~14_combout ;
wire \Mux20~15_combout ;
wire \Mux20~16_combout ;
wire \Reg[21][10]~feeder_combout ;
wire \Reg[21][10]~q ;
wire \Reg[29][10]~feeder_combout ;
wire \Reg[29][10]~q ;
wire \Reg[17][10]~q ;
wire \Reg[25][10]~feeder_combout ;
wire \Reg[25][10]~q ;
wire \Mux21~0_combout ;
wire \Mux21~1_combout ;
wire \Reg[26][10]~q ;
wire \Reg[18][10]~q ;
wire \Reg[22][10]~q ;
wire \Mux21~2_combout ;
wire \Mux21~3_combout ;
wire \Reg[20][10]~q ;
wire \Reg[16][10]~feeder_combout ;
wire \Reg[16][10]~q ;
wire \Mux21~4_combout ;
wire \Reg[28][10]~q ;
wire \Reg[24][10]~feeder_combout ;
wire \Reg[24][10]~q ;
wire \Mux21~5_combout ;
wire \Mux21~6_combout ;
wire \Reg[27][10]~q ;
wire \Reg[19][10]~q ;
wire \Mux21~7_combout ;
wire \Reg[23][10]~q ;
wire \Reg[31][10]~q ;
wire \Mux21~8_combout ;
wire \Reg[7][10]~q ;
wire \Reg[5][10]~q ;
wire \Reg[4][10]~q ;
wire \Mux21~10_combout ;
wire \Reg[6][10]~q ;
wire \Mux21~11_combout ;
wire \Reg[13][10]~q ;
wire \Mux21~17_combout ;
wire \Reg[14][10]~q ;
wire \Reg[15][10]~q ;
wire \Mux21~18_combout ;
wire \Reg[2][10]~q ;
wire \Reg[3][10]~q ;
wire \Reg[1][10]~q ;
wire \Mux21~14_combout ;
wire \Mux21~15_combout ;
wire \Reg[11][10]~q ;
wire \Reg[8][10]~q ;
wire \Reg[10][10]~q ;
wire \Mux21~12_combout ;
wire \Mux21~13_combout ;
wire \Mux21~16_combout ;
wire \Reg[25][9]~q ;
wire \Reg[29][9]~q ;
wire \Reg[21][9]~q ;
wire \Reg[17][9]~q ;
wire \Mux22~0_combout ;
wire \Mux22~1_combout ;
wire \Reg[30][9]~q ;
wire \Reg[18][9]~q ;
wire \Reg[26][9]~feeder_combout ;
wire \Reg[26][9]~q ;
wire \Mux22~2_combout ;
wire \Mux22~3_combout ;
wire \Reg[20][9]~feeder_combout ;
wire \Reg[20][9]~q ;
wire \Reg[24][9]~q ;
wire \Mux22~4_combout ;
wire \Mux22~5_combout ;
wire \Mux22~6_combout ;
wire \Reg[31][9]~feeder_combout ;
wire \Reg[31][9]~q ;
wire \Reg[27][9]~q ;
wire \Reg[19][9]~q ;
wire \Reg[23][9]~feeder_combout ;
wire \Reg[23][9]~q ;
wire \Mux22~7_combout ;
wire \Mux22~8_combout ;
wire \Reg[14][9]~q ;
wire \Reg[15][9]~feeder_combout ;
wire \Reg[15][9]~q ;
wire \Reg[13][9]~q ;
wire \Reg[12][9]~q ;
wire \Mux22~17_combout ;
wire \Mux22~18_combout ;
wire \Reg[11][9]~q ;
wire \Reg[10][9]~q ;
wire \Reg[8][9]~q ;
wire \Mux22~10_combout ;
wire \Reg[9][9]~q ;
wire \Mux22~11_combout ;
wire \Reg[6][9]~q ;
wire \Reg[7][9]~q ;
wire \Reg[4][9]~q ;
wire \Reg[5][9]~q ;
wire \Mux22~12_combout ;
wire \Mux22~13_combout ;
wire \Reg[2][9]~feeder_combout ;
wire \Reg[2][9]~q ;
wire \Mux22~15_combout ;
wire \Mux22~16_combout ;
wire \Mux59~0_combout ;
wire \Mux59~1_combout ;
wire \Mux59~7_combout ;
wire \Mux59~8_combout ;
wire \Reg[26][4]~q ;
wire \Reg[18][4]~feeder_combout ;
wire \Reg[18][4]~q ;
wire \Mux59~2_combout ;
wire \Mux59~3_combout ;
wire \Mux59~4_combout ;
wire \Mux59~5_combout ;
wire \Mux59~6_combout ;
wire \Mux59~17_combout ;
wire \Mux59~18_combout ;
wire \Mux59~15_combout ;
wire \Mux59~13_combout ;
wire \Mux59~16_combout ;
wire \Mux59~10_combout ;
wire \Mux59~11_combout ;
wire \Reg[31][31]~feeder_combout ;
wire \Reg[31][31]~q ;
wire \Reg[27][31]~q ;
wire \Reg[23][31]~q ;
wire \Mux0~7_combout ;
wire \Mux0~8_combout ;
wire \Reg[25][31]~feeder_combout ;
wire \Reg[25][31]~q ;
wire \Reg[29][31]~q ;
wire \Reg[17][31]~feeder_combout ;
wire \Reg[17][31]~q ;
wire \Reg[21][31]~q ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \Reg[22][31]~feeder_combout ;
wire \Reg[22][31]~q ;
wire \Reg[26][31]~q ;
wire \Reg[18][31]~q ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \Reg[20][31]~feeder_combout ;
wire \Reg[20][31]~q ;
wire \Reg[28][31]~q ;
wire \Mux0~5_combout ;
wire \Mux0~6_combout ;
wire \Reg[15][31]~q ;
wire \Reg[12][31]~q ;
wire \Reg[13][31]~q ;
wire \Mux0~17_combout ;
wire \Reg[14][31]~q ;
wire \Mux0~18_combout ;
wire \Reg[11][31]~q ;
wire \Reg[9][31]~q ;
wire \Reg[10][31]~q ;
wire \Mux0~10_combout ;
wire \Mux0~11_combout ;
wire \Reg[2][31]~feeder_combout ;
wire \Reg[2][31]~q ;
wire \Reg[3][31]~q ;
wire \Reg[1][31]~q ;
wire \Mux0~14_combout ;
wire \Mux0~15_combout ;
wire \Reg[6][31]~q ;
wire \Reg[7][31]~q ;
wire \Reg[4][31]~q ;
wire \Reg[5][31]~q ;
wire \Mux0~12_combout ;
wire \Mux0~13_combout ;
wire \Mux0~16_combout ;
wire \Reg[29][29]~feeder_combout ;
wire \Reg[29][29]~q ;
wire \Reg[25][29]~feeder_combout ;
wire \Reg[25][29]~q ;
wire \Reg[21][29]~feeder_combout ;
wire \Reg[21][29]~q ;
wire \Reg[17][29]~q ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \Reg[23][29]~feeder_combout ;
wire \Reg[23][29]~q ;
wire \Reg[19][29]~q ;
wire \Mux2~7_combout ;
wire \Reg[31][29]~q ;
wire \Reg[27][29]~q ;
wire \Mux2~8_combout ;
wire \Reg[22][29]~q ;
wire \Reg[30][29]~q ;
wire \Reg[18][29]~q ;
wire \Reg[26][29]~q ;
wire \Mux2~2_combout ;
wire \Mux2~3_combout ;
wire \Reg[28][29]~q ;
wire \Reg[24][29]~q ;
wire \Mux2~4_combout ;
wire \Mux2~5_combout ;
wire \Mux2~6_combout ;
wire \Reg[2][29]~q ;
wire \Reg[3][29]~q ;
wire \Mux2~14_combout ;
wire \Mux2~15_combout ;
wire \Reg[4][29]~q ;
wire \Reg[5][29]~q ;
wire \Mux2~12_combout ;
wire \Reg[6][29]~q ;
wire \Reg[7][29]~feeder_combout ;
wire \Reg[7][29]~q ;
wire \Mux2~13_combout ;
wire \Mux2~16_combout ;
wire \Reg[15][29]~q ;
wire \Reg[14][29]~q ;
wire \Reg[12][29]~q ;
wire \Reg[13][29]~q ;
wire \Mux2~17_combout ;
wire \Mux2~18_combout ;
wire \Reg[11][29]~q ;
wire \Reg[9][29]~q ;
wire \Reg[10][29]~q ;
wire \Reg[8][29]~q ;
wire \Mux2~10_combout ;
wire \Mux2~11_combout ;
wire \Reg[21][30]~q ;
wire \Reg[29][30]~q ;
wire \Reg[25][30]~q ;
wire \Reg[17][30]~q ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Reg[24][30]~q ;
wire \Reg[28][30]~q ;
wire \Reg[16][30]~feeder_combout ;
wire \Reg[16][30]~q ;
wire \Reg[20][30]~q ;
wire \Mux1~4_combout ;
wire \Mux1~5_combout ;
wire \Reg[22][30]~q ;
wire \Reg[18][30]~q ;
wire \Mux1~2_combout ;
wire \Reg[30][30]~q ;
wire \Reg[26][30]~feeder_combout ;
wire \Reg[26][30]~q ;
wire \Mux1~3_combout ;
wire \Mux1~6_combout ;
wire \Reg[31][30]~q ;
wire \Reg[23][30]~q ;
wire \Reg[19][30]~q ;
wire \Mux1~7_combout ;
wire \Mux1~8_combout ;
wire \Reg[6][30]~feeder_combout ;
wire \Reg[6][30]~q ;
wire \Reg[5][30]~q ;
wire \Reg[4][30]~q ;
wire \Mux1~10_combout ;
wire \Reg[7][30]~q ;
wire \Mux1~11_combout ;
wire \Reg[15][30]~q ;
wire \Reg[13][30]~feeder_combout ;
wire \Reg[13][30]~q ;
wire \Reg[12][30]~q ;
wire \Mux1~17_combout ;
wire \Reg[14][30]~q ;
wire \Mux1~18_combout ;
wire \Reg[2][30]~q ;
wire \Mux1~15_combout ;
wire \Reg[11][30]~q ;
wire \Reg[9][30]~q ;
wire \Mux1~13_combout ;
wire \Mux1~16_combout ;
wire \Reg[31][28]~q ;
wire \Reg[23][28]~q ;
wire \Reg[19][28]~q ;
wire \Reg[27][28]~feeder_combout ;
wire \Reg[27][28]~q ;
wire \Mux3~7_combout ;
wire \Mux3~8_combout ;
wire \Reg[29][28]~feeder_combout ;
wire \Reg[29][28]~q ;
wire \Reg[21][28]~feeder_combout ;
wire \Reg[21][28]~q ;
wire \Reg[17][28]~feeder_combout ;
wire \Reg[17][28]~q ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \Reg[28][28]~q ;
wire \Reg[24][28]~feeder_combout ;
wire \Reg[24][28]~q ;
wire \Reg[20][28]~q ;
wire \Reg[16][28]~q ;
wire \Mux3~4_combout ;
wire \Mux3~5_combout ;
wire \Reg[26][28]~q ;
wire \Reg[30][28]~q ;
wire \Reg[22][28]~q ;
wire \Reg[18][28]~feeder_combout ;
wire \Reg[18][28]~q ;
wire \Mux3~2_combout ;
wire \Mux3~3_combout ;
wire \Mux3~6_combout ;
wire \Reg[6][28]~feeder_combout ;
wire \Reg[6][28]~q ;
wire \Reg[4][28]~q ;
wire \Reg[5][28]~q ;
wire \Mux3~10_combout ;
wire \Reg[7][28]~q ;
wire \Mux3~11_combout ;
wire \Reg[15][28]~q ;
wire \Reg[12][28]~q ;
wire \Reg[13][28]~q ;
wire \Mux3~17_combout ;
wire \Reg[14][28]~q ;
wire \Mux3~18_combout ;
wire \Reg[9][28]~q ;
wire \Reg[11][28]~q ;
wire \Mux3~13_combout ;
wire \Reg[1][28]~q ;
wire \Reg[3][28]~q ;
wire \Mux3~14_combout ;
wire \Reg[2][28]~q ;
wire \Mux3~15_combout ;
wire \Mux3~16_combout ;
wire \Reg[23][26]~q ;
wire \Reg[31][26]~feeder_combout ;
wire \Reg[31][26]~q ;
wire \Reg[19][26]~q ;
wire \Mux5~7_combout ;
wire \Mux5~8_combout ;
wire \Reg[16][26]~feeder_combout ;
wire \Reg[16][26]~q ;
wire \Reg[20][26]~q ;
wire \Mux5~4_combout ;
wire \Reg[28][26]~q ;
wire \Reg[24][26]~q ;
wire \Mux5~5_combout ;
wire \Reg[18][26]~q ;
wire \Reg[22][26]~feeder_combout ;
wire \Reg[22][26]~q ;
wire \Mux5~2_combout ;
wire \Reg[26][26]~q ;
wire \Mux5~3_combout ;
wire \Mux5~6_combout ;
wire \Reg[25][26]~q ;
wire \Reg[17][26]~q ;
wire \Mux5~0_combout ;
wire \Reg[29][26]~q ;
wire \Reg[21][26]~q ;
wire \Mux5~1_combout ;
wire \Reg[12][26]~feeder_combout ;
wire \Reg[12][26]~q ;
wire \Reg[13][26]~q ;
wire \Mux5~17_combout ;
wire \Reg[15][26]~q ;
wire \Reg[14][26]~q ;
wire \Mux5~18_combout ;
wire \Reg[7][26]~q ;
wire \Reg[6][26]~q ;
wire \Reg[5][26]~q ;
wire \Mux5~10_combout ;
wire \Mux5~11_combout ;
wire \Reg[3][26]~q ;
wire \Reg[1][26]~q ;
wire \Mux5~14_combout ;
wire \Reg[2][26]~q ;
wire \Mux5~15_combout ;
wire \Reg[11][26]~feeder_combout ;
wire \Reg[11][26]~q ;
wire \Reg[8][26]~q ;
wire \Reg[10][26]~q ;
wire \Mux5~12_combout ;
wire \Reg[9][26]~feeder_combout ;
wire \Reg[9][26]~q ;
wire \Mux5~13_combout ;
wire \Mux5~16_combout ;
wire \Reg[25][27]~q ;
wire \Reg[29][27]~q ;
wire \Reg[17][27]~q ;
wire \Reg[21][27]~q ;
wire \Mux4~0_combout ;
wire \Mux4~1_combout ;
wire \Reg[27][27]~q ;
wire \Reg[23][27]~feeder_combout ;
wire \Reg[23][27]~q ;
wire \Reg[19][27]~q ;
wire \Mux4~7_combout ;
wire \Reg[31][27]~q ;
wire \Mux4~8_combout ;
wire \Reg[20][27]~feeder_combout ;
wire \Reg[20][27]~q ;
wire \Reg[24][27]~q ;
wire \Mux4~4_combout ;
wire \Mux4~5_combout ;
wire \Reg[22][27]~q ;
wire \Reg[18][27]~q ;
wire \Reg[26][27]~feeder_combout ;
wire \Reg[26][27]~q ;
wire \Mux4~2_combout ;
wire \Mux4~3_combout ;
wire \Mux4~6_combout ;
wire \Reg[11][27]~q ;
wire \Reg[9][27]~q ;
wire \Reg[10][27]~q ;
wire \Reg[8][27]~q ;
wire \Mux4~10_combout ;
wire \Mux4~11_combout ;
wire \Reg[14][27]~feeder_combout ;
wire \Reg[14][27]~q ;
wire \Reg[12][27]~q ;
wire \Mux4~17_combout ;
wire \Reg[15][27]~feeder_combout ;
wire \Reg[15][27]~q ;
wire \Mux4~18_combout ;
wire \Reg[6][27]~q ;
wire \Reg[7][27]~q ;
wire \Reg[5][27]~q ;
wire \Reg[4][27]~q ;
wire \Mux4~12_combout ;
wire \Mux4~13_combout ;
wire \Reg[3][27]~q ;
wire \Reg[1][27]~q ;
wire \Mux4~14_combout ;
wire \Reg[2][27]~q ;
wire \Mux4~15_combout ;
wire \Mux4~16_combout ;
wire \Reg[31][25]~feeder_combout ;
wire \Reg[31][25]~q ;
wire \Reg[27][25]~q ;
wire \Reg[23][25]~q ;
wire \Reg[19][25]~q ;
wire \Mux6~7_combout ;
wire \Mux6~8_combout ;
wire \Reg[22][25]~q ;
wire \Reg[30][25]~q ;
wire \Reg[18][25]~q ;
wire \Reg[26][25]~feeder_combout ;
wire \Reg[26][25]~q ;
wire \Mux6~2_combout ;
wire \Mux6~3_combout ;
wire \Reg[28][25]~q ;
wire \Reg[20][25]~q ;
wire \Reg[24][25]~q ;
wire \Mux6~4_combout ;
wire \Mux6~5_combout ;
wire \Mux6~6_combout ;
wire \Reg[25][25]~q ;
wire \Reg[29][25]~q ;
wire \Reg[17][25]~q ;
wire \Reg[21][25]~q ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \Reg[9][25]~feeder_combout ;
wire \Reg[9][25]~q ;
wire \Reg[11][25]~q ;
wire \Reg[10][25]~q ;
wire \Mux6~10_combout ;
wire \Mux6~11_combout ;
wire \Reg[13][25]~q ;
wire \Reg[12][25]~feeder_combout ;
wire \Reg[12][25]~q ;
wire \Mux6~17_combout ;
wire \Reg[14][25]~q ;
wire \Reg[15][25]~feeder_combout ;
wire \Reg[15][25]~q ;
wire \Mux6~18_combout ;
wire \Reg[3][25]~q ;
wire \Reg[1][25]~q ;
wire \Mux6~14_combout ;
wire \Reg[2][25]~q ;
wire \Mux6~15_combout ;
wire \Reg[7][25]~q ;
wire \Reg[4][25]~q ;
wire \Reg[5][25]~q ;
wire \Mux6~12_combout ;
wire \Mux6~13_combout ;
wire \Mux6~16_combout ;
wire \Reg[18][24]~feeder_combout ;
wire \Reg[18][24]~q ;
wire \Reg[22][24]~feeder_combout ;
wire \Reg[22][24]~q ;
wire \Mux7~2_combout ;
wire \Reg[26][24]~q ;
wire \Reg[30][24]~feeder_combout ;
wire \Reg[30][24]~q ;
wire \Mux7~3_combout ;
wire \Reg[16][24]~q ;
wire \Mux7~4_combout ;
wire \Reg[24][24]~q ;
wire \Mux7~5_combout ;
wire \Mux7~6_combout ;
wire \Reg[21][24]~q ;
wire \Reg[29][24]~q ;
wire \Reg[25][24]~q ;
wire \Reg[17][24]~q ;
wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \Reg[31][24]~q ;
wire \Reg[27][24]~q ;
wire \Reg[19][24]~q ;
wire \Mux7~7_combout ;
wire \Reg[23][24]~q ;
wire \Mux7~8_combout ;
wire \Reg[5][24]~q ;
wire \Mux7~10_combout ;
wire \Reg[6][24]~q ;
wire \Reg[7][24]~feeder_combout ;
wire \Reg[7][24]~q ;
wire \Mux7~11_combout ;
wire \Reg[14][24]~q ;
wire \Reg[15][24]~q ;
wire \Reg[12][24]~q ;
wire \Reg[13][24]~q ;
wire \Mux7~17_combout ;
wire \Mux7~18_combout ;
wire \Reg[1][24]~q ;
wire \Mux7~14_combout ;
wire \Reg[2][24]~feeder_combout ;
wire \Reg[2][24]~q ;
wire \Mux7~15_combout ;
wire \Reg[10][24]~q ;
wire \Reg[8][24]~q ;
wire \Mux7~12_combout ;
wire \Reg[11][24]~q ;
wire \Mux7~13_combout ;
wire \Mux7~16_combout ;
wire \Reg[31][22]~q ;
wire \Reg[23][22]~q ;
wire \Reg[27][22]~q ;
wire \Reg[19][22]~q ;
wire \Mux9~7_combout ;
wire \Mux9~8_combout ;
wire \Reg[16][22]~q ;
wire \Mux9~4_combout ;
wire \Reg[28][22]~q ;
wire \Reg[24][22]~q ;
wire \Mux9~5_combout ;
wire \Reg[30][22]~feeder_combout ;
wire \Reg[30][22]~q ;
wire \Reg[18][22]~q ;
wire \Reg[22][22]~q ;
wire \Mux9~2_combout ;
wire \Reg[26][22]~q ;
wire \Mux9~3_combout ;
wire \Mux9~6_combout ;
wire \Reg[21][22]~q ;
wire \Reg[29][22]~q ;
wire \Reg[17][22]~feeder_combout ;
wire \Reg[17][22]~q ;
wire \Mux9~0_combout ;
wire \Mux9~1_combout ;
wire \Reg[12][22]~q ;
wire \Reg[13][22]~q ;
wire \Mux9~17_combout ;
wire \Reg[15][22]~q ;
wire \Reg[14][22]~q ;
wire \Mux9~18_combout ;
wire \Reg[1][22]~feeder_combout ;
wire \Reg[1][22]~q ;
wire \Reg[3][22]~q ;
wire \Mux9~14_combout ;
wire \Reg[2][22]~q ;
wire \Mux9~15_combout ;
wire \Reg[11][22]~q ;
wire \Reg[10][22]~q ;
wire \Reg[8][22]~q ;
wire \Mux9~12_combout ;
wire \Mux9~13_combout ;
wire \Mux9~16_combout ;
wire \Reg[7][22]~q ;
wire \Reg[4][22]~q ;
wire \Reg[5][22]~q ;
wire \Mux9~10_combout ;
wire \Reg[6][22]~q ;
wire \Mux9~11_combout ;
wire \Reg[19][23]~q ;
wire \Reg[23][23]~q ;
wire \Mux8~7_combout ;
wire \Reg[27][23]~q ;
wire \Reg[31][23]~q ;
wire \Mux8~8_combout ;
wire \Reg[29][23]~feeder_combout ;
wire \Reg[29][23]~q ;
wire \Reg[17][23]~feeder_combout ;
wire \Reg[17][23]~q ;
wire \Mux8~0_combout ;
wire \Reg[25][23]~feeder_combout ;
wire \Reg[25][23]~q ;
wire \Mux8~1_combout ;
wire \Reg[22][23]~q ;
wire \Reg[26][23]~q ;
wire \Reg[18][23]~q ;
wire \Mux8~2_combout ;
wire \Mux8~3_combout ;
wire \Reg[28][23]~q ;
wire \Reg[16][23]~q ;
wire \Reg[24][23]~feeder_combout ;
wire \Reg[24][23]~q ;
wire \Mux8~4_combout ;
wire \Reg[20][23]~q ;
wire \Mux8~5_combout ;
wire \Mux8~6_combout ;
wire \Reg[15][23]~feeder_combout ;
wire \Reg[15][23]~q ;
wire \Reg[14][23]~q ;
wire \Reg[13][23]~q ;
wire \Reg[12][23]~q ;
wire \Mux8~17_combout ;
wire \Mux8~18_combout ;
wire \Reg[1][23]~q ;
wire \Mux8~14_combout ;
wire \Mux8~15_combout ;
wire \Reg[6][23]~feeder_combout ;
wire \Reg[6][23]~q ;
wire \Reg[7][23]~q ;
wire \Reg[5][23]~q ;
wire \Reg[4][23]~q ;
wire \Mux8~12_combout ;
wire \Mux8~13_combout ;
wire \Mux8~16_combout ;
wire \Reg[11][23]~q ;
wire \Reg[9][23]~q ;
wire \Reg[10][23]~q ;
wire \Mux8~10_combout ;
wire \Mux8~11_combout ;
wire \Reg[28][21]~q ;
wire \Reg[16][21]~q ;
wire \Mux10~4_combout ;
wire \Mux10~5_combout ;
wire \Reg[18][21]~q ;
wire \Mux10~2_combout ;
wire \Reg[22][21]~q ;
wire \Mux10~3_combout ;
wire \Mux10~6_combout ;
wire \Reg[27][21]~q ;
wire \Reg[31][21]~q ;
wire \Reg[23][21]~feeder_combout ;
wire \Reg[23][21]~q ;
wire \Reg[19][21]~q ;
wire \Mux10~7_combout ;
wire \Mux10~8_combout ;
wire \Reg[17][21]~q ;
wire \Reg[21][21]~q ;
wire \Mux10~0_combout ;
wire \Reg[29][21]~q ;
wire \Reg[25][21]~q ;
wire \Mux10~1_combout ;
wire \Reg[13][21]~q ;
wire \Reg[12][21]~q ;
wire \Mux10~17_combout ;
wire \Reg[14][21]~q ;
wire \Reg[15][21]~feeder_combout ;
wire \Reg[15][21]~q ;
wire \Mux10~18_combout ;
wire \Reg[6][21]~q ;
wire \Reg[7][21]~q ;
wire \Mux10~13_combout ;
wire \Reg[2][21]~q ;
wire \Reg[3][21]~q ;
wire \Reg[1][21]~q ;
wire \Mux10~14_combout ;
wire \Mux10~15_combout ;
wire \Mux10~16_combout ;
wire \Reg[11][21]~q ;
wire \Reg[8][21]~q ;
wire \Reg[10][21]~q ;
wire \Mux10~10_combout ;
wire \Reg[9][21]~q ;
wire \Mux10~11_combout ;
wire \Reg[30][20]~q ;
wire \Reg[18][20]~q ;
wire \Reg[22][20]~feeder_combout ;
wire \Reg[22][20]~q ;
wire \Mux11~2_combout ;
wire \Reg[26][20]~q ;
wire \Mux11~3_combout ;
wire \Reg[16][20]~q ;
wire \Mux11~4_combout ;
wire \Reg[28][20]~q ;
wire \Mux11~5_combout ;
wire \Mux11~6_combout ;
wire \Reg[23][20]~q ;
wire \Reg[31][20]~feeder_combout ;
wire \Reg[31][20]~q ;
wire \Reg[19][20]~q ;
wire \Reg[27][20]~feeder_combout ;
wire \Reg[27][20]~q ;
wire \Mux11~7_combout ;
wire \Mux11~8_combout ;
wire \Reg[21][20]~feeder_combout ;
wire \Reg[21][20]~q ;
wire \Reg[29][20]~q ;
wire \Reg[17][20]~q ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \Reg[14][20]~q ;
wire \Reg[12][20]~q ;
wire \Reg[13][20]~q ;
wire \Mux11~17_combout ;
wire \Reg[15][20]~q ;
wire \Mux11~18_combout ;
wire \Reg[7][20]~q ;
wire \Reg[6][20]~q ;
wire \Reg[5][20]~q ;
wire \Mux11~10_combout ;
wire \Mux11~11_combout ;
wire \Reg[2][20]~q ;
wire \Mux11~15_combout ;
wire \Reg[9][20]~q ;
wire \Reg[11][20]~q ;
wire \Reg[10][20]~q ;
wire \Reg[8][20]~q ;
wire \Mux11~12_combout ;
wire \Mux11~13_combout ;
wire \Mux11~16_combout ;
wire \Reg[18][18]~q ;
wire \Reg[22][18]~feeder_combout ;
wire \Reg[22][18]~q ;
wire \Mux13~2_combout ;
wire \Reg[30][18]~q ;
wire \Reg[26][18]~q ;
wire \Mux13~3_combout ;
wire \Reg[24][18]~q ;
wire \Reg[28][18]~q ;
wire \Mux13~5_combout ;
wire \Mux13~6_combout ;
wire \Reg[31][18]~feeder_combout ;
wire \Reg[31][18]~q ;
wire \Reg[23][18]~q ;
wire \Reg[19][18]~q ;
wire \Reg[27][18]~feeder_combout ;
wire \Reg[27][18]~q ;
wire \Mux13~7_combout ;
wire \Mux13~8_combout ;
wire \Reg[21][18]~feeder_combout ;
wire \Reg[21][18]~q ;
wire \Reg[29][18]~q ;
wire \Reg[25][18]~feeder_combout ;
wire \Reg[25][18]~q ;
wire \Reg[17][18]~q ;
wire \Mux13~0_combout ;
wire \Mux13~1_combout ;
wire \Reg[14][18]~q ;
wire \Reg[15][18]~q ;
wire \Reg[13][18]~q ;
wire \Reg[12][18]~q ;
wire \Mux13~17_combout ;
wire \Mux13~18_combout ;
wire \Reg[5][18]~q ;
wire \Reg[4][18]~q ;
wire \Mux13~10_combout ;
wire \Reg[6][18]~q ;
wire \Reg[7][18]~q ;
wire \Mux13~11_combout ;
wire \Reg[9][18]~q ;
wire \Reg[11][18]~q ;
wire \Reg[10][18]~q ;
wire \Reg[8][18]~q ;
wire \Mux13~12_combout ;
wire \Mux13~13_combout ;
wire \Reg[1][18]~q ;
wire \Reg[3][18]~q ;
wire \Mux13~14_combout ;
wire \Reg[2][18]~q ;
wire \Mux13~15_combout ;
wire \Mux13~16_combout ;
wire \Reg[27][19]~q ;
wire \Reg[31][19]~q ;
wire \Reg[23][19]~feeder_combout ;
wire \Reg[23][19]~q ;
wire \Reg[19][19]~q ;
wire \Mux12~7_combout ;
wire \Mux12~8_combout ;
wire \Reg[17][19]~q ;
wire \Reg[21][19]~q ;
wire \Mux12~0_combout ;
wire \Reg[29][19]~q ;
wire \Reg[25][19]~q ;
wire \Mux12~1_combout ;
wire \Reg[22][19]~q ;
wire \Reg[26][19]~q ;
wire \Mux12~2_combout ;
wire \Mux12~3_combout ;
wire \Reg[20][19]~q ;
wire \Reg[16][19]~q ;
wire \Mux12~4_combout ;
wire \Mux12~5_combout ;
wire \Mux12~6_combout ;
wire \Reg[11][19]~q ;
wire \Reg[8][19]~q ;
wire \Reg[10][19]~q ;
wire \Mux12~10_combout ;
wire \Reg[9][19]~q ;
wire \Mux12~11_combout ;
wire \Reg[12][19]~q ;
wire \Reg[13][19]~q ;
wire \Mux12~17_combout ;
wire \Reg[15][19]~feeder_combout ;
wire \Reg[15][19]~q ;
wire \Reg[14][19]~q ;
wire \Mux12~18_combout ;
wire \Reg[6][19]~q ;
wire \Reg[7][19]~q ;
wire \Reg[4][19]~q ;
wire \Reg[5][19]~q ;
wire \Mux12~12_combout ;
wire \Mux12~13_combout ;
wire \Reg[1][19]~q ;
wire \Reg[3][19]~q ;
wire \Mux12~14_combout ;
wire \Reg[2][19]~q ;
wire \Mux12~15_combout ;
wire \Mux12~16_combout ;
wire \Reg[31][17]~q ;
wire \Reg[23][17]~feeder_combout ;
wire \Reg[23][17]~q ;
wire \Reg[19][17]~q ;
wire \Mux14~7_combout ;
wire \Reg[27][17]~q ;
wire \Mux14~8_combout ;
wire \Reg[28][17]~q ;
wire \Reg[24][17]~q ;
wire \Reg[16][17]~q ;
wire \Mux14~4_combout ;
wire \Mux14~5_combout ;
wire \Reg[22][17]~q ;
wire \Reg[26][17]~q ;
wire \Reg[18][17]~q ;
wire \Mux14~2_combout ;
wire \Mux14~3_combout ;
wire \Mux14~6_combout ;
wire \Reg[29][17]~q ;
wire \Reg[25][17]~q ;
wire \Reg[17][17]~q ;
wire \Reg[21][17]~q ;
wire \Mux14~0_combout ;
wire \Mux14~1_combout ;
wire \Reg[6][17]~q ;
wire \Reg[7][17]~q ;
wire \Mux14~13_combout ;
wire \Reg[1][17]~q ;
wire \Reg[3][17]~q ;
wire \Mux14~14_combout ;
wire \Reg[2][17]~q ;
wire \Mux14~15_combout ;
wire \Mux14~16_combout ;
wire \Reg[11][17]~q ;
wire \Reg[9][17]~q ;
wire \Reg[10][17]~q ;
wire \Reg[8][17]~q ;
wire \Mux14~10_combout ;
wire \Mux14~11_combout ;
wire \Reg[14][17]~feeder_combout ;
wire \Reg[14][17]~q ;
wire \Reg[15][17]~feeder_combout ;
wire \Reg[15][17]~q ;
wire \Reg[12][17]~q ;
wire \Reg[13][17]~q ;
wire \Mux14~17_combout ;
wire \Mux14~18_combout ;
wire \Mux32~0_combout ;
wire \Mux32~1_combout ;
wire \Reg[30][31]~q ;
wire \Mux32~3_combout ;
wire \Reg[16][31]~q ;
wire \Mux32~4_combout ;
wire \Mux32~5_combout ;
wire \Mux32~6_combout ;
wire \Reg[19][31]~q ;
wire \Mux32~7_combout ;
wire \Mux32~8_combout ;
wire \Mux32~17_combout ;
wire \Mux32~18_combout ;
wire \Mux32~10_combout ;
wire \Mux32~11_combout ;
wire \Mux32~15_combout ;
wire \Mux32~13_combout ;
wire \Mux32~16_combout ;
wire \Reg[18][16]~q ;
wire \Mux47~2_combout ;
wire \Reg[22][16]~q ;
wire \Mux47~3_combout ;
wire \Reg[20][16]~q ;
wire \Mux47~4_combout ;
wire \Mux47~5_combout ;
wire \Mux47~6_combout ;
wire \Mux47~7_combout ;
wire \Mux47~8_combout ;
wire \Mux47~0_combout ;
wire \Mux47~1_combout ;
wire \Mux47~17_combout ;
wire \Mux47~18_combout ;
wire \Mux47~10_combout ;
wire \Mux47~11_combout ;
wire \Mux47~14_combout ;
wire \Mux47~15_combout ;
wire \Mux47~13_combout ;
wire \Mux47~16_combout ;
wire \Mux46~7_combout ;
wire \Mux46~8_combout ;
wire \Mux46~0_combout ;
wire \Mux46~1_combout ;
wire \Reg[20][17]~feeder_combout ;
wire \Reg[20][17]~q ;
wire \Mux46~4_combout ;
wire \Mux46~5_combout ;
wire \Reg[30][17]~feeder_combout ;
wire \Reg[30][17]~q ;
wire \Mux46~2_combout ;
wire \Mux46~3_combout ;
wire \Mux46~6_combout ;
wire \Mux46~17_combout ;
wire \Mux46~18_combout ;
wire \Mux46~15_combout ;
wire \Mux46~12_combout ;
wire \Mux46~13_combout ;
wire \Mux46~16_combout ;
wire \Reg[5][17]~q ;
wire \Reg[4][17]~q ;
wire \Mux46~10_combout ;
wire \Mux46~11_combout ;
wire \Reg[20][18]~q ;
wire \Reg[16][18]~q ;
wire \Mux45~4_combout ;
wire \Mux45~5_combout ;
wire \Mux45~2_combout ;
wire \Mux45~3_combout ;
wire \Mux45~6_combout ;
wire \Mux45~7_combout ;
wire \Mux45~8_combout ;
wire \Mux45~0_combout ;
wire \Mux45~1_combout ;
wire \Mux45~10_combout ;
wire \Mux45~11_combout ;
wire \Mux45~17_combout ;
wire \Mux45~18_combout ;
wire \Mux45~13_combout ;
wire \Mux45~15_combout ;
wire \Mux45~16_combout ;
wire \Mux44~0_combout ;
wire \Mux44~1_combout ;
wire \Mux44~7_combout ;
wire \Mux44~8_combout ;
wire \Reg[24][19]~q ;
wire \Mux44~4_combout ;
wire \Mux44~5_combout ;
wire \Reg[30][19]~q ;
wire \Reg[18][19]~q ;
wire \Mux44~2_combout ;
wire \Mux44~3_combout ;
wire \Mux44~6_combout ;
wire \Mux44~12_combout ;
wire \Mux44~13_combout ;
wire \Mux44~14_combout ;
wire \Mux44~15_combout ;
wire \Mux44~16_combout ;
wire \Mux44~17_combout ;
wire \Mux44~18_combout ;
wire \Mux44~10_combout ;
wire \Mux44~11_combout ;
wire \Mux43~7_combout ;
wire \Mux43~8_combout ;
wire \Mux43~0_combout ;
wire \Reg[25][20]~q ;
wire \Mux43~1_combout ;
wire \Mux43~2_combout ;
wire \Mux43~3_combout ;
wire \Reg[24][20]~q ;
wire \Mux43~4_combout ;
wire \Reg[20][20]~q ;
wire \Mux43~5_combout ;
wire \Mux43~6_combout ;
wire \Mux43~17_combout ;
wire \Mux43~18_combout ;
wire \Mux43~10_combout ;
wire \Mux43~11_combout ;
wire \Mux43~15_combout ;
wire \Mux43~13_combout ;
wire \Mux43~16_combout ;
wire \Mux42~7_combout ;
wire \Mux42~8_combout ;
wire \Mux42~0_combout ;
wire \Mux42~1_combout ;
wire \Reg[20][21]~q ;
wire \Mux42~4_combout ;
wire \Reg[24][21]~q ;
wire \Mux42~5_combout ;
wire \Reg[30][21]~q ;
wire \Mux42~2_combout ;
wire \Mux42~3_combout ;
wire \Mux42~6_combout ;
wire \Mux42~17_combout ;
wire \Mux42~18_combout ;
wire \Reg[5][21]~q ;
wire \Mux42~10_combout ;
wire \Mux42~11_combout ;
wire \Mux42~15_combout ;
wire \Mux42~12_combout ;
wire \Mux42~13_combout ;
wire \Mux42~16_combout ;
wire \Reg[20][22]~feeder_combout ;
wire \Reg[20][22]~q ;
wire \Mux41~4_combout ;
wire \Mux41~5_combout ;
wire \Mux41~2_combout ;
wire \Mux41~3_combout ;
wire \Mux41~6_combout ;
wire \Mux41~7_combout ;
wire \Mux41~8_combout ;
wire \Mux41~0_combout ;
wire \Reg[25][22]~q ;
wire \Mux41~1_combout ;
wire \Mux41~14_combout ;
wire \Mux41~15_combout ;
wire \Mux41~12_combout ;
wire \Mux41~13_combout ;
wire \Mux41~16_combout ;
wire \Reg[9][22]~feeder_combout ;
wire \Reg[9][22]~q ;
wire \Mux41~10_combout ;
wire \Mux41~11_combout ;
wire \Mux41~17_combout ;
wire \Mux41~18_combout ;
wire \Reg[21][23]~feeder_combout ;
wire \Reg[21][23]~q ;
wire \Mux40~0_combout ;
wire \Mux40~1_combout ;
wire \Mux40~7_combout ;
wire \Mux40~8_combout ;
wire \Reg[30][23]~q ;
wire \Mux40~2_combout ;
wire \Mux40~3_combout ;
wire \Mux40~5_combout ;
wire \Mux40~6_combout ;
wire \Mux40~10_combout ;
wire \Mux40~11_combout ;
wire \Reg[2][23]~q ;
wire \Mux40~15_combout ;
wire \Reg[8][23]~q ;
wire \Mux40~12_combout ;
wire \Mux40~13_combout ;
wire \Mux40~16_combout ;
wire \Mux40~17_combout ;
wire \Mux40~18_combout ;
wire \Mux39~7_combout ;
wire \Mux39~8_combout ;
wire \Mux39~4_combout ;
wire \Reg[28][24]~q ;
wire \Reg[20][24]~feeder_combout ;
wire \Reg[20][24]~q ;
wire \Mux39~5_combout ;
wire \Mux39~2_combout ;
wire \Mux39~3_combout ;
wire \Mux39~6_combout ;
wire \Mux39~0_combout ;
wire \Mux39~1_combout ;
wire \Mux39~17_combout ;
wire \Mux39~18_combout ;
wire \Mux39~15_combout ;
wire \Reg[4][24]~q ;
wire \Mux39~12_combout ;
wire \Mux39~13_combout ;
wire \Mux39~16_combout ;
wire \Mux39~10_combout ;
wire \Reg[9][24]~q ;
wire \Mux39~11_combout ;
wire \Mux38~7_combout ;
wire \Mux38~8_combout ;
wire \Reg[16][25]~q ;
wire \Mux38~4_combout ;
wire \Mux38~5_combout ;
wire \Mux38~2_combout ;
wire \Mux38~3_combout ;
wire \Mux38~6_combout ;
wire \Mux38~0_combout ;
wire \Mux38~1_combout ;
wire \Mux38~17_combout ;
wire \Mux38~18_combout ;
wire \Reg[6][25]~q ;
wire \Mux38~10_combout ;
wire \Mux38~11_combout ;
wire \Reg[8][25]~q ;
wire \Mux38~12_combout ;
wire \Mux38~13_combout ;
wire \Mux38~14_combout ;
wire \Mux38~15_combout ;
wire \Mux38~16_combout ;
wire \Mux37~0_combout ;
wire \Mux37~1_combout ;
wire \Reg[27][26]~feeder_combout ;
wire \Reg[27][26]~q ;
wire \Mux37~7_combout ;
wire \Mux37~8_combout ;
wire \Mux37~4_combout ;
wire \Mux37~5_combout ;
wire \Mux37~2_combout ;
wire \Mux37~3_combout ;
wire \Mux37~6_combout ;
wire \Mux37~14_combout ;
wire \Mux37~15_combout ;
wire \Mux37~13_combout ;
wire \Mux37~16_combout ;
wire \Mux37~10_combout ;
wire \Mux37~11_combout ;
wire \Mux37~17_combout ;
wire \Mux37~18_combout ;
wire \Reg[19][5]~q ;
wire \Mux58~7_combout ;
wire \Mux58~8_combout ;
wire \Mux58~0_combout ;
wire \Mux58~1_combout ;
wire \Mux58~3_combout ;
wire \Mux58~4_combout ;
wire \Mux58~5_combout ;
wire \Mux58~6_combout ;
wire \Mux58~10_combout ;
wire \Reg[6][5]~q ;
wire \Mux58~11_combout ;
wire \Reg[12][5]~q ;
wire \Mux58~17_combout ;
wire \Mux58~18_combout ;
wire \Mux58~14_combout ;
wire \Mux58~15_combout ;
wire \Reg[8][5]~q ;
wire \Mux58~12_combout ;
wire \Mux58~13_combout ;
wire \Mux58~16_combout ;
wire \Mux57~7_combout ;
wire \Mux57~8_combout ;
wire \Reg[17][6]~q ;
wire \Mux57~0_combout ;
wire \Mux57~1_combout ;
wire \Mux57~4_combout ;
wire \Mux57~5_combout ;
wire \Reg[30][6]~q ;
wire \Mux57~2_combout ;
wire \Mux57~3_combout ;
wire \Mux57~6_combout ;
wire \Mux57~10_combout ;
wire \Mux57~11_combout ;
wire \Mux57~17_combout ;
wire \Mux57~18_combout ;
wire \Mux57~12_combout ;
wire \Mux57~13_combout ;
wire \Reg[1][6]~q ;
wire \Mux57~14_combout ;
wire \Mux57~15_combout ;
wire \Mux57~16_combout ;
wire \Reg[24][7]~feeder_combout ;
wire \Reg[24][7]~q ;
wire \Reg[16][7]~q ;
wire \Mux56~4_combout ;
wire \Mux56~5_combout ;
wire \Mux56~2_combout ;
wire \Reg[30][7]~q ;
wire \Mux56~3_combout ;
wire \Mux56~6_combout ;
wire \Mux56~0_combout ;
wire \Reg[21][7]~feeder_combout ;
wire \Reg[21][7]~q ;
wire \Mux56~1_combout ;
wire \Mux56~7_combout ;
wire \Mux56~8_combout ;
wire \Reg[5][7]~q ;
wire \Reg[4][7]~q ;
wire \Mux56~10_combout ;
wire \Mux56~11_combout ;
wire \Reg[12][7]~q ;
wire \Mux56~17_combout ;
wire \Mux56~18_combout ;
wire \Reg[8][7]~q ;
wire \Mux56~12_combout ;
wire \Mux56~13_combout ;
wire \Mux56~14_combout ;
wire \Mux56~15_combout ;
wire \Mux56~16_combout ;
wire \Reg[19][8]~feeder_combout ;
wire \Reg[19][8]~q ;
wire \Mux55~7_combout ;
wire \Mux55~8_combout ;
wire \Mux55~0_combout ;
wire \Mux55~1_combout ;
wire \Reg[28][8]~q ;
wire \Mux55~4_combout ;
wire \Mux55~5_combout ;
wire \Mux55~2_combout ;
wire \Mux55~3_combout ;
wire \Mux55~6_combout ;
wire \Mux55~17_combout ;
wire \Mux55~18_combout ;
wire \Mux55~10_combout ;
wire \Reg[9][8]~feeder_combout ;
wire \Reg[9][8]~q ;
wire \Mux55~11_combout ;
wire \Mux55~14_combout ;
wire \Mux55~15_combout ;
wire \Mux55~12_combout ;
wire \Mux55~13_combout ;
wire \Mux55~16_combout ;
wire \Mux36~7_combout ;
wire \Mux36~8_combout ;
wire \Mux36~0_combout ;
wire \Mux36~1_combout ;
wire \Reg[16][27]~q ;
wire \Mux36~4_combout ;
wire \Mux36~5_combout ;
wire \Mux36~2_combout ;
wire \Reg[30][27]~feeder_combout ;
wire \Reg[30][27]~q ;
wire \Mux36~3_combout ;
wire \Mux36~6_combout ;
wire \Reg[13][27]~feeder_combout ;
wire \Reg[13][27]~q ;
wire \Mux36~17_combout ;
wire \Mux36~18_combout ;
wire \Mux36~10_combout ;
wire \Mux36~11_combout ;
wire \Mux36~12_combout ;
wire \Mux36~13_combout ;
wire \Mux36~14_combout ;
wire \Mux36~15_combout ;
wire \Mux36~16_combout ;
wire \Reg[25][28]~feeder_combout ;
wire \Reg[25][28]~q ;
wire \Mux35~0_combout ;
wire \Mux35~1_combout ;
wire \Mux35~7_combout ;
wire \Mux35~8_combout ;
wire \Mux35~2_combout ;
wire \Mux35~3_combout ;
wire \Mux35~5_combout ;
wire \Mux35~6_combout ;
wire \Mux35~17_combout ;
wire \Mux35~18_combout ;
wire \Reg[8][28]~q ;
wire \Reg[10][28]~q ;
wire \Mux35~10_combout ;
wire \Mux35~11_combout ;
wire \Mux35~15_combout ;
wire \Mux35~13_combout ;
wire \Mux35~16_combout ;
wire \Mux34~7_combout ;
wire \Mux34~8_combout ;
wire \Mux34~0_combout ;
wire \Mux34~1_combout ;
wire \Mux34~2_combout ;
wire \Mux34~3_combout ;
wire \Reg[16][29]~q ;
wire \Mux34~4_combout ;
wire \Mux34~5_combout ;
wire \Mux34~6_combout ;
wire \Mux34~10_combout ;
wire \Mux34~11_combout ;
wire \Reg[1][29]~q ;
wire \Mux34~14_combout ;
wire \Mux34~15_combout ;
wire \Mux34~12_combout ;
wire \Mux34~13_combout ;
wire \Mux34~16_combout ;
wire \Mux34~17_combout ;
wire \Mux34~18_combout ;
wire \Mux33~7_combout ;
wire \Reg[27][30]~feeder_combout ;
wire \Reg[27][30]~q ;
wire \Mux33~8_combout ;
wire \Mux33~5_combout ;
wire \Mux33~2_combout ;
wire \Mux33~3_combout ;
wire \Mux33~6_combout ;
wire \Mux33~0_combout ;
wire \Mux33~1_combout ;
wire \Mux33~17_combout ;
wire \Mux33~18_combout ;
wire \Reg[8][30]~q ;
wire \Reg[10][30]~q ;
wire \Mux33~10_combout ;
wire \Mux33~11_combout ;
wire \Reg[1][30]~q ;
wire \Mux33~14_combout ;
wire \Mux33~15_combout ;
wire \Mux33~13_combout ;
wire \Mux33~16_combout ;
wire \Mux54~7_combout ;
wire \Mux54~8_combout ;
wire \Mux54~0_combout ;
wire \Mux54~1_combout ;
wire \Reg[16][9]~q ;
wire \Mux54~4_combout ;
wire \Reg[28][9]~q ;
wire \Mux54~5_combout ;
wire \Reg[22][9]~q ;
wire \Mux54~2_combout ;
wire \Mux54~3_combout ;
wire \Mux54~6_combout ;
wire \Mux54~10_combout ;
wire \Mux54~11_combout ;
wire \Mux54~17_combout ;
wire \Mux54~18_combout ;
wire \Reg[1][9]~q ;
wire \Mux54~14_combout ;
wire \Mux54~15_combout ;
wire \Mux54~12_combout ;
wire \Mux54~13_combout ;
wire \Mux54~16_combout ;
wire \Mux49~7_combout ;
wire \Mux49~8_combout ;
wire \Mux49~0_combout ;
wire \Mux49~1_combout ;
wire \Reg[16][14]~q ;
wire \Mux49~4_combout ;
wire \Reg[20][14]~q ;
wire \Mux49~5_combout ;
wire \Mux49~2_combout ;
wire \Mux49~3_combout ;
wire \Mux49~6_combout ;
wire \Mux49~14_combout ;
wire \Mux49~15_combout ;
wire \Mux49~13_combout ;
wire \Mux49~16_combout ;
wire \Mux49~10_combout ;
wire \Mux49~11_combout ;
wire \Mux49~17_combout ;
wire \Mux49~18_combout ;
wire \Mux48~7_combout ;
wire \Mux48~8_combout ;
wire \Mux48~0_combout ;
wire \Mux48~1_combout ;
wire \Mux48~4_combout ;
wire \Mux48~5_combout ;
wire \Reg[18][15]~q ;
wire \Mux48~2_combout ;
wire \Mux48~3_combout ;
wire \Mux48~6_combout ;
wire \Mux48~13_combout ;
wire \Mux48~14_combout ;
wire \Mux48~15_combout ;
wire \Mux48~16_combout ;
wire \Mux48~17_combout ;
wire \Mux48~18_combout ;
wire \Reg[5][15]~q ;
wire \Reg[4][15]~q ;
wire \Mux48~10_combout ;
wire \Mux48~11_combout ;
wire \Mux53~7_combout ;
wire \Mux53~8_combout ;
wire \Mux53~4_combout ;
wire \Mux53~5_combout ;
wire \Reg[30][10]~q ;
wire \Mux53~3_combout ;
wire \Mux53~6_combout ;
wire \Mux53~0_combout ;
wire \Mux53~1_combout ;
wire \Reg[12][10]~q ;
wire \Mux53~17_combout ;
wire \Mux53~18_combout ;
wire \Mux53~12_combout ;
wire \Mux53~13_combout ;
wire \Mux53~14_combout ;
wire \Mux53~15_combout ;
wire \Mux53~16_combout ;
wire \Mux53~10_combout ;
wire \Reg[9][10]~feeder_combout ;
wire \Reg[9][10]~q ;
wire \Mux53~11_combout ;
wire \Mux52~7_combout ;
wire \Mux52~8_combout ;
wire \Mux52~3_combout ;
wire \Reg[16][11]~q ;
wire \Mux52~4_combout ;
wire \Reg[24][11]~q ;
wire \Mux52~5_combout ;
wire \Mux52~6_combout ;
wire \Mux52~0_combout ;
wire \Mux52~1_combout ;
wire \Mux52~14_combout ;
wire \Mux52~15_combout ;
wire \Reg[8][11]~q ;
wire \Mux52~12_combout ;
wire \Mux52~13_combout ;
wire \Mux52~16_combout ;
wire \Mux52~10_combout ;
wire \Mux52~11_combout ;
wire \Reg[12][11]~q ;
wire \Mux52~17_combout ;
wire \Mux52~18_combout ;
wire \Mux51~0_combout ;
wire \Mux51~1_combout ;
wire \Mux51~7_combout ;
wire \Mux51~8_combout ;
wire \Reg[18][12]~q ;
wire \Mux51~2_combout ;
wire \Mux51~3_combout ;
wire \Reg[24][12]~feeder_combout ;
wire \Reg[24][12]~q ;
wire \Mux51~4_combout ;
wire \Mux51~5_combout ;
wire \Mux51~6_combout ;
wire \Mux51~17_combout ;
wire \Mux51~18_combout ;
wire \Mux51~10_combout ;
wire \Mux51~11_combout ;
wire \Mux51~13_combout ;
wire \Mux51~15_combout ;
wire \Mux51~16_combout ;
wire \Mux50~0_combout ;
wire \Mux50~1_combout ;
wire \Mux50~7_combout ;
wire \Mux50~8_combout ;
wire \Mux50~4_combout ;
wire \Reg[28][13]~feeder_combout ;
wire \Reg[28][13]~q ;
wire \Mux50~5_combout ;
wire \Reg[22][13]~feeder_combout ;
wire \Reg[22][13]~q ;
wire \Mux50~2_combout ;
wire \Mux50~3_combout ;
wire \Mux50~6_combout ;
wire \Mux50~12_combout ;
wire \Mux50~13_combout ;
wire \Mux50~14_combout ;
wire \Mux50~15_combout ;
wire \Mux50~16_combout ;
wire \Mux50~17_combout ;
wire \Mux50~18_combout ;
wire \Reg[4][13]~q ;
wire \Reg[5][13]~q ;
wire \Mux50~10_combout ;
wire \Mux50~11_combout ;


// Location: LCCOMB_X59_Y39_N24
cycloneive_lcell_comb \Mux62~14 (
// Equation(s):
// \Mux62~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][1]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][1]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[3][1]~q ),
	.datad(\Reg[1][1]~q ),
	.cin(gnd),
	.combout(\Mux62~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~14 .lut_mask = 16'hA280;
defparam \Mux62~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N1
dffeas \Reg[3][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][4] .is_wysiwyg = "true";
defparam \Reg[3][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N3
dffeas \Reg[1][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][4] .is_wysiwyg = "true";
defparam \Reg[1][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N2
cycloneive_lcell_comb \Mux27~14 (
// Equation(s):
// \Mux27~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][4]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][4]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[1][4]~q ),
	.datad(\Reg[3][4]~q ),
	.cin(gnd),
	.combout(\Mux27~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~14 .lut_mask = 16'hA820;
defparam \Mux27~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N27
dffeas \Reg[1][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][3] .is_wysiwyg = "true";
defparam \Reg[1][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N26
cycloneive_lcell_comb \Mux28~14 (
// Equation(s):
// \Mux28~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][3]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][3]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[1][3]~q ),
	.datad(\Reg[3][3]~q ),
	.cin(gnd),
	.combout(\Mux28~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~14 .lut_mask = 16'hA820;
defparam \Mux28~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N26
cycloneive_lcell_comb \Mux61~2 (
// Equation(s):
// \Mux61~2_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[26][2]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[18][2]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[18][2]~q ),
	.datad(\Reg[26][2]~q ),
	.cin(gnd),
	.combout(\Mux61~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~2 .lut_mask = 16'hDC98;
defparam \Mux61~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N14
cycloneive_lcell_comb \Mux61~12 (
// Equation(s):
// \Mux61~12_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17) # ((\Reg[5][2]~q )))) # (!ifid_ifinstr_o_16 & (!ifid_ifinstr_o_17 & (\Reg[4][2]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[4][2]~q ),
	.datad(\Reg[5][2]~q ),
	.cin(gnd),
	.combout(\Mux61~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~12 .lut_mask = 16'hBA98;
defparam \Mux61~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N10
cycloneive_lcell_comb \Mux24~4 (
// Equation(s):
// \Mux24~4_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[24][7]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & (\Reg[16][7]~q )))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[16][7]~q ),
	.datad(\Reg[24][7]~q ),
	.cin(gnd),
	.combout(\Mux24~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~4 .lut_mask = 16'hBA98;
defparam \Mux24~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N10
cycloneive_lcell_comb \Mux24~12 (
// Equation(s):
// \Mux24~12_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[5][7]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[4][7]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[5][7]~q ),
	.datac(\Reg[4][7]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux24~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~12 .lut_mask = 16'hEE50;
defparam \Mux24~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N1
dffeas \Reg[3][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][6] .is_wysiwyg = "true";
defparam \Reg[3][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N0
cycloneive_lcell_comb \Mux25~14 (
// Equation(s):
// \Mux25~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][6]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][6]~q ))))

	.dataa(\Reg[1][6]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[3][6]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux25~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~14 .lut_mask = 16'hC088;
defparam \Mux25~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N26
cycloneive_lcell_comb \Mux60~2 (
// Equation(s):
// \Mux60~2_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Reg[22][3]~q ))) # (!ifid_ifinstr_o_18 & (\Reg[18][3]~q ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[18][3]~q ),
	.datad(\Reg[22][3]~q ),
	.cin(gnd),
	.combout(\Mux60~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~2 .lut_mask = 16'hDC98;
defparam \Mux60~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N2
cycloneive_lcell_comb \Mux15~2 (
// Equation(s):
// \Mux15~2_combout  = (ifid_ifinstr_o_23 & (((\Reg[22][16]~q ) # (ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (\Reg[18][16]~q  & ((!ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[18][16]~q ),
	.datac(\Reg[22][16]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux15~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~2 .lut_mask = 16'hAAE4;
defparam \Mux15~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N31
dffeas \Reg[28][16] (
	.clk(!CLK),
	.d(\Reg[28][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][16] .is_wysiwyg = "true";
defparam \Reg[28][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N31
dffeas \Reg[8][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][15] .is_wysiwyg = "true";
defparam \Reg[8][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N18
cycloneive_lcell_comb \Mux16~12 (
// Equation(s):
// \Mux16~12_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[5][15]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[4][15]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[4][15]~q ),
	.datad(\Reg[5][15]~q ),
	.cin(gnd),
	.combout(\Mux16~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~12 .lut_mask = 16'hDC98;
defparam \Mux16~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y36_N7
dffeas \Reg[30][14] (
	.clk(!CLK),
	.d(\Reg[30][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][14] .is_wysiwyg = "true";
defparam \Reg[30][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N16
cycloneive_lcell_comb \Mux17~4 (
// Equation(s):
// \Mux17~4_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & (\Reg[20][14]~q )) # (!ifid_ifinstr_o_23 & ((\Reg[16][14]~q )))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[20][14]~q ),
	.datad(\Reg[16][14]~q ),
	.cin(gnd),
	.combout(\Mux17~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~4 .lut_mask = 16'hD9C8;
defparam \Mux17~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N22
cycloneive_lcell_comb \Mux18~12 (
// Equation(s):
// \Mux18~12_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[5][13]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[4][13]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[4][13]~q ),
	.datad(\Reg[5][13]~q ),
	.cin(gnd),
	.combout(\Mux18~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~12 .lut_mask = 16'hDC98;
defparam \Mux18~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y31_N29
dffeas \Reg[22][11] (
	.clk(!CLK),
	.d(\Reg[22][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][11] .is_wysiwyg = "true";
defparam \Reg[22][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N16
cycloneive_lcell_comb \Mux20~4 (
// Equation(s):
// \Mux20~4_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Reg[24][11]~q ))) # (!ifid_ifinstr_o_24 & (\Reg[16][11]~q ))))

	.dataa(\Reg[16][11]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[24][11]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux20~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~4 .lut_mask = 16'hFC22;
defparam \Mux20~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y36_N27
dffeas \Reg[3][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][9] .is_wysiwyg = "true";
defparam \Reg[3][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N26
cycloneive_lcell_comb \Mux22~14 (
// Equation(s):
// \Mux22~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[3][9]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[1][9]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[3][9]~q ),
	.datad(\Reg[1][9]~q ),
	.cin(gnd),
	.combout(\Mux22~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~14 .lut_mask = 16'hA280;
defparam \Mux22~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N18
cycloneive_lcell_comb \Mux59~12 (
// Equation(s):
// \Mux59~12_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17) # ((\Reg[5][4]~q )))) # (!ifid_ifinstr_o_16 & (!ifid_ifinstr_o_17 & (\Reg[4][4]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[4][4]~q ),
	.datad(\Reg[5][4]~q ),
	.cin(gnd),
	.combout(\Mux59~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~12 .lut_mask = 16'hBA98;
defparam \Mux59~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N0
cycloneive_lcell_comb \Mux59~14 (
// Equation(s):
// \Mux59~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][4]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][4]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[3][4]~q ),
	.datad(\Reg[1][4]~q ),
	.cin(gnd),
	.combout(\Mux59~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~14 .lut_mask = 16'hA280;
defparam \Mux59~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y32_N25
dffeas \Reg[24][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][31] .is_wysiwyg = "true";
defparam \Reg[24][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N24
cycloneive_lcell_comb \Mux0~4 (
// Equation(s):
// \Mux0~4_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[24][31]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & ((\Reg[16][31]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[24][31]~q ),
	.datad(\Reg[16][31]~q ),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~4 .lut_mask = 16'hB9A8;
defparam \Mux0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N27
dffeas \Reg[8][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][31] .is_wysiwyg = "true";
defparam \Reg[8][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y34_N19
dffeas \Reg[20][29] (
	.clk(!CLK),
	.d(\Reg[20][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][29] .is_wysiwyg = "true";
defparam \Reg[20][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N14
cycloneive_lcell_comb \Mux1~12 (
// Equation(s):
// \Mux1~12_combout  = (ifid_ifinstr_o_21 & (ifid_ifinstr_o_22)) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[10][30]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[8][30]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[8][30]~q ),
	.datad(\Reg[10][30]~q ),
	.cin(gnd),
	.combout(\Mux1~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~12 .lut_mask = 16'hDC98;
defparam \Mux1~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N27
dffeas \Reg[3][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][30] .is_wysiwyg = "true";
defparam \Reg[3][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N26
cycloneive_lcell_comb \Mux1~14 (
// Equation(s):
// \Mux1~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[3][30]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[1][30]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[3][30]~q ),
	.datad(\Reg[1][30]~q ),
	.cin(gnd),
	.combout(\Mux1~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~14 .lut_mask = 16'hC480;
defparam \Mux1~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N14
cycloneive_lcell_comb \Mux3~12 (
// Equation(s):
// \Mux3~12_combout  = (ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21) # ((\Reg[10][28]~q )))) # (!ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & (\Reg[8][28]~q )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[8][28]~q ),
	.datad(\Reg[10][28]~q ),
	.cin(gnd),
	.combout(\Mux3~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~12 .lut_mask = 16'hBA98;
defparam \Mux3~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N13
dffeas \Reg[30][26] (
	.clk(!CLK),
	.d(\Reg[30][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][26] .is_wysiwyg = "true";
defparam \Reg[30][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N27
dffeas \Reg[4][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][26] .is_wysiwyg = "true";
defparam \Reg[4][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N13
dffeas \Reg[28][27] (
	.clk(!CLK),
	.d(\Reg[28][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][27] .is_wysiwyg = "true";
defparam \Reg[28][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y38_N13
dffeas \Reg[3][24] (
	.clk(!CLK),
	.d(\Reg[3][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][24] .is_wysiwyg = "true";
defparam \Reg[3][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N23
dffeas \Reg[3][23] (
	.clk(!CLK),
	.d(\Reg[3][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][23] .is_wysiwyg = "true";
defparam \Reg[3][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N27
dffeas \Reg[26][21] (
	.clk(!CLK),
	.d(\Reg[26][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][21] .is_wysiwyg = "true";
defparam \Reg[26][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y39_N27
dffeas \Reg[4][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][21] .is_wysiwyg = "true";
defparam \Reg[4][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N26
cycloneive_lcell_comb \Mux10~12 (
// Equation(s):
// \Mux10~12_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[5][21]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[4][21]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[4][21]~q ),
	.datad(\Reg[5][21]~q ),
	.cin(gnd),
	.combout(\Mux10~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~12 .lut_mask = 16'hDC98;
defparam \Mux10~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y39_N23
dffeas \Reg[4][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][20] .is_wysiwyg = "true";
defparam \Reg[4][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N15
dffeas \Reg[3][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][20] .is_wysiwyg = "true";
defparam \Reg[3][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N1
dffeas \Reg[1][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][20] .is_wysiwyg = "true";
defparam \Reg[1][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N0
cycloneive_lcell_comb \Mux11~14 (
// Equation(s):
// \Mux11~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[3][20]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[1][20]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[3][20]~q ),
	.datac(\Reg[1][20]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux11~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~14 .lut_mask = 16'h88A0;
defparam \Mux11~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N28
cycloneive_lcell_comb \Mux13~4 (
// Equation(s):
// \Mux13~4_combout  = (ifid_ifinstr_o_23 & ((\Reg[20][18]~q ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((\Reg[16][18]~q  & !ifid_ifinstr_o_24))))

	.dataa(\Reg[20][18]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[16][18]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux13~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~4 .lut_mask = 16'hCCB8;
defparam \Mux13~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N27
dffeas \Reg[28][19] (
	.clk(!CLK),
	.d(\Reg[28][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][19] .is_wysiwyg = "true";
defparam \Reg[28][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N2
cycloneive_lcell_comb \Mux14~12 (
// Equation(s):
// \Mux14~12_combout  = (ifid_ifinstr_o_21 & ((\Reg[5][17]~q ) # ((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & (((\Reg[4][17]~q  & !ifid_ifinstr_o_22))))

	.dataa(\Reg[5][17]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[4][17]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux14~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~12 .lut_mask = 16'hCCB8;
defparam \Mux14~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N2
cycloneive_lcell_comb \Mux32~2 (
// Equation(s):
// \Mux32~2_combout  = (ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19) # ((\Reg[22][31]~q )))) # (!ifid_ifinstr_o_18 & (!ifid_ifinstr_o_19 & (\Reg[18][31]~q )))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[18][31]~q ),
	.datad(\Reg[22][31]~q ),
	.cin(gnd),
	.combout(\Mux32~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~2 .lut_mask = 16'hBA98;
defparam \Mux32~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N26
cycloneive_lcell_comb \Mux32~12 (
// Equation(s):
// \Mux32~12_combout  = (ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16) # ((\Reg[10][31]~q )))) # (!ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & (\Reg[8][31]~q )))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[8][31]~q ),
	.datad(\Reg[10][31]~q ),
	.cin(gnd),
	.combout(\Mux32~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~12 .lut_mask = 16'hBA98;
defparam \Mux32~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N6
cycloneive_lcell_comb \Mux32~14 (
// Equation(s):
// \Mux32~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][31]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][31]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[3][31]~q ),
	.datac(\Reg[1][31]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux32~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~14 .lut_mask = 16'h88A0;
defparam \Mux32~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N10
cycloneive_lcell_comb \Mux47~12 (
// Equation(s):
// \Mux47~12_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17) # ((\Reg[5][16]~q )))) # (!ifid_ifinstr_o_16 & (!ifid_ifinstr_o_17 & (\Reg[4][16]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[4][16]~q ),
	.datad(\Reg[5][16]~q ),
	.cin(gnd),
	.combout(\Mux47~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~12 .lut_mask = 16'hBA98;
defparam \Mux47~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N10
cycloneive_lcell_comb \Mux46~14 (
// Equation(s):
// \Mux46~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][17]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][17]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[3][17]~q ),
	.datad(\Reg[1][17]~q ),
	.cin(gnd),
	.combout(\Mux46~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~14 .lut_mask = 16'hA280;
defparam \Mux46~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N2
cycloneive_lcell_comb \Mux45~12 (
// Equation(s):
// \Mux45~12_combout  = (ifid_ifinstr_o_16 & ((\Reg[5][18]~q ) # ((ifid_ifinstr_o_17)))) # (!ifid_ifinstr_o_16 & (((\Reg[4][18]~q  & !ifid_ifinstr_o_17))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[5][18]~q ),
	.datac(\Reg[4][18]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux45~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~12 .lut_mask = 16'hAAD8;
defparam \Mux45~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N12
cycloneive_lcell_comb \Mux45~14 (
// Equation(s):
// \Mux45~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[3][18]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[1][18]~q ))))

	.dataa(\Reg[1][18]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[3][18]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux45~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~14 .lut_mask = 16'hE200;
defparam \Mux45~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N22
cycloneive_lcell_comb \Mux43~12 (
// Equation(s):
// \Mux43~12_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[5][20]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[4][20]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[4][20]~q ),
	.datad(\Reg[5][20]~q ),
	.cin(gnd),
	.combout(\Mux43~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~12 .lut_mask = 16'hDC98;
defparam \Mux43~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N14
cycloneive_lcell_comb \Mux43~14 (
// Equation(s):
// \Mux43~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][20]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][20]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[3][20]~q ),
	.datad(\Reg[1][20]~q ),
	.cin(gnd),
	.combout(\Mux43~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~14 .lut_mask = 16'hA280;
defparam \Mux43~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N18
cycloneive_lcell_comb \Mux42~14 (
// Equation(s):
// \Mux42~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][21]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][21]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[3][21]~q ),
	.datad(\Reg[1][21]~q ),
	.cin(gnd),
	.combout(\Mux42~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~14 .lut_mask = 16'hA280;
defparam \Mux42~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N20
cycloneive_lcell_comb \Mux40~4 (
// Equation(s):
// \Mux40~4_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[20][23]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[16][23]~q )))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[20][23]~q ),
	.datad(\Reg[16][23]~q ),
	.cin(gnd),
	.combout(\Mux40~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~4 .lut_mask = 16'hD9C8;
defparam \Mux40~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N26
cycloneive_lcell_comb \Mux40~14 (
// Equation(s):
// \Mux40~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][23]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][23]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[3][23]~q ),
	.datad(\Reg[1][23]~q ),
	.cin(gnd),
	.combout(\Mux40~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~14 .lut_mask = 16'hA280;
defparam \Mux40~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N26
cycloneive_lcell_comb \Mux39~14 (
// Equation(s):
// \Mux39~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][24]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][24]~q )))))

	.dataa(\Reg[3][24]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[1][24]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux39~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~14 .lut_mask = 16'hB800;
defparam \Mux39~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N26
cycloneive_lcell_comb \Mux37~12 (
// Equation(s):
// \Mux37~12_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[5][26]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[4][26]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[5][26]~q ),
	.datac(\Reg[4][26]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux37~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~12 .lut_mask = 16'hEE50;
defparam \Mux37~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N12
cycloneive_lcell_comb \Mux58~2 (
// Equation(s):
// \Mux58~2_combout  = (ifid_ifinstr_o_18 & ((\Reg[22][5]~q ) # ((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (((\Reg[18][5]~q  & !ifid_ifinstr_o_19))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[22][5]~q ),
	.datac(\Reg[18][5]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux58~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~2 .lut_mask = 16'hAAD8;
defparam \Mux58~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N8
cycloneive_lcell_comb \Mux35~4 (
// Equation(s):
// \Mux35~4_combout  = (ifid_ifinstr_o_19 & ((\Reg[24][28]~q ) # ((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & (((\Reg[16][28]~q  & !ifid_ifinstr_o_18))))

	.dataa(\Reg[24][28]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[16][28]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux35~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~4 .lut_mask = 16'hCCB8;
defparam \Mux35~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N14
cycloneive_lcell_comb \Mux35~12 (
// Equation(s):
// \Mux35~12_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[5][28]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[4][28]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[4][28]~q ),
	.datad(\Reg[5][28]~q ),
	.cin(gnd),
	.combout(\Mux35~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~12 .lut_mask = 16'hDC98;
defparam \Mux35~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N10
cycloneive_lcell_comb \Mux35~14 (
// Equation(s):
// \Mux35~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[3][28]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[1][28]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[1][28]~q ),
	.datac(\Reg[3][28]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux35~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~14 .lut_mask = 16'hE400;
defparam \Mux35~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N16
cycloneive_lcell_comb \Mux33~4 (
// Equation(s):
// \Mux33~4_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[24][30]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[16][30]~q ))))

	.dataa(\Reg[16][30]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[24][30]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux33~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~4 .lut_mask = 16'hFC22;
defparam \Mux33~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N26
cycloneive_lcell_comb \Mux33~12 (
// Equation(s):
// \Mux33~12_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[5][30]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[4][30]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[5][30]~q ),
	.datac(\Reg[4][30]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux33~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~12 .lut_mask = 16'hEE50;
defparam \Mux33~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N10
cycloneive_lcell_comb \Mux49~12 (
// Equation(s):
// \Mux49~12_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[5][14]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[4][14]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[5][14]~q ),
	.datac(\Reg[4][14]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux49~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~12 .lut_mask = 16'hEE50;
defparam \Mux49~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N30
cycloneive_lcell_comb \Mux48~12 (
// Equation(s):
// \Mux48~12_combout  = (ifid_ifinstr_o_16 & (((ifid_ifinstr_o_17)))) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[10][15]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[8][15]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[10][15]~q ),
	.datac(\Reg[8][15]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux48~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~12 .lut_mask = 16'hEE50;
defparam \Mux48~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N30
cycloneive_lcell_comb \Mux53~2 (
// Equation(s):
// \Mux53~2_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[26][10]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[18][10]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[18][10]~q ),
	.datad(\Reg[26][10]~q ),
	.cin(gnd),
	.combout(\Mux53~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~2 .lut_mask = 16'hDC98;
defparam \Mux53~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N18
cycloneive_lcell_comb \Mux52~2 (
// Equation(s):
// \Mux52~2_combout  = (ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19) # ((\Reg[22][11]~q )))) # (!ifid_ifinstr_o_18 & (!ifid_ifinstr_o_19 & (\Reg[18][11]~q )))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[18][11]~q ),
	.datad(\Reg[22][11]~q ),
	.cin(gnd),
	.combout(\Mux52~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~2 .lut_mask = 16'hBA98;
defparam \Mux52~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N6
cycloneive_lcell_comb \Mux51~12 (
// Equation(s):
// \Mux51~12_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[5][12]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[4][12]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[4][12]~q ),
	.datad(\Reg[5][12]~q ),
	.cin(gnd),
	.combout(\Mux51~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~12 .lut_mask = 16'hDC98;
defparam \Mux51~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N2
cycloneive_lcell_comb \Mux51~14 (
// Equation(s):
// \Mux51~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[3][12]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[1][12]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[1][12]~q ),
	.datad(\Reg[3][12]~q ),
	.cin(gnd),
	.combout(\Mux51~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~14 .lut_mask = 16'hA820;
defparam \Mux51~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N30
cycloneive_lcell_comb \Reg[28][16]~feeder (
// Equation(s):
// \Reg[28][16]~feeder_combout  = \wdat~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat9),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[28][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[28][16]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[28][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N6
cycloneive_lcell_comb \Reg[30][14]~feeder (
// Equation(s):
// \Reg[30][14]~feeder_combout  = \wdat~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat11),
	.cin(gnd),
	.combout(\Reg[30][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[30][14]~feeder .lut_mask = 16'hFF00;
defparam \Reg[30][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N28
cycloneive_lcell_comb \Reg[22][11]~feeder (
// Equation(s):
// \Reg[22][11]~feeder_combout  = \wdat~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat14),
	.cin(gnd),
	.combout(\Reg[22][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[22][11]~feeder .lut_mask = 16'hFF00;
defparam \Reg[22][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N18
cycloneive_lcell_comb \Reg[20][29]~feeder (
// Equation(s):
// \Reg[20][29]~feeder_combout  = \wdat~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat18),
	.cin(gnd),
	.combout(\Reg[20][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[20][29]~feeder .lut_mask = 16'hFF00;
defparam \Reg[20][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N12
cycloneive_lcell_comb \Reg[30][26]~feeder (
// Equation(s):
// \Reg[30][26]~feeder_combout  = \wdat~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat21),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[30][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[30][26]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[30][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N12
cycloneive_lcell_comb \Reg[28][27]~feeder (
// Equation(s):
// \Reg[28][27]~feeder_combout  = \wdat~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat22),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[28][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[28][27]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[28][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N12
cycloneive_lcell_comb \Reg[3][24]~feeder (
// Equation(s):
// \Reg[3][24]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat24),
	.cin(gnd),
	.combout(\Reg[3][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[3][24]~feeder .lut_mask = 16'hFF00;
defparam \Reg[3][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N22
cycloneive_lcell_comb \Reg[3][23]~feeder (
// Equation(s):
// \Reg[3][23]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat26),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[3][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[3][23]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[3][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N26
cycloneive_lcell_comb \Reg[26][21]~feeder (
// Equation(s):
// \Reg[26][21]~feeder_combout  = \wdat~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat27),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[26][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[26][21]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[26][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N26
cycloneive_lcell_comb \Reg[28][19]~feeder (
// Equation(s):
// \Reg[28][19]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat30),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[28][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[28][19]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[28][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N4
cycloneive_lcell_comb \Mux62~9 (
// Equation(s):
// Mux62 = (ifid_ifinstr_o_16 & ((\Mux62~6_combout  & ((\Mux62~8_combout ))) # (!\Mux62~6_combout  & (\Mux62~1_combout )))) # (!ifid_ifinstr_o_16 & (((\Mux62~6_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux62~1_combout ),
	.datac(\Mux62~6_combout ),
	.datad(\Mux62~8_combout ),
	.cin(gnd),
	.combout(Mux62),
	.cout());
// synopsys translate_off
defparam \Mux62~9 .lut_mask = 16'hF858;
defparam \Mux62~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N18
cycloneive_lcell_comb \Mux62~19 (
// Equation(s):
// Mux621 = (ifid_ifinstr_o_18 & ((\Mux62~16_combout  & (\Mux62~18_combout )) # (!\Mux62~16_combout  & ((\Mux62~11_combout ))))) # (!ifid_ifinstr_o_18 & (((\Mux62~16_combout ))))

	.dataa(\Mux62~18_combout ),
	.datab(\Mux62~11_combout ),
	.datac(ifid_ifinstr_o_18),
	.datad(\Mux62~16_combout ),
	.cin(gnd),
	.combout(Mux621),
	.cout());
// synopsys translate_off
defparam \Mux62~19 .lut_mask = 16'hAFC0;
defparam \Mux62~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N2
cycloneive_lcell_comb \Mux30~9 (
// Equation(s):
// Mux30 = (ifid_ifinstr_o_21 & ((\Mux30~6_combout  & ((\Mux30~8_combout ))) # (!\Mux30~6_combout  & (\Mux30~1_combout )))) # (!ifid_ifinstr_o_21 & (((\Mux30~6_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux30~1_combout ),
	.datac(\Mux30~6_combout ),
	.datad(\Mux30~8_combout ),
	.cin(gnd),
	.combout(Mux30),
	.cout());
// synopsys translate_off
defparam \Mux30~9 .lut_mask = 16'hF858;
defparam \Mux30~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N8
cycloneive_lcell_comb \Mux30~19 (
// Equation(s):
// Mux301 = (\Mux30~16_combout  & (((\Mux30~18_combout ) # (!ifid_ifinstr_o_24)))) # (!\Mux30~16_combout  & (\Mux30~11_combout  & (ifid_ifinstr_o_24)))

	.dataa(\Mux30~11_combout ),
	.datab(\Mux30~16_combout ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Mux30~18_combout ),
	.cin(gnd),
	.combout(Mux301),
	.cout());
// synopsys translate_off
defparam \Mux30~19 .lut_mask = 16'hEC2C;
defparam \Mux30~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N22
cycloneive_lcell_comb \Mux63~9 (
// Equation(s):
// Mux63 = (ifid_ifinstr_o_16 & ((\Mux63~6_combout  & ((\Mux63~8_combout ))) # (!\Mux63~6_combout  & (\Mux63~1_combout )))) # (!ifid_ifinstr_o_16 & (((\Mux63~6_combout ))))

	.dataa(\Mux63~1_combout ),
	.datab(\Mux63~8_combout ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux63~6_combout ),
	.cin(gnd),
	.combout(Mux63),
	.cout());
// synopsys translate_off
defparam \Mux63~9 .lut_mask = 16'hCFA0;
defparam \Mux63~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N18
cycloneive_lcell_comb \Mux63~19 (
// Equation(s):
// Mux631 = (\Mux63~16_combout  & ((\Mux63~18_combout ) # ((!ifid_ifinstr_o_19)))) # (!\Mux63~16_combout  & (((\Mux63~11_combout  & ifid_ifinstr_o_19))))

	.dataa(\Mux63~18_combout ),
	.datab(\Mux63~16_combout ),
	.datac(\Mux63~11_combout ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(Mux631),
	.cout());
// synopsys translate_off
defparam \Mux63~19 .lut_mask = 16'hB8CC;
defparam \Mux63~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N18
cycloneive_lcell_comb \Mux31~9 (
// Equation(s):
// Mux31 = (ifid_ifinstr_o_21 & ((\Mux31~6_combout  & ((\Mux31~8_combout ))) # (!\Mux31~6_combout  & (\Mux31~1_combout )))) # (!ifid_ifinstr_o_21 & (((\Mux31~6_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux31~1_combout ),
	.datac(\Mux31~8_combout ),
	.datad(\Mux31~6_combout ),
	.cin(gnd),
	.combout(Mux31),
	.cout());
// synopsys translate_off
defparam \Mux31~9 .lut_mask = 16'hF588;
defparam \Mux31~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N20
cycloneive_lcell_comb \Mux31~19 (
// Equation(s):
// Mux311 = (ifid_ifinstr_o_23 & ((\Mux31~16_combout  & (\Mux31~18_combout )) # (!\Mux31~16_combout  & ((\Mux31~11_combout ))))) # (!ifid_ifinstr_o_23 & (((\Mux31~16_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux31~18_combout ),
	.datac(\Mux31~16_combout ),
	.datad(\Mux31~11_combout ),
	.cin(gnd),
	.combout(Mux311),
	.cout());
// synopsys translate_off
defparam \Mux31~19 .lut_mask = 16'hDAD0;
defparam \Mux31~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N10
cycloneive_lcell_comb \Mux29~9 (
// Equation(s):
// Mux29 = (ifid_ifinstr_o_21 & ((\Mux29~6_combout  & ((\Mux29~8_combout ))) # (!\Mux29~6_combout  & (\Mux29~1_combout )))) # (!ifid_ifinstr_o_21 & (((\Mux29~6_combout ))))

	.dataa(\Mux29~1_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux29~8_combout ),
	.datad(\Mux29~6_combout ),
	.cin(gnd),
	.combout(Mux29),
	.cout());
// synopsys translate_off
defparam \Mux29~9 .lut_mask = 16'hF388;
defparam \Mux29~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N6
cycloneive_lcell_comb \Mux29~19 (
// Equation(s):
// Mux291 = (ifid_ifinstr_o_23 & ((\Mux29~16_combout  & ((\Mux29~18_combout ))) # (!\Mux29~16_combout  & (\Mux29~11_combout )))) # (!ifid_ifinstr_o_23 & (((\Mux29~16_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux29~11_combout ),
	.datac(\Mux29~18_combout ),
	.datad(\Mux29~16_combout ),
	.cin(gnd),
	.combout(Mux291),
	.cout());
// synopsys translate_off
defparam \Mux29~19 .lut_mask = 16'hF588;
defparam \Mux29~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N30
cycloneive_lcell_comb \Mux27~9 (
// Equation(s):
// Mux27 = (ifid_ifinstr_o_21 & ((\Mux27~6_combout  & ((\Mux27~8_combout ))) # (!\Mux27~6_combout  & (\Mux27~1_combout )))) # (!ifid_ifinstr_o_21 & (((\Mux27~6_combout ))))

	.dataa(\Mux27~1_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux27~6_combout ),
	.datad(\Mux27~8_combout ),
	.cin(gnd),
	.combout(Mux27),
	.cout());
// synopsys translate_off
defparam \Mux27~9 .lut_mask = 16'hF838;
defparam \Mux27~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N0
cycloneive_lcell_comb \Mux27~19 (
// Equation(s):
// Mux271 = (\Mux27~16_combout  & (((\Mux27~18_combout )) # (!ifid_ifinstr_o_23))) # (!\Mux27~16_combout  & (ifid_ifinstr_o_23 & (\Mux27~11_combout )))

	.dataa(\Mux27~16_combout ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Mux27~11_combout ),
	.datad(\Mux27~18_combout ),
	.cin(gnd),
	.combout(Mux271),
	.cout());
// synopsys translate_off
defparam \Mux27~19 .lut_mask = 16'hEA62;
defparam \Mux27~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N26
cycloneive_lcell_comb \Mux28~9 (
// Equation(s):
// Mux28 = (ifid_ifinstr_o_21 & ((\Mux28~6_combout  & (\Mux28~8_combout )) # (!\Mux28~6_combout  & ((\Mux28~1_combout ))))) # (!ifid_ifinstr_o_21 & (((\Mux28~6_combout ))))

	.dataa(\Mux28~8_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux28~1_combout ),
	.datad(\Mux28~6_combout ),
	.cin(gnd),
	.combout(Mux28),
	.cout());
// synopsys translate_off
defparam \Mux28~9 .lut_mask = 16'hBBC0;
defparam \Mux28~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N24
cycloneive_lcell_comb \Mux28~19 (
// Equation(s):
// Mux281 = (\Mux28~16_combout  & ((\Mux28~18_combout ) # ((!ifid_ifinstr_o_24)))) # (!\Mux28~16_combout  & (((ifid_ifinstr_o_24 & \Mux28~11_combout ))))

	.dataa(\Mux28~16_combout ),
	.datab(\Mux28~18_combout ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Mux28~11_combout ),
	.cin(gnd),
	.combout(Mux281),
	.cout());
// synopsys translate_off
defparam \Mux28~19 .lut_mask = 16'hDA8A;
defparam \Mux28~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N8
cycloneive_lcell_comb \Mux61~9 (
// Equation(s):
// Mux61 = (ifid_ifinstr_o_16 & ((\Mux61~6_combout  & (\Mux61~8_combout )) # (!\Mux61~6_combout  & ((\Mux61~1_combout ))))) # (!ifid_ifinstr_o_16 & (\Mux61~6_combout ))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux61~6_combout ),
	.datac(\Mux61~8_combout ),
	.datad(\Mux61~1_combout ),
	.cin(gnd),
	.combout(Mux61),
	.cout());
// synopsys translate_off
defparam \Mux61~9 .lut_mask = 16'hE6C4;
defparam \Mux61~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N28
cycloneive_lcell_comb \Mux61~19 (
// Equation(s):
// Mux611 = (ifid_ifinstr_o_19 & ((\Mux61~16_combout  & ((\Mux61~18_combout ))) # (!\Mux61~16_combout  & (\Mux61~11_combout )))) # (!ifid_ifinstr_o_19 & (((\Mux61~16_combout ))))

	.dataa(\Mux61~11_combout ),
	.datab(\Mux61~18_combout ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux61~16_combout ),
	.cin(gnd),
	.combout(Mux611),
	.cout());
// synopsys translate_off
defparam \Mux61~19 .lut_mask = 16'hCFA0;
defparam \Mux61~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N22
cycloneive_lcell_comb \Mux23~9 (
// Equation(s):
// Mux23 = (ifid_ifinstr_o_21 & ((\Mux23~6_combout  & (\Mux23~8_combout )) # (!\Mux23~6_combout  & ((\Mux23~1_combout ))))) # (!ifid_ifinstr_o_21 & (\Mux23~6_combout ))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux23~6_combout ),
	.datac(\Mux23~8_combout ),
	.datad(\Mux23~1_combout ),
	.cin(gnd),
	.combout(Mux23),
	.cout());
// synopsys translate_off
defparam \Mux23~9 .lut_mask = 16'hE6C4;
defparam \Mux23~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N12
cycloneive_lcell_comb \Mux23~19 (
// Equation(s):
// Mux231 = (ifid_ifinstr_o_23 & ((\Mux23~16_combout  & ((\Mux23~18_combout ))) # (!\Mux23~16_combout  & (\Mux23~11_combout )))) # (!ifid_ifinstr_o_23 & (((\Mux23~16_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux23~11_combout ),
	.datac(\Mux23~18_combout ),
	.datad(\Mux23~16_combout ),
	.cin(gnd),
	.combout(Mux231),
	.cout());
// synopsys translate_off
defparam \Mux23~19 .lut_mask = 16'hF588;
defparam \Mux23~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N10
cycloneive_lcell_comb \Mux24~9 (
// Equation(s):
// Mux24 = (ifid_ifinstr_o_21 & ((\Mux24~6_combout  & (\Mux24~8_combout )) # (!\Mux24~6_combout  & ((\Mux24~1_combout ))))) # (!ifid_ifinstr_o_21 & (((\Mux24~6_combout ))))

	.dataa(\Mux24~8_combout ),
	.datab(\Mux24~1_combout ),
	.datac(ifid_ifinstr_o_21),
	.datad(\Mux24~6_combout ),
	.cin(gnd),
	.combout(Mux24),
	.cout());
// synopsys translate_off
defparam \Mux24~9 .lut_mask = 16'hAFC0;
defparam \Mux24~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N8
cycloneive_lcell_comb \Mux24~19 (
// Equation(s):
// Mux241 = (\Mux24~16_combout  & (((\Mux24~18_combout )) # (!ifid_ifinstr_o_24))) # (!\Mux24~16_combout  & (ifid_ifinstr_o_24 & ((\Mux24~11_combout ))))

	.dataa(\Mux24~16_combout ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Mux24~18_combout ),
	.datad(\Mux24~11_combout ),
	.cin(gnd),
	.combout(Mux241),
	.cout());
// synopsys translate_off
defparam \Mux24~19 .lut_mask = 16'hE6A2;
defparam \Mux24~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N0
cycloneive_lcell_comb \Mux25~9 (
// Equation(s):
// Mux25 = (\Mux25~6_combout  & (((\Mux25~8_combout ) # (!ifid_ifinstr_o_21)))) # (!\Mux25~6_combout  & (\Mux25~1_combout  & (ifid_ifinstr_o_21)))

	.dataa(\Mux25~6_combout ),
	.datab(\Mux25~1_combout ),
	.datac(ifid_ifinstr_o_21),
	.datad(\Mux25~8_combout ),
	.cin(gnd),
	.combout(Mux25),
	.cout());
// synopsys translate_off
defparam \Mux25~9 .lut_mask = 16'hEA4A;
defparam \Mux25~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N8
cycloneive_lcell_comb \Mux25~19 (
// Equation(s):
// Mux251 = (ifid_ifinstr_o_23 & ((\Mux25~16_combout  & (\Mux25~18_combout )) # (!\Mux25~16_combout  & ((\Mux25~11_combout ))))) # (!ifid_ifinstr_o_23 & (((\Mux25~16_combout ))))

	.dataa(\Mux25~18_combout ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Mux25~11_combout ),
	.datad(\Mux25~16_combout ),
	.cin(gnd),
	.combout(Mux251),
	.cout());
// synopsys translate_off
defparam \Mux25~19 .lut_mask = 16'hBBC0;
defparam \Mux25~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N28
cycloneive_lcell_comb \Mux26~9 (
// Equation(s):
// Mux26 = (ifid_ifinstr_o_21 & ((\Mux26~6_combout  & (\Mux26~8_combout )) # (!\Mux26~6_combout  & ((\Mux26~1_combout ))))) # (!ifid_ifinstr_o_21 & (((\Mux26~6_combout ))))

	.dataa(\Mux26~8_combout ),
	.datab(\Mux26~1_combout ),
	.datac(ifid_ifinstr_o_21),
	.datad(\Mux26~6_combout ),
	.cin(gnd),
	.combout(Mux26),
	.cout());
// synopsys translate_off
defparam \Mux26~9 .lut_mask = 16'hAFC0;
defparam \Mux26~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N22
cycloneive_lcell_comb \Mux26~19 (
// Equation(s):
// Mux261 = (\Mux26~16_combout  & (((\Mux26~18_combout ) # (!ifid_ifinstr_o_24)))) # (!\Mux26~16_combout  & (\Mux26~11_combout  & (ifid_ifinstr_o_24)))

	.dataa(\Mux26~16_combout ),
	.datab(\Mux26~11_combout ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Mux26~18_combout ),
	.cin(gnd),
	.combout(Mux261),
	.cout());
// synopsys translate_off
defparam \Mux26~19 .lut_mask = 16'hEA4A;
defparam \Mux26~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N14
cycloneive_lcell_comb \Mux60~9 (
// Equation(s):
// Mux60 = (\Mux60~6_combout  & ((\Mux60~8_combout ) # ((!ifid_ifinstr_o_16)))) # (!\Mux60~6_combout  & (((\Mux60~1_combout  & ifid_ifinstr_o_16))))

	.dataa(\Mux60~8_combout ),
	.datab(\Mux60~1_combout ),
	.datac(\Mux60~6_combout ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(Mux60),
	.cout());
// synopsys translate_off
defparam \Mux60~9 .lut_mask = 16'hACF0;
defparam \Mux60~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N28
cycloneive_lcell_comb \Mux60~19 (
// Equation(s):
// Mux601 = (ifid_ifinstr_o_18 & ((\Mux60~16_combout  & ((\Mux60~18_combout ))) # (!\Mux60~16_combout  & (\Mux60~11_combout )))) # (!ifid_ifinstr_o_18 & (((\Mux60~16_combout ))))

	.dataa(\Mux60~11_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Mux60~18_combout ),
	.datad(\Mux60~16_combout ),
	.cin(gnd),
	.combout(Mux601),
	.cout());
// synopsys translate_off
defparam \Mux60~19 .lut_mask = 16'hF388;
defparam \Mux60~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N24
cycloneive_lcell_comb \Mux15~9 (
// Equation(s):
// Mux15 = (ifid_ifinstr_o_21 & ((\Mux15~6_combout  & (\Mux15~8_combout )) # (!\Mux15~6_combout  & ((\Mux15~1_combout ))))) # (!ifid_ifinstr_o_21 & (((\Mux15~6_combout ))))

	.dataa(\Mux15~8_combout ),
	.datab(\Mux15~1_combout ),
	.datac(ifid_ifinstr_o_21),
	.datad(\Mux15~6_combout ),
	.cin(gnd),
	.combout(Mux15),
	.cout());
// synopsys translate_off
defparam \Mux15~9 .lut_mask = 16'hAFC0;
defparam \Mux15~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N14
cycloneive_lcell_comb \Mux15~19 (
// Equation(s):
// Mux151 = (ifid_ifinstr_o_23 & ((\Mux15~16_combout  & (\Mux15~18_combout )) # (!\Mux15~16_combout  & ((\Mux15~11_combout ))))) # (!ifid_ifinstr_o_23 & (((\Mux15~16_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux15~18_combout ),
	.datac(\Mux15~11_combout ),
	.datad(\Mux15~16_combout ),
	.cin(gnd),
	.combout(Mux151),
	.cout());
// synopsys translate_off
defparam \Mux15~19 .lut_mask = 16'hDDA0;
defparam \Mux15~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N12
cycloneive_lcell_comb \Mux16~9 (
// Equation(s):
// Mux16 = (ifid_ifinstr_o_21 & ((\Mux16~6_combout  & ((\Mux16~8_combout ))) # (!\Mux16~6_combout  & (\Mux16~1_combout )))) # (!ifid_ifinstr_o_21 & (((\Mux16~6_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux16~1_combout ),
	.datac(\Mux16~8_combout ),
	.datad(\Mux16~6_combout ),
	.cin(gnd),
	.combout(Mux16),
	.cout());
// synopsys translate_off
defparam \Mux16~9 .lut_mask = 16'hF588;
defparam \Mux16~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N22
cycloneive_lcell_comb \Mux16~19 (
// Equation(s):
// Mux161 = (ifid_ifinstr_o_24 & ((\Mux16~16_combout  & (\Mux16~18_combout )) # (!\Mux16~16_combout  & ((\Mux16~11_combout ))))) # (!ifid_ifinstr_o_24 & (\Mux16~16_combout ))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux16~16_combout ),
	.datac(\Mux16~18_combout ),
	.datad(\Mux16~11_combout ),
	.cin(gnd),
	.combout(Mux161),
	.cout());
// synopsys translate_off
defparam \Mux16~19 .lut_mask = 16'hE6C4;
defparam \Mux16~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N6
cycloneive_lcell_comb \Mux17~9 (
// Equation(s):
// Mux17 = (ifid_ifinstr_o_21 & ((\Mux17~6_combout  & ((\Mux17~8_combout ))) # (!\Mux17~6_combout  & (\Mux17~1_combout )))) # (!ifid_ifinstr_o_21 & (((\Mux17~6_combout ))))

	.dataa(\Mux17~1_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux17~6_combout ),
	.datad(\Mux17~8_combout ),
	.cin(gnd),
	.combout(Mux17),
	.cout());
// synopsys translate_off
defparam \Mux17~9 .lut_mask = 16'hF838;
defparam \Mux17~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N18
cycloneive_lcell_comb \Mux17~19 (
// Equation(s):
// Mux171 = (ifid_ifinstr_o_23 & ((\Mux17~16_combout  & (\Mux17~18_combout )) # (!\Mux17~16_combout  & ((\Mux17~11_combout ))))) # (!ifid_ifinstr_o_23 & (((\Mux17~16_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux17~18_combout ),
	.datac(\Mux17~11_combout ),
	.datad(\Mux17~16_combout ),
	.cin(gnd),
	.combout(Mux171),
	.cout());
// synopsys translate_off
defparam \Mux17~19 .lut_mask = 16'hDDA0;
defparam \Mux17~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N6
cycloneive_lcell_comb \Mux18~9 (
// Equation(s):
// Mux18 = (ifid_ifinstr_o_21 & ((\Mux18~6_combout  & (\Mux18~8_combout )) # (!\Mux18~6_combout  & ((\Mux18~1_combout ))))) # (!ifid_ifinstr_o_21 & (((\Mux18~6_combout ))))

	.dataa(\Mux18~8_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux18~1_combout ),
	.datad(\Mux18~6_combout ),
	.cin(gnd),
	.combout(Mux18),
	.cout());
// synopsys translate_off
defparam \Mux18~9 .lut_mask = 16'hBBC0;
defparam \Mux18~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N4
cycloneive_lcell_comb \Mux18~19 (
// Equation(s):
// Mux181 = (\Mux18~16_combout  & (((\Mux18~18_combout )) # (!ifid_ifinstr_o_24))) # (!\Mux18~16_combout  & (ifid_ifinstr_o_24 & ((\Mux18~11_combout ))))

	.dataa(\Mux18~16_combout ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Mux18~18_combout ),
	.datad(\Mux18~11_combout ),
	.cin(gnd),
	.combout(Mux181),
	.cout());
// synopsys translate_off
defparam \Mux18~19 .lut_mask = 16'hE6A2;
defparam \Mux18~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N8
cycloneive_lcell_comb \Mux19~9 (
// Equation(s):
// Mux19 = (ifid_ifinstr_o_21 & ((\Mux19~6_combout  & ((\Mux19~8_combout ))) # (!\Mux19~6_combout  & (\Mux19~1_combout )))) # (!ifid_ifinstr_o_21 & (((\Mux19~6_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux19~1_combout ),
	.datac(\Mux19~8_combout ),
	.datad(\Mux19~6_combout ),
	.cin(gnd),
	.combout(Mux19),
	.cout());
// synopsys translate_off
defparam \Mux19~9 .lut_mask = 16'hF588;
defparam \Mux19~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N14
cycloneive_lcell_comb \Mux19~19 (
// Equation(s):
// Mux191 = (ifid_ifinstr_o_23 & ((\Mux19~16_combout  & (\Mux19~18_combout )) # (!\Mux19~16_combout  & ((\Mux19~11_combout ))))) # (!ifid_ifinstr_o_23 & (((\Mux19~16_combout ))))

	.dataa(\Mux19~18_combout ),
	.datab(\Mux19~11_combout ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux19~16_combout ),
	.cin(gnd),
	.combout(Mux191),
	.cout());
// synopsys translate_off
defparam \Mux19~19 .lut_mask = 16'hAFC0;
defparam \Mux19~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N12
cycloneive_lcell_comb \Mux20~9 (
// Equation(s):
// Mux20 = (\Mux20~6_combout  & (((\Mux20~8_combout ) # (!ifid_ifinstr_o_21)))) # (!\Mux20~6_combout  & (\Mux20~1_combout  & ((ifid_ifinstr_o_21))))

	.dataa(\Mux20~6_combout ),
	.datab(\Mux20~1_combout ),
	.datac(\Mux20~8_combout ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(Mux20),
	.cout());
// synopsys translate_off
defparam \Mux20~9 .lut_mask = 16'hE4AA;
defparam \Mux20~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N20
cycloneive_lcell_comb \Mux20~19 (
// Equation(s):
// Mux201 = (ifid_ifinstr_o_24 & ((\Mux20~16_combout  & (\Mux20~18_combout )) # (!\Mux20~16_combout  & ((\Mux20~11_combout ))))) # (!ifid_ifinstr_o_24 & (((\Mux20~16_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux20~18_combout ),
	.datac(\Mux20~11_combout ),
	.datad(\Mux20~16_combout ),
	.cin(gnd),
	.combout(Mux201),
	.cout());
// synopsys translate_off
defparam \Mux20~19 .lut_mask = 16'hDDA0;
defparam \Mux20~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N6
cycloneive_lcell_comb \Mux21~9 (
// Equation(s):
// Mux21 = (ifid_ifinstr_o_21 & ((\Mux21~6_combout  & ((\Mux21~8_combout ))) # (!\Mux21~6_combout  & (\Mux21~1_combout )))) # (!ifid_ifinstr_o_21 & (((\Mux21~6_combout ))))

	.dataa(\Mux21~1_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux21~6_combout ),
	.datad(\Mux21~8_combout ),
	.cin(gnd),
	.combout(Mux21),
	.cout());
// synopsys translate_off
defparam \Mux21~9 .lut_mask = 16'hF838;
defparam \Mux21~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N20
cycloneive_lcell_comb \Mux21~19 (
// Equation(s):
// Mux211 = (ifid_ifinstr_o_23 & ((\Mux21~16_combout  & ((\Mux21~18_combout ))) # (!\Mux21~16_combout  & (\Mux21~11_combout )))) # (!ifid_ifinstr_o_23 & (((\Mux21~16_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux21~11_combout ),
	.datac(\Mux21~18_combout ),
	.datad(\Mux21~16_combout ),
	.cin(gnd),
	.combout(Mux211),
	.cout());
// synopsys translate_off
defparam \Mux21~19 .lut_mask = 16'hF588;
defparam \Mux21~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N28
cycloneive_lcell_comb \Mux22~9 (
// Equation(s):
// Mux22 = (\Mux22~6_combout  & (((\Mux22~8_combout ) # (!ifid_ifinstr_o_21)))) # (!\Mux22~6_combout  & (\Mux22~1_combout  & ((ifid_ifinstr_o_21))))

	.dataa(\Mux22~1_combout ),
	.datab(\Mux22~6_combout ),
	.datac(\Mux22~8_combout ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(Mux22),
	.cout());
// synopsys translate_off
defparam \Mux22~9 .lut_mask = 16'hE2CC;
defparam \Mux22~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N22
cycloneive_lcell_comb \Mux22~19 (
// Equation(s):
// Mux221 = (ifid_ifinstr_o_24 & ((\Mux22~16_combout  & (\Mux22~18_combout )) # (!\Mux22~16_combout  & ((\Mux22~11_combout ))))) # (!ifid_ifinstr_o_24 & (((\Mux22~16_combout ))))

	.dataa(\Mux22~18_combout ),
	.datab(\Mux22~11_combout ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Mux22~16_combout ),
	.cin(gnd),
	.combout(Mux221),
	.cout());
// synopsys translate_off
defparam \Mux22~19 .lut_mask = 16'hAFC0;
defparam \Mux22~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N10
cycloneive_lcell_comb \Mux59~9 (
// Equation(s):
// Mux59 = (ifid_ifinstr_o_16 & ((\Mux59~6_combout  & ((\Mux59~8_combout ))) # (!\Mux59~6_combout  & (\Mux59~1_combout )))) # (!ifid_ifinstr_o_16 & (((\Mux59~6_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux59~1_combout ),
	.datac(\Mux59~8_combout ),
	.datad(\Mux59~6_combout ),
	.cin(gnd),
	.combout(Mux59),
	.cout());
// synopsys translate_off
defparam \Mux59~9 .lut_mask = 16'hF588;
defparam \Mux59~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N18
cycloneive_lcell_comb \Mux59~19 (
// Equation(s):
// Mux591 = (ifid_ifinstr_o_19 & ((\Mux59~16_combout  & (\Mux59~18_combout )) # (!\Mux59~16_combout  & ((\Mux59~11_combout ))))) # (!ifid_ifinstr_o_19 & (((\Mux59~16_combout ))))

	.dataa(\Mux59~18_combout ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Mux59~16_combout ),
	.datad(\Mux59~11_combout ),
	.cin(gnd),
	.combout(Mux591),
	.cout());
// synopsys translate_off
defparam \Mux59~19 .lut_mask = 16'hBCB0;
defparam \Mux59~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N30
cycloneive_lcell_comb \Mux0~9 (
// Equation(s):
// Mux0 = (ifid_ifinstr_o_21 & ((\Mux0~6_combout  & (\Mux0~8_combout )) # (!\Mux0~6_combout  & ((\Mux0~1_combout ))))) # (!ifid_ifinstr_o_21 & (((\Mux0~6_combout ))))

	.dataa(\Mux0~8_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux0~1_combout ),
	.datad(\Mux0~6_combout ),
	.cin(gnd),
	.combout(Mux0),
	.cout());
// synopsys translate_off
defparam \Mux0~9 .lut_mask = 16'hBBC0;
defparam \Mux0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N18
cycloneive_lcell_comb \Mux0~19 (
// Equation(s):
// Mux01 = (ifid_ifinstr_o_24 & ((\Mux0~16_combout  & (\Mux0~18_combout )) # (!\Mux0~16_combout  & ((\Mux0~11_combout ))))) # (!ifid_ifinstr_o_24 & (((\Mux0~16_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux0~18_combout ),
	.datac(\Mux0~11_combout ),
	.datad(\Mux0~16_combout ),
	.cin(gnd),
	.combout(Mux01),
	.cout());
// synopsys translate_off
defparam \Mux0~19 .lut_mask = 16'hDDA0;
defparam \Mux0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N2
cycloneive_lcell_comb \Mux2~9 (
// Equation(s):
// Mux2 = (ifid_ifinstr_o_21 & ((\Mux2~6_combout  & ((\Mux2~8_combout ))) # (!\Mux2~6_combout  & (\Mux2~1_combout )))) # (!ifid_ifinstr_o_21 & (((\Mux2~6_combout ))))

	.dataa(\Mux2~1_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux2~8_combout ),
	.datad(\Mux2~6_combout ),
	.cin(gnd),
	.combout(Mux2),
	.cout());
// synopsys translate_off
defparam \Mux2~9 .lut_mask = 16'hF388;
defparam \Mux2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N26
cycloneive_lcell_comb \Mux2~19 (
// Equation(s):
// Mux210 = (\Mux2~16_combout  & ((\Mux2~18_combout ) # ((!ifid_ifinstr_o_24)))) # (!\Mux2~16_combout  & (((\Mux2~11_combout  & ifid_ifinstr_o_24))))

	.dataa(\Mux2~16_combout ),
	.datab(\Mux2~18_combout ),
	.datac(\Mux2~11_combout ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(Mux210),
	.cout());
// synopsys translate_off
defparam \Mux2~19 .lut_mask = 16'hD8AA;
defparam \Mux2~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N6
cycloneive_lcell_comb \Mux1~9 (
// Equation(s):
// Mux1 = (ifid_ifinstr_o_21 & ((\Mux1~6_combout  & ((\Mux1~8_combout ))) # (!\Mux1~6_combout  & (\Mux1~1_combout )))) # (!ifid_ifinstr_o_21 & (((\Mux1~6_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux1~1_combout ),
	.datac(\Mux1~6_combout ),
	.datad(\Mux1~8_combout ),
	.cin(gnd),
	.combout(Mux1),
	.cout());
// synopsys translate_off
defparam \Mux1~9 .lut_mask = 16'hF858;
defparam \Mux1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N30
cycloneive_lcell_comb \Mux1~19 (
// Equation(s):
// Mux11 = (ifid_ifinstr_o_23 & ((\Mux1~16_combout  & ((\Mux1~18_combout ))) # (!\Mux1~16_combout  & (\Mux1~11_combout )))) # (!ifid_ifinstr_o_23 & (((\Mux1~16_combout ))))

	.dataa(\Mux1~11_combout ),
	.datab(\Mux1~18_combout ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux1~16_combout ),
	.cin(gnd),
	.combout(Mux11),
	.cout());
// synopsys translate_off
defparam \Mux1~19 .lut_mask = 16'hCFA0;
defparam \Mux1~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N24
cycloneive_lcell_comb \Mux3~9 (
// Equation(s):
// Mux3 = (ifid_ifinstr_o_21 & ((\Mux3~6_combout  & (\Mux3~8_combout )) # (!\Mux3~6_combout  & ((\Mux3~1_combout ))))) # (!ifid_ifinstr_o_21 & (((\Mux3~6_combout ))))

	.dataa(\Mux3~8_combout ),
	.datab(\Mux3~1_combout ),
	.datac(ifid_ifinstr_o_21),
	.datad(\Mux3~6_combout ),
	.cin(gnd),
	.combout(Mux3),
	.cout());
// synopsys translate_off
defparam \Mux3~9 .lut_mask = 16'hAFC0;
defparam \Mux3~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N4
cycloneive_lcell_comb \Mux3~19 (
// Equation(s):
// Mux32 = (ifid_ifinstr_o_23 & ((\Mux3~16_combout  & ((\Mux3~18_combout ))) # (!\Mux3~16_combout  & (\Mux3~11_combout )))) # (!ifid_ifinstr_o_23 & (((\Mux3~16_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux3~11_combout ),
	.datac(\Mux3~18_combout ),
	.datad(\Mux3~16_combout ),
	.cin(gnd),
	.combout(Mux32),
	.cout());
// synopsys translate_off
defparam \Mux3~19 .lut_mask = 16'hF588;
defparam \Mux3~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N6
cycloneive_lcell_comb \Mux5~9 (
// Equation(s):
// Mux5 = (ifid_ifinstr_o_21 & ((\Mux5~6_combout  & (\Mux5~8_combout )) # (!\Mux5~6_combout  & ((\Mux5~1_combout ))))) # (!ifid_ifinstr_o_21 & (((\Mux5~6_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux5~8_combout ),
	.datac(\Mux5~6_combout ),
	.datad(\Mux5~1_combout ),
	.cin(gnd),
	.combout(Mux5),
	.cout());
// synopsys translate_off
defparam \Mux5~9 .lut_mask = 16'hDAD0;
defparam \Mux5~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N30
cycloneive_lcell_comb \Mux5~19 (
// Equation(s):
// Mux51 = (ifid_ifinstr_o_23 & ((\Mux5~16_combout  & (\Mux5~18_combout )) # (!\Mux5~16_combout  & ((\Mux5~11_combout ))))) # (!ifid_ifinstr_o_23 & (((\Mux5~16_combout ))))

	.dataa(\Mux5~18_combout ),
	.datab(\Mux5~11_combout ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux5~16_combout ),
	.cin(gnd),
	.combout(Mux51),
	.cout());
// synopsys translate_off
defparam \Mux5~19 .lut_mask = 16'hAFC0;
defparam \Mux5~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N12
cycloneive_lcell_comb \Mux4~9 (
// Equation(s):
// Mux4 = (ifid_ifinstr_o_21 & ((\Mux4~6_combout  & ((\Mux4~8_combout ))) # (!\Mux4~6_combout  & (\Mux4~1_combout )))) # (!ifid_ifinstr_o_21 & (((\Mux4~6_combout ))))

	.dataa(\Mux4~1_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux4~8_combout ),
	.datad(\Mux4~6_combout ),
	.cin(gnd),
	.combout(Mux4),
	.cout());
// synopsys translate_off
defparam \Mux4~9 .lut_mask = 16'hF388;
defparam \Mux4~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N0
cycloneive_lcell_comb \Mux4~19 (
// Equation(s):
// Mux41 = (ifid_ifinstr_o_24 & ((\Mux4~16_combout  & ((\Mux4~18_combout ))) # (!\Mux4~16_combout  & (\Mux4~11_combout )))) # (!ifid_ifinstr_o_24 & (((\Mux4~16_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux4~11_combout ),
	.datac(\Mux4~18_combout ),
	.datad(\Mux4~16_combout ),
	.cin(gnd),
	.combout(Mux41),
	.cout());
// synopsys translate_off
defparam \Mux4~19 .lut_mask = 16'hF588;
defparam \Mux4~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N24
cycloneive_lcell_comb \Mux6~9 (
// Equation(s):
// Mux6 = (ifid_ifinstr_o_21 & ((\Mux6~6_combout  & (\Mux6~8_combout )) # (!\Mux6~6_combout  & ((\Mux6~1_combout ))))) # (!ifid_ifinstr_o_21 & (((\Mux6~6_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux6~8_combout ),
	.datac(\Mux6~6_combout ),
	.datad(\Mux6~1_combout ),
	.cin(gnd),
	.combout(Mux6),
	.cout());
// synopsys translate_off
defparam \Mux6~9 .lut_mask = 16'hDAD0;
defparam \Mux6~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N4
cycloneive_lcell_comb \Mux6~19 (
// Equation(s):
// Mux64 = (ifid_ifinstr_o_24 & ((\Mux6~16_combout  & ((\Mux6~18_combout ))) # (!\Mux6~16_combout  & (\Mux6~11_combout )))) # (!ifid_ifinstr_o_24 & (((\Mux6~16_combout ))))

	.dataa(\Mux6~11_combout ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Mux6~18_combout ),
	.datad(\Mux6~16_combout ),
	.cin(gnd),
	.combout(Mux64),
	.cout());
// synopsys translate_off
defparam \Mux6~19 .lut_mask = 16'hF388;
defparam \Mux6~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N28
cycloneive_lcell_comb \Mux7~9 (
// Equation(s):
// Mux7 = (\Mux7~6_combout  & (((\Mux7~8_combout )) # (!ifid_ifinstr_o_21))) # (!\Mux7~6_combout  & (ifid_ifinstr_o_21 & (\Mux7~1_combout )))

	.dataa(\Mux7~6_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux7~1_combout ),
	.datad(\Mux7~8_combout ),
	.cin(gnd),
	.combout(Mux7),
	.cout());
// synopsys translate_off
defparam \Mux7~9 .lut_mask = 16'hEA62;
defparam \Mux7~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N12
cycloneive_lcell_comb \Mux7~19 (
// Equation(s):
// Mux71 = (ifid_ifinstr_o_23 & ((\Mux7~16_combout  & ((\Mux7~18_combout ))) # (!\Mux7~16_combout  & (\Mux7~11_combout )))) # (!ifid_ifinstr_o_23 & (((\Mux7~16_combout ))))

	.dataa(\Mux7~11_combout ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Mux7~18_combout ),
	.datad(\Mux7~16_combout ),
	.cin(gnd),
	.combout(Mux71),
	.cout());
// synopsys translate_off
defparam \Mux7~19 .lut_mask = 16'hF388;
defparam \Mux7~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N4
cycloneive_lcell_comb \Mux9~9 (
// Equation(s):
// Mux9 = (ifid_ifinstr_o_21 & ((\Mux9~6_combout  & (\Mux9~8_combout )) # (!\Mux9~6_combout  & ((\Mux9~1_combout ))))) # (!ifid_ifinstr_o_21 & (((\Mux9~6_combout ))))

	.dataa(\Mux9~8_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux9~6_combout ),
	.datad(\Mux9~1_combout ),
	.cin(gnd),
	.combout(Mux9),
	.cout());
// synopsys translate_off
defparam \Mux9~9 .lut_mask = 16'hBCB0;
defparam \Mux9~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N24
cycloneive_lcell_comb \Mux9~19 (
// Equation(s):
// Mux91 = (\Mux9~16_combout  & ((\Mux9~18_combout ) # ((!ifid_ifinstr_o_23)))) # (!\Mux9~16_combout  & (((\Mux9~11_combout  & ifid_ifinstr_o_23))))

	.dataa(\Mux9~18_combout ),
	.datab(\Mux9~16_combout ),
	.datac(\Mux9~11_combout ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(Mux91),
	.cout());
// synopsys translate_off
defparam \Mux9~19 .lut_mask = 16'hB8CC;
defparam \Mux9~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N2
cycloneive_lcell_comb \Mux8~9 (
// Equation(s):
// Mux8 = (ifid_ifinstr_o_21 & ((\Mux8~6_combout  & (\Mux8~8_combout )) # (!\Mux8~6_combout  & ((\Mux8~1_combout ))))) # (!ifid_ifinstr_o_21 & (((\Mux8~6_combout ))))

	.dataa(\Mux8~8_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux8~1_combout ),
	.datad(\Mux8~6_combout ),
	.cin(gnd),
	.combout(Mux8),
	.cout());
// synopsys translate_off
defparam \Mux8~9 .lut_mask = 16'hBBC0;
defparam \Mux8~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N10
cycloneive_lcell_comb \Mux8~19 (
// Equation(s):
// Mux81 = (\Mux8~16_combout  & ((\Mux8~18_combout ) # ((!ifid_ifinstr_o_24)))) # (!\Mux8~16_combout  & (((ifid_ifinstr_o_24 & \Mux8~11_combout ))))

	.dataa(\Mux8~18_combout ),
	.datab(\Mux8~16_combout ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Mux8~11_combout ),
	.cin(gnd),
	.combout(Mux81),
	.cout());
// synopsys translate_off
defparam \Mux8~19 .lut_mask = 16'hBC8C;
defparam \Mux8~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N16
cycloneive_lcell_comb \Mux10~9 (
// Equation(s):
// Mux10 = (\Mux10~6_combout  & ((\Mux10~8_combout ) # ((!ifid_ifinstr_o_21)))) # (!\Mux10~6_combout  & (((ifid_ifinstr_o_21 & \Mux10~1_combout ))))

	.dataa(\Mux10~6_combout ),
	.datab(\Mux10~8_combout ),
	.datac(ifid_ifinstr_o_21),
	.datad(\Mux10~1_combout ),
	.cin(gnd),
	.combout(Mux10),
	.cout());
// synopsys translate_off
defparam \Mux10~9 .lut_mask = 16'hDA8A;
defparam \Mux10~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N6
cycloneive_lcell_comb \Mux10~19 (
// Equation(s):
// Mux101 = (ifid_ifinstr_o_24 & ((\Mux10~16_combout  & (\Mux10~18_combout )) # (!\Mux10~16_combout  & ((\Mux10~11_combout ))))) # (!ifid_ifinstr_o_24 & (((\Mux10~16_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux10~18_combout ),
	.datac(\Mux10~16_combout ),
	.datad(\Mux10~11_combout ),
	.cin(gnd),
	.combout(Mux101),
	.cout());
// synopsys translate_off
defparam \Mux10~19 .lut_mask = 16'hDAD0;
defparam \Mux10~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N14
cycloneive_lcell_comb \Mux11~9 (
// Equation(s):
// Mux111 = (\Mux11~6_combout  & (((\Mux11~8_combout )) # (!ifid_ifinstr_o_21))) # (!\Mux11~6_combout  & (ifid_ifinstr_o_21 & ((\Mux11~1_combout ))))

	.dataa(\Mux11~6_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux11~8_combout ),
	.datad(\Mux11~1_combout ),
	.cin(gnd),
	.combout(Mux111),
	.cout());
// synopsys translate_off
defparam \Mux11~9 .lut_mask = 16'hE6A2;
defparam \Mux11~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N28
cycloneive_lcell_comb \Mux11~19 (
// Equation(s):
// Mux112 = (ifid_ifinstr_o_23 & ((\Mux11~16_combout  & (\Mux11~18_combout )) # (!\Mux11~16_combout  & ((\Mux11~11_combout ))))) # (!ifid_ifinstr_o_23 & (((\Mux11~16_combout ))))

	.dataa(\Mux11~18_combout ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Mux11~11_combout ),
	.datad(\Mux11~16_combout ),
	.cin(gnd),
	.combout(Mux112),
	.cout());
// synopsys translate_off
defparam \Mux11~19 .lut_mask = 16'hBBC0;
defparam \Mux11~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N26
cycloneive_lcell_comb \Mux13~9 (
// Equation(s):
// Mux13 = (\Mux13~6_combout  & (((\Mux13~8_combout )) # (!ifid_ifinstr_o_21))) # (!\Mux13~6_combout  & (ifid_ifinstr_o_21 & ((\Mux13~1_combout ))))

	.dataa(\Mux13~6_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux13~8_combout ),
	.datad(\Mux13~1_combout ),
	.cin(gnd),
	.combout(Mux13),
	.cout());
// synopsys translate_off
defparam \Mux13~9 .lut_mask = 16'hE6A2;
defparam \Mux13~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N24
cycloneive_lcell_comb \Mux13~19 (
// Equation(s):
// Mux131 = (\Mux13~16_combout  & ((\Mux13~18_combout ) # ((!ifid_ifinstr_o_23)))) # (!\Mux13~16_combout  & (((\Mux13~11_combout  & ifid_ifinstr_o_23))))

	.dataa(\Mux13~18_combout ),
	.datab(\Mux13~11_combout ),
	.datac(\Mux13~16_combout ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(Mux131),
	.cout());
// synopsys translate_off
defparam \Mux13~19 .lut_mask = 16'hACF0;
defparam \Mux13~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N12
cycloneive_lcell_comb \Mux12~9 (
// Equation(s):
// Mux12 = (ifid_ifinstr_o_21 & ((\Mux12~6_combout  & (\Mux12~8_combout )) # (!\Mux12~6_combout  & ((\Mux12~1_combout ))))) # (!ifid_ifinstr_o_21 & (((\Mux12~6_combout ))))

	.dataa(\Mux12~8_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux12~1_combout ),
	.datad(\Mux12~6_combout ),
	.cin(gnd),
	.combout(Mux12),
	.cout());
// synopsys translate_off
defparam \Mux12~9 .lut_mask = 16'hBBC0;
defparam \Mux12~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N18
cycloneive_lcell_comb \Mux12~19 (
// Equation(s):
// Mux121 = (ifid_ifinstr_o_24 & ((\Mux12~16_combout  & ((\Mux12~18_combout ))) # (!\Mux12~16_combout  & (\Mux12~11_combout )))) # (!ifid_ifinstr_o_24 & (((\Mux12~16_combout ))))

	.dataa(\Mux12~11_combout ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Mux12~18_combout ),
	.datad(\Mux12~16_combout ),
	.cin(gnd),
	.combout(Mux121),
	.cout());
// synopsys translate_off
defparam \Mux12~19 .lut_mask = 16'hF388;
defparam \Mux12~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N10
cycloneive_lcell_comb \Mux14~9 (
// Equation(s):
// Mux14 = (ifid_ifinstr_o_21 & ((\Mux14~6_combout  & (\Mux14~8_combout )) # (!\Mux14~6_combout  & ((\Mux14~1_combout ))))) # (!ifid_ifinstr_o_21 & (((\Mux14~6_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux14~8_combout ),
	.datac(\Mux14~6_combout ),
	.datad(\Mux14~1_combout ),
	.cin(gnd),
	.combout(Mux14),
	.cout());
// synopsys translate_off
defparam \Mux14~9 .lut_mask = 16'hDAD0;
defparam \Mux14~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N2
cycloneive_lcell_comb \Mux14~19 (
// Equation(s):
// Mux141 = (ifid_ifinstr_o_24 & ((\Mux14~16_combout  & ((\Mux14~18_combout ))) # (!\Mux14~16_combout  & (\Mux14~11_combout )))) # (!ifid_ifinstr_o_24 & (\Mux14~16_combout ))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux14~16_combout ),
	.datac(\Mux14~11_combout ),
	.datad(\Mux14~18_combout ),
	.cin(gnd),
	.combout(Mux141),
	.cout());
// synopsys translate_off
defparam \Mux14~19 .lut_mask = 16'hEC64;
defparam \Mux14~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N20
cycloneive_lcell_comb \Mux32~9 (
// Equation(s):
// Mux321 = (ifid_ifinstr_o_16 & ((\Mux32~6_combout  & ((\Mux32~8_combout ))) # (!\Mux32~6_combout  & (\Mux32~1_combout )))) # (!ifid_ifinstr_o_16 & (((\Mux32~6_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux32~1_combout ),
	.datac(\Mux32~6_combout ),
	.datad(\Mux32~8_combout ),
	.cin(gnd),
	.combout(Mux321),
	.cout());
// synopsys translate_off
defparam \Mux32~9 .lut_mask = 16'hF858;
defparam \Mux32~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N26
cycloneive_lcell_comb \Mux32~19 (
// Equation(s):
// Mux322 = (ifid_ifinstr_o_18 & ((\Mux32~16_combout  & (\Mux32~18_combout )) # (!\Mux32~16_combout  & ((\Mux32~11_combout ))))) # (!ifid_ifinstr_o_18 & (((\Mux32~16_combout ))))

	.dataa(\Mux32~18_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Mux32~11_combout ),
	.datad(\Mux32~16_combout ),
	.cin(gnd),
	.combout(Mux322),
	.cout());
// synopsys translate_off
defparam \Mux32~19 .lut_mask = 16'hBBC0;
defparam \Mux32~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N12
cycloneive_lcell_comb \Mux47~9 (
// Equation(s):
// Mux47 = (\Mux47~6_combout  & ((\Mux47~8_combout ) # ((!ifid_ifinstr_o_16)))) # (!\Mux47~6_combout  & (((ifid_ifinstr_o_16 & \Mux47~1_combout ))))

	.dataa(\Mux47~6_combout ),
	.datab(\Mux47~8_combout ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux47~1_combout ),
	.cin(gnd),
	.combout(Mux47),
	.cout());
// synopsys translate_off
defparam \Mux47~9 .lut_mask = 16'hDA8A;
defparam \Mux47~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N30
cycloneive_lcell_comb \Mux47~19 (
// Equation(s):
// Mux471 = (ifid_ifinstr_o_19 & ((\Mux47~16_combout  & (\Mux47~18_combout )) # (!\Mux47~16_combout  & ((\Mux47~11_combout ))))) # (!ifid_ifinstr_o_19 & (((\Mux47~16_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Mux47~18_combout ),
	.datac(\Mux47~11_combout ),
	.datad(\Mux47~16_combout ),
	.cin(gnd),
	.combout(Mux471),
	.cout());
// synopsys translate_off
defparam \Mux47~19 .lut_mask = 16'hDDA0;
defparam \Mux47~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N16
cycloneive_lcell_comb \Mux46~9 (
// Equation(s):
// Mux46 = (ifid_ifinstr_o_16 & ((\Mux46~6_combout  & (\Mux46~8_combout )) # (!\Mux46~6_combout  & ((\Mux46~1_combout ))))) # (!ifid_ifinstr_o_16 & (((\Mux46~6_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux46~8_combout ),
	.datac(\Mux46~1_combout ),
	.datad(\Mux46~6_combout ),
	.cin(gnd),
	.combout(Mux46),
	.cout());
// synopsys translate_off
defparam \Mux46~9 .lut_mask = 16'hDDA0;
defparam \Mux46~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N30
cycloneive_lcell_comb \Mux46~19 (
// Equation(s):
// Mux461 = (\Mux46~16_combout  & ((\Mux46~18_combout ) # ((!ifid_ifinstr_o_18)))) # (!\Mux46~16_combout  & (((\Mux46~11_combout  & ifid_ifinstr_o_18))))

	.dataa(\Mux46~18_combout ),
	.datab(\Mux46~16_combout ),
	.datac(\Mux46~11_combout ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(Mux461),
	.cout());
// synopsys translate_off
defparam \Mux46~19 .lut_mask = 16'hB8CC;
defparam \Mux46~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N28
cycloneive_lcell_comb \Mux45~9 (
// Equation(s):
// Mux45 = (\Mux45~6_combout  & (((\Mux45~8_combout )) # (!ifid_ifinstr_o_16))) # (!\Mux45~6_combout  & (ifid_ifinstr_o_16 & ((\Mux45~1_combout ))))

	.dataa(\Mux45~6_combout ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux45~8_combout ),
	.datad(\Mux45~1_combout ),
	.cin(gnd),
	.combout(Mux45),
	.cout());
// synopsys translate_off
defparam \Mux45~9 .lut_mask = 16'hE6A2;
defparam \Mux45~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N12
cycloneive_lcell_comb \Mux45~19 (
// Equation(s):
// Mux451 = (ifid_ifinstr_o_19 & ((\Mux45~16_combout  & ((\Mux45~18_combout ))) # (!\Mux45~16_combout  & (\Mux45~11_combout )))) # (!ifid_ifinstr_o_19 & (((\Mux45~16_combout ))))

	.dataa(\Mux45~11_combout ),
	.datab(\Mux45~18_combout ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux45~16_combout ),
	.cin(gnd),
	.combout(Mux451),
	.cout());
// synopsys translate_off
defparam \Mux45~19 .lut_mask = 16'hCFA0;
defparam \Mux45~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N4
cycloneive_lcell_comb \Mux44~9 (
// Equation(s):
// Mux44 = (ifid_ifinstr_o_16 & ((\Mux44~6_combout  & ((\Mux44~8_combout ))) # (!\Mux44~6_combout  & (\Mux44~1_combout )))) # (!ifid_ifinstr_o_16 & (((\Mux44~6_combout ))))

	.dataa(\Mux44~1_combout ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux44~8_combout ),
	.datad(\Mux44~6_combout ),
	.cin(gnd),
	.combout(Mux44),
	.cout());
// synopsys translate_off
defparam \Mux44~9 .lut_mask = 16'hF388;
defparam \Mux44~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N16
cycloneive_lcell_comb \Mux44~19 (
// Equation(s):
// Mux441 = (ifid_ifinstr_o_18 & ((\Mux44~16_combout  & (\Mux44~18_combout )) # (!\Mux44~16_combout  & ((\Mux44~11_combout ))))) # (!ifid_ifinstr_o_18 & (\Mux44~16_combout ))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux44~16_combout ),
	.datac(\Mux44~18_combout ),
	.datad(\Mux44~11_combout ),
	.cin(gnd),
	.combout(Mux441),
	.cout());
// synopsys translate_off
defparam \Mux44~19 .lut_mask = 16'hE6C4;
defparam \Mux44~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N6
cycloneive_lcell_comb \Mux43~9 (
// Equation(s):
// Mux43 = (\Mux43~6_combout  & ((\Mux43~8_combout ) # ((!ifid_ifinstr_o_16)))) # (!\Mux43~6_combout  & (((\Mux43~1_combout  & ifid_ifinstr_o_16))))

	.dataa(\Mux43~8_combout ),
	.datab(\Mux43~1_combout ),
	.datac(\Mux43~6_combout ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(Mux43),
	.cout());
// synopsys translate_off
defparam \Mux43~9 .lut_mask = 16'hACF0;
defparam \Mux43~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N30
cycloneive_lcell_comb \Mux43~19 (
// Equation(s):
// Mux431 = (ifid_ifinstr_o_19 & ((\Mux43~16_combout  & (\Mux43~18_combout )) # (!\Mux43~16_combout  & ((\Mux43~11_combout ))))) # (!ifid_ifinstr_o_19 & (((\Mux43~16_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Mux43~18_combout ),
	.datac(\Mux43~11_combout ),
	.datad(\Mux43~16_combout ),
	.cin(gnd),
	.combout(Mux431),
	.cout());
// synopsys translate_off
defparam \Mux43~19 .lut_mask = 16'hDDA0;
defparam \Mux43~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N22
cycloneive_lcell_comb \Mux42~9 (
// Equation(s):
// Mux42 = (ifid_ifinstr_o_16 & ((\Mux42~6_combout  & (\Mux42~8_combout )) # (!\Mux42~6_combout  & ((\Mux42~1_combout ))))) # (!ifid_ifinstr_o_16 & (((\Mux42~6_combout ))))

	.dataa(\Mux42~8_combout ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux42~1_combout ),
	.datad(\Mux42~6_combout ),
	.cin(gnd),
	.combout(Mux42),
	.cout());
// synopsys translate_off
defparam \Mux42~9 .lut_mask = 16'hBBC0;
defparam \Mux42~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N0
cycloneive_lcell_comb \Mux42~19 (
// Equation(s):
// Mux421 = (ifid_ifinstr_o_18 & ((\Mux42~16_combout  & (\Mux42~18_combout )) # (!\Mux42~16_combout  & ((\Mux42~11_combout ))))) # (!ifid_ifinstr_o_18 & (((\Mux42~16_combout ))))

	.dataa(\Mux42~18_combout ),
	.datab(\Mux42~11_combout ),
	.datac(ifid_ifinstr_o_18),
	.datad(\Mux42~16_combout ),
	.cin(gnd),
	.combout(Mux421),
	.cout());
// synopsys translate_off
defparam \Mux42~19 .lut_mask = 16'hAFC0;
defparam \Mux42~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N30
cycloneive_lcell_comb \Mux41~9 (
// Equation(s):
// Mux411 = (\Mux41~6_combout  & ((\Mux41~8_combout ) # ((!ifid_ifinstr_o_16)))) # (!\Mux41~6_combout  & (((\Mux41~1_combout  & ifid_ifinstr_o_16))))

	.dataa(\Mux41~6_combout ),
	.datab(\Mux41~8_combout ),
	.datac(\Mux41~1_combout ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(Mux411),
	.cout());
// synopsys translate_off
defparam \Mux41~9 .lut_mask = 16'hD8AA;
defparam \Mux41~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N16
cycloneive_lcell_comb \Mux41~19 (
// Equation(s):
// Mux412 = (\Mux41~16_combout  & (((\Mux41~18_combout ) # (!ifid_ifinstr_o_19)))) # (!\Mux41~16_combout  & (\Mux41~11_combout  & ((ifid_ifinstr_o_19))))

	.dataa(\Mux41~16_combout ),
	.datab(\Mux41~11_combout ),
	.datac(\Mux41~18_combout ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(Mux412),
	.cout());
// synopsys translate_off
defparam \Mux41~19 .lut_mask = 16'hE4AA;
defparam \Mux41~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N0
cycloneive_lcell_comb \Mux40~9 (
// Equation(s):
// Mux40 = (\Mux40~6_combout  & (((\Mux40~8_combout ) # (!ifid_ifinstr_o_16)))) # (!\Mux40~6_combout  & (\Mux40~1_combout  & ((ifid_ifinstr_o_16))))

	.dataa(\Mux40~1_combout ),
	.datab(\Mux40~8_combout ),
	.datac(\Mux40~6_combout ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(Mux40),
	.cout());
// synopsys translate_off
defparam \Mux40~9 .lut_mask = 16'hCAF0;
defparam \Mux40~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N16
cycloneive_lcell_comb \Mux40~19 (
// Equation(s):
// Mux401 = (ifid_ifinstr_o_18 & ((\Mux40~16_combout  & ((\Mux40~18_combout ))) # (!\Mux40~16_combout  & (\Mux40~11_combout )))) # (!ifid_ifinstr_o_18 & (((\Mux40~16_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux40~11_combout ),
	.datac(\Mux40~16_combout ),
	.datad(\Mux40~18_combout ),
	.cin(gnd),
	.combout(Mux401),
	.cout());
// synopsys translate_off
defparam \Mux40~19 .lut_mask = 16'hF858;
defparam \Mux40~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N6
cycloneive_lcell_comb \Mux39~9 (
// Equation(s):
// Mux39 = (\Mux39~6_combout  & ((\Mux39~8_combout ) # ((!ifid_ifinstr_o_16)))) # (!\Mux39~6_combout  & (((\Mux39~1_combout  & ifid_ifinstr_o_16))))

	.dataa(\Mux39~8_combout ),
	.datab(\Mux39~6_combout ),
	.datac(\Mux39~1_combout ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(Mux39),
	.cout());
// synopsys translate_off
defparam \Mux39~9 .lut_mask = 16'hB8CC;
defparam \Mux39~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N2
cycloneive_lcell_comb \Mux39~19 (
// Equation(s):
// Mux391 = (\Mux39~16_combout  & ((\Mux39~18_combout ) # ((!ifid_ifinstr_o_19)))) # (!\Mux39~16_combout  & (((ifid_ifinstr_o_19 & \Mux39~11_combout ))))

	.dataa(\Mux39~18_combout ),
	.datab(\Mux39~16_combout ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux39~11_combout ),
	.cin(gnd),
	.combout(Mux391),
	.cout());
// synopsys translate_off
defparam \Mux39~19 .lut_mask = 16'hBC8C;
defparam \Mux39~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N4
cycloneive_lcell_comb \Mux38~9 (
// Equation(s):
// Mux38 = (\Mux38~6_combout  & ((\Mux38~8_combout ) # ((!ifid_ifinstr_o_16)))) # (!\Mux38~6_combout  & (((ifid_ifinstr_o_16 & \Mux38~1_combout ))))

	.dataa(\Mux38~8_combout ),
	.datab(\Mux38~6_combout ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux38~1_combout ),
	.cin(gnd),
	.combout(Mux38),
	.cout());
// synopsys translate_off
defparam \Mux38~9 .lut_mask = 16'hBC8C;
defparam \Mux38~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N24
cycloneive_lcell_comb \Mux38~19 (
// Equation(s):
// Mux381 = (ifid_ifinstr_o_18 & ((\Mux38~16_combout  & (\Mux38~18_combout )) # (!\Mux38~16_combout  & ((\Mux38~11_combout ))))) # (!ifid_ifinstr_o_18 & (((\Mux38~16_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux38~18_combout ),
	.datac(\Mux38~11_combout ),
	.datad(\Mux38~16_combout ),
	.cin(gnd),
	.combout(Mux381),
	.cout());
// synopsys translate_off
defparam \Mux38~19 .lut_mask = 16'hDDA0;
defparam \Mux38~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N28
cycloneive_lcell_comb \Mux37~9 (
// Equation(s):
// Mux37 = (ifid_ifinstr_o_16 & ((\Mux37~6_combout  & ((\Mux37~8_combout ))) # (!\Mux37~6_combout  & (\Mux37~1_combout )))) # (!ifid_ifinstr_o_16 & (((\Mux37~6_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux37~1_combout ),
	.datac(\Mux37~8_combout ),
	.datad(\Mux37~6_combout ),
	.cin(gnd),
	.combout(Mux37),
	.cout());
// synopsys translate_off
defparam \Mux37~9 .lut_mask = 16'hF588;
defparam \Mux37~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N8
cycloneive_lcell_comb \Mux37~19 (
// Equation(s):
// Mux371 = (\Mux37~16_combout  & (((\Mux37~18_combout ) # (!ifid_ifinstr_o_19)))) # (!\Mux37~16_combout  & (\Mux37~11_combout  & (ifid_ifinstr_o_19)))

	.dataa(\Mux37~16_combout ),
	.datab(\Mux37~11_combout ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux37~18_combout ),
	.cin(gnd),
	.combout(Mux371),
	.cout());
// synopsys translate_off
defparam \Mux37~19 .lut_mask = 16'hEA4A;
defparam \Mux37~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N20
cycloneive_lcell_comb \Mux58~9 (
// Equation(s):
// Mux58 = (ifid_ifinstr_o_16 & ((\Mux58~6_combout  & (\Mux58~8_combout )) # (!\Mux58~6_combout  & ((\Mux58~1_combout ))))) # (!ifid_ifinstr_o_16 & (((\Mux58~6_combout ))))

	.dataa(\Mux58~8_combout ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux58~1_combout ),
	.datad(\Mux58~6_combout ),
	.cin(gnd),
	.combout(Mux58),
	.cout());
// synopsys translate_off
defparam \Mux58~9 .lut_mask = 16'hBBC0;
defparam \Mux58~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N26
cycloneive_lcell_comb \Mux58~19 (
// Equation(s):
// Mux581 = (ifid_ifinstr_o_18 & ((\Mux58~16_combout  & ((\Mux58~18_combout ))) # (!\Mux58~16_combout  & (\Mux58~11_combout )))) # (!ifid_ifinstr_o_18 & (((\Mux58~16_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux58~11_combout ),
	.datac(\Mux58~18_combout ),
	.datad(\Mux58~16_combout ),
	.cin(gnd),
	.combout(Mux581),
	.cout());
// synopsys translate_off
defparam \Mux58~19 .lut_mask = 16'hF588;
defparam \Mux58~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N0
cycloneive_lcell_comb \Mux57~9 (
// Equation(s):
// Mux57 = (ifid_ifinstr_o_16 & ((\Mux57~6_combout  & (\Mux57~8_combout )) # (!\Mux57~6_combout  & ((\Mux57~1_combout ))))) # (!ifid_ifinstr_o_16 & (((\Mux57~6_combout ))))

	.dataa(\Mux57~8_combout ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux57~1_combout ),
	.datad(\Mux57~6_combout ),
	.cin(gnd),
	.combout(Mux57),
	.cout());
// synopsys translate_off
defparam \Mux57~9 .lut_mask = 16'hBBC0;
defparam \Mux57~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N22
cycloneive_lcell_comb \Mux57~19 (
// Equation(s):
// Mux571 = (ifid_ifinstr_o_19 & ((\Mux57~16_combout  & ((\Mux57~18_combout ))) # (!\Mux57~16_combout  & (\Mux57~11_combout )))) # (!ifid_ifinstr_o_19 & (((\Mux57~16_combout ))))

	.dataa(\Mux57~11_combout ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Mux57~18_combout ),
	.datad(\Mux57~16_combout ),
	.cin(gnd),
	.combout(Mux571),
	.cout());
// synopsys translate_off
defparam \Mux57~19 .lut_mask = 16'hF388;
defparam \Mux57~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N10
cycloneive_lcell_comb \Mux56~9 (
// Equation(s):
// Mux56 = (\Mux56~6_combout  & (((\Mux56~8_combout )) # (!ifid_ifinstr_o_16))) # (!\Mux56~6_combout  & (ifid_ifinstr_o_16 & (\Mux56~1_combout )))

	.dataa(\Mux56~6_combout ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux56~1_combout ),
	.datad(\Mux56~8_combout ),
	.cin(gnd),
	.combout(Mux56),
	.cout());
// synopsys translate_off
defparam \Mux56~9 .lut_mask = 16'hEA62;
defparam \Mux56~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N22
cycloneive_lcell_comb \Mux56~19 (
// Equation(s):
// Mux561 = (ifid_ifinstr_o_18 & ((\Mux56~16_combout  & ((\Mux56~18_combout ))) # (!\Mux56~16_combout  & (\Mux56~11_combout )))) # (!ifid_ifinstr_o_18 & (((\Mux56~16_combout ))))

	.dataa(\Mux56~11_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Mux56~18_combout ),
	.datad(\Mux56~16_combout ),
	.cin(gnd),
	.combout(Mux561),
	.cout());
// synopsys translate_off
defparam \Mux56~19 .lut_mask = 16'hF388;
defparam \Mux56~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N18
cycloneive_lcell_comb \Mux55~9 (
// Equation(s):
// Mux55 = (ifid_ifinstr_o_16 & ((\Mux55~6_combout  & (\Mux55~8_combout )) # (!\Mux55~6_combout  & ((\Mux55~1_combout ))))) # (!ifid_ifinstr_o_16 & (((\Mux55~6_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux55~8_combout ),
	.datac(\Mux55~1_combout ),
	.datad(\Mux55~6_combout ),
	.cin(gnd),
	.combout(Mux55),
	.cout());
// synopsys translate_off
defparam \Mux55~9 .lut_mask = 16'hDDA0;
defparam \Mux55~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N0
cycloneive_lcell_comb \Mux55~19 (
// Equation(s):
// Mux551 = (ifid_ifinstr_o_19 & ((\Mux55~16_combout  & (\Mux55~18_combout )) # (!\Mux55~16_combout  & ((\Mux55~11_combout ))))) # (!ifid_ifinstr_o_19 & (((\Mux55~16_combout ))))

	.dataa(\Mux55~18_combout ),
	.datab(\Mux55~11_combout ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux55~16_combout ),
	.cin(gnd),
	.combout(Mux551),
	.cout());
// synopsys translate_off
defparam \Mux55~19 .lut_mask = 16'hAFC0;
defparam \Mux55~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N30
cycloneive_lcell_comb \Mux36~9 (
// Equation(s):
// Mux36 = (ifid_ifinstr_o_16 & ((\Mux36~6_combout  & (\Mux36~8_combout )) # (!\Mux36~6_combout  & ((\Mux36~1_combout ))))) # (!ifid_ifinstr_o_16 & (((\Mux36~6_combout ))))

	.dataa(\Mux36~8_combout ),
	.datab(\Mux36~1_combout ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux36~6_combout ),
	.cin(gnd),
	.combout(Mux36),
	.cout());
// synopsys translate_off
defparam \Mux36~9 .lut_mask = 16'hAFC0;
defparam \Mux36~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N10
cycloneive_lcell_comb \Mux36~19 (
// Equation(s):
// Mux361 = (ifid_ifinstr_o_18 & ((\Mux36~16_combout  & (\Mux36~18_combout )) # (!\Mux36~16_combout  & ((\Mux36~11_combout ))))) # (!ifid_ifinstr_o_18 & (((\Mux36~16_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux36~18_combout ),
	.datac(\Mux36~11_combout ),
	.datad(\Mux36~16_combout ),
	.cin(gnd),
	.combout(Mux361),
	.cout());
// synopsys translate_off
defparam \Mux36~19 .lut_mask = 16'hDDA0;
defparam \Mux36~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N0
cycloneive_lcell_comb \Mux35~9 (
// Equation(s):
// Mux35 = (ifid_ifinstr_o_16 & ((\Mux35~6_combout  & ((\Mux35~8_combout ))) # (!\Mux35~6_combout  & (\Mux35~1_combout )))) # (!ifid_ifinstr_o_16 & (((\Mux35~6_combout ))))

	.dataa(\Mux35~1_combout ),
	.datab(\Mux35~8_combout ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux35~6_combout ),
	.cin(gnd),
	.combout(Mux35),
	.cout());
// synopsys translate_off
defparam \Mux35~9 .lut_mask = 16'hCFA0;
defparam \Mux35~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N24
cycloneive_lcell_comb \Mux35~19 (
// Equation(s):
// Mux351 = (ifid_ifinstr_o_19 & ((\Mux35~16_combout  & (\Mux35~18_combout )) # (!\Mux35~16_combout  & ((\Mux35~11_combout ))))) # (!ifid_ifinstr_o_19 & (((\Mux35~16_combout ))))

	.dataa(\Mux35~18_combout ),
	.datab(\Mux35~11_combout ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux35~16_combout ),
	.cin(gnd),
	.combout(Mux351),
	.cout());
// synopsys translate_off
defparam \Mux35~19 .lut_mask = 16'hAFC0;
defparam \Mux35~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N10
cycloneive_lcell_comb \Mux34~9 (
// Equation(s):
// Mux34 = (ifid_ifinstr_o_16 & ((\Mux34~6_combout  & (\Mux34~8_combout )) # (!\Mux34~6_combout  & ((\Mux34~1_combout ))))) # (!ifid_ifinstr_o_16 & (((\Mux34~6_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux34~8_combout ),
	.datac(\Mux34~1_combout ),
	.datad(\Mux34~6_combout ),
	.cin(gnd),
	.combout(Mux34),
	.cout());
// synopsys translate_off
defparam \Mux34~9 .lut_mask = 16'hDDA0;
defparam \Mux34~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N18
cycloneive_lcell_comb \Mux34~19 (
// Equation(s):
// Mux341 = (ifid_ifinstr_o_18 & ((\Mux34~16_combout  & ((\Mux34~18_combout ))) # (!\Mux34~16_combout  & (\Mux34~11_combout )))) # (!ifid_ifinstr_o_18 & (((\Mux34~16_combout ))))

	.dataa(\Mux34~11_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Mux34~16_combout ),
	.datad(\Mux34~18_combout ),
	.cin(gnd),
	.combout(Mux341),
	.cout());
// synopsys translate_off
defparam \Mux34~19 .lut_mask = 16'hF838;
defparam \Mux34~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N4
cycloneive_lcell_comb \Mux33~9 (
// Equation(s):
// Mux33 = (ifid_ifinstr_o_16 & ((\Mux33~6_combout  & (\Mux33~8_combout )) # (!\Mux33~6_combout  & ((\Mux33~1_combout ))))) # (!ifid_ifinstr_o_16 & (((\Mux33~6_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux33~8_combout ),
	.datac(\Mux33~6_combout ),
	.datad(\Mux33~1_combout ),
	.cin(gnd),
	.combout(Mux33),
	.cout());
// synopsys translate_off
defparam \Mux33~9 .lut_mask = 16'hDAD0;
defparam \Mux33~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N24
cycloneive_lcell_comb \Mux33~19 (
// Equation(s):
// Mux331 = (ifid_ifinstr_o_19 & ((\Mux33~16_combout  & (\Mux33~18_combout )) # (!\Mux33~16_combout  & ((\Mux33~11_combout ))))) # (!ifid_ifinstr_o_19 & (((\Mux33~16_combout ))))

	.dataa(\Mux33~18_combout ),
	.datab(\Mux33~11_combout ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux33~16_combout ),
	.cin(gnd),
	.combout(Mux331),
	.cout());
// synopsys translate_off
defparam \Mux33~19 .lut_mask = 16'hAFC0;
defparam \Mux33~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N26
cycloneive_lcell_comb \Mux54~9 (
// Equation(s):
// Mux54 = (ifid_ifinstr_o_16 & ((\Mux54~6_combout  & (\Mux54~8_combout )) # (!\Mux54~6_combout  & ((\Mux54~1_combout ))))) # (!ifid_ifinstr_o_16 & (((\Mux54~6_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux54~8_combout ),
	.datac(\Mux54~1_combout ),
	.datad(\Mux54~6_combout ),
	.cin(gnd),
	.combout(Mux54),
	.cout());
// synopsys translate_off
defparam \Mux54~9 .lut_mask = 16'hDDA0;
defparam \Mux54~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N26
cycloneive_lcell_comb \Mux54~19 (
// Equation(s):
// Mux541 = (ifid_ifinstr_o_18 & ((\Mux54~16_combout  & ((\Mux54~18_combout ))) # (!\Mux54~16_combout  & (\Mux54~11_combout )))) # (!ifid_ifinstr_o_18 & (((\Mux54~16_combout ))))

	.dataa(\Mux54~11_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Mux54~18_combout ),
	.datad(\Mux54~16_combout ),
	.cin(gnd),
	.combout(Mux541),
	.cout());
// synopsys translate_off
defparam \Mux54~19 .lut_mask = 16'hF388;
defparam \Mux54~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N28
cycloneive_lcell_comb \Mux49~9 (
// Equation(s):
// Mux49 = (ifid_ifinstr_o_16 & ((\Mux49~6_combout  & (\Mux49~8_combout )) # (!\Mux49~6_combout  & ((\Mux49~1_combout ))))) # (!ifid_ifinstr_o_16 & (((\Mux49~6_combout ))))

	.dataa(\Mux49~8_combout ),
	.datab(\Mux49~1_combout ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux49~6_combout ),
	.cin(gnd),
	.combout(Mux49),
	.cout());
// synopsys translate_off
defparam \Mux49~9 .lut_mask = 16'hAFC0;
defparam \Mux49~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N18
cycloneive_lcell_comb \Mux49~19 (
// Equation(s):
// Mux491 = (\Mux49~16_combout  & (((\Mux49~18_combout )) # (!ifid_ifinstr_o_19))) # (!\Mux49~16_combout  & (ifid_ifinstr_o_19 & (\Mux49~11_combout )))

	.dataa(\Mux49~16_combout ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Mux49~11_combout ),
	.datad(\Mux49~18_combout ),
	.cin(gnd),
	.combout(Mux491),
	.cout());
// synopsys translate_off
defparam \Mux49~19 .lut_mask = 16'hEA62;
defparam \Mux49~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N20
cycloneive_lcell_comb \Mux48~9 (
// Equation(s):
// Mux48 = (ifid_ifinstr_o_16 & ((\Mux48~6_combout  & (\Mux48~8_combout )) # (!\Mux48~6_combout  & ((\Mux48~1_combout ))))) # (!ifid_ifinstr_o_16 & (((\Mux48~6_combout ))))

	.dataa(\Mux48~8_combout ),
	.datab(\Mux48~1_combout ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux48~6_combout ),
	.cin(gnd),
	.combout(Mux48),
	.cout());
// synopsys translate_off
defparam \Mux48~9 .lut_mask = 16'hAFC0;
defparam \Mux48~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N16
cycloneive_lcell_comb \Mux48~19 (
// Equation(s):
// Mux481 = (\Mux48~16_combout  & ((\Mux48~18_combout ) # ((!ifid_ifinstr_o_18)))) # (!\Mux48~16_combout  & (((\Mux48~11_combout  & ifid_ifinstr_o_18))))

	.dataa(\Mux48~16_combout ),
	.datab(\Mux48~18_combout ),
	.datac(\Mux48~11_combout ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(Mux481),
	.cout());
// synopsys translate_off
defparam \Mux48~19 .lut_mask = 16'hD8AA;
defparam \Mux48~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N2
cycloneive_lcell_comb \Mux53~9 (
// Equation(s):
// Mux53 = (\Mux53~6_combout  & ((\Mux53~8_combout ) # ((!ifid_ifinstr_o_16)))) # (!\Mux53~6_combout  & (((ifid_ifinstr_o_16 & \Mux53~1_combout ))))

	.dataa(\Mux53~8_combout ),
	.datab(\Mux53~6_combout ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux53~1_combout ),
	.cin(gnd),
	.combout(Mux53),
	.cout());
// synopsys translate_off
defparam \Mux53~9 .lut_mask = 16'hBC8C;
defparam \Mux53~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N26
cycloneive_lcell_comb \Mux53~19 (
// Equation(s):
// Mux531 = (ifid_ifinstr_o_19 & ((\Mux53~16_combout  & (\Mux53~18_combout )) # (!\Mux53~16_combout  & ((\Mux53~11_combout ))))) # (!ifid_ifinstr_o_19 & (((\Mux53~16_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Mux53~18_combout ),
	.datac(\Mux53~16_combout ),
	.datad(\Mux53~11_combout ),
	.cin(gnd),
	.combout(Mux531),
	.cout());
// synopsys translate_off
defparam \Mux53~19 .lut_mask = 16'hDAD0;
defparam \Mux53~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N20
cycloneive_lcell_comb \Mux52~9 (
// Equation(s):
// Mux52 = (\Mux52~6_combout  & ((\Mux52~8_combout ) # ((!ifid_ifinstr_o_16)))) # (!\Mux52~6_combout  & (((ifid_ifinstr_o_16 & \Mux52~1_combout ))))

	.dataa(\Mux52~8_combout ),
	.datab(\Mux52~6_combout ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux52~1_combout ),
	.cin(gnd),
	.combout(Mux52),
	.cout());
// synopsys translate_off
defparam \Mux52~9 .lut_mask = 16'hBC8C;
defparam \Mux52~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N26
cycloneive_lcell_comb \Mux52~19 (
// Equation(s):
// Mux521 = (ifid_ifinstr_o_18 & ((\Mux52~16_combout  & ((\Mux52~18_combout ))) # (!\Mux52~16_combout  & (\Mux52~11_combout )))) # (!ifid_ifinstr_o_18 & (\Mux52~16_combout ))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux52~16_combout ),
	.datac(\Mux52~11_combout ),
	.datad(\Mux52~18_combout ),
	.cin(gnd),
	.combout(Mux521),
	.cout());
// synopsys translate_off
defparam \Mux52~19 .lut_mask = 16'hEC64;
defparam \Mux52~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N6
cycloneive_lcell_comb \Mux51~9 (
// Equation(s):
// Mux511 = (\Mux51~6_combout  & (((\Mux51~8_combout ) # (!ifid_ifinstr_o_16)))) # (!\Mux51~6_combout  & (\Mux51~1_combout  & ((ifid_ifinstr_o_16))))

	.dataa(\Mux51~1_combout ),
	.datab(\Mux51~8_combout ),
	.datac(\Mux51~6_combout ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(Mux511),
	.cout());
// synopsys translate_off
defparam \Mux51~9 .lut_mask = 16'hCAF0;
defparam \Mux51~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N6
cycloneive_lcell_comb \Mux51~19 (
// Equation(s):
// Mux512 = (ifid_ifinstr_o_19 & ((\Mux51~16_combout  & (\Mux51~18_combout )) # (!\Mux51~16_combout  & ((\Mux51~11_combout ))))) # (!ifid_ifinstr_o_19 & (((\Mux51~16_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Mux51~18_combout ),
	.datac(\Mux51~11_combout ),
	.datad(\Mux51~16_combout ),
	.cin(gnd),
	.combout(Mux512),
	.cout());
// synopsys translate_off
defparam \Mux51~19 .lut_mask = 16'hDDA0;
defparam \Mux51~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N16
cycloneive_lcell_comb \Mux50~9 (
// Equation(s):
// Mux50 = (ifid_ifinstr_o_16 & ((\Mux50~6_combout  & ((\Mux50~8_combout ))) # (!\Mux50~6_combout  & (\Mux50~1_combout )))) # (!ifid_ifinstr_o_16 & (((\Mux50~6_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux50~1_combout ),
	.datac(\Mux50~8_combout ),
	.datad(\Mux50~6_combout ),
	.cin(gnd),
	.combout(Mux50),
	.cout());
// synopsys translate_off
defparam \Mux50~9 .lut_mask = 16'hF588;
defparam \Mux50~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N26
cycloneive_lcell_comb \Mux50~19 (
// Equation(s):
// Mux501 = (\Mux50~16_combout  & (((\Mux50~18_combout )) # (!ifid_ifinstr_o_18))) # (!\Mux50~16_combout  & (ifid_ifinstr_o_18 & ((\Mux50~11_combout ))))

	.dataa(\Mux50~16_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Mux50~18_combout ),
	.datad(\Mux50~11_combout ),
	.cin(gnd),
	.combout(Mux501),
	.cout());
// synopsys translate_off
defparam \Mux50~19 .lut_mask = 16'hE6A2;
defparam \Mux50~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N10
cycloneive_lcell_comb \Reg[21][1]~feeder (
// Equation(s):
// \Reg[21][1]~feeder_combout  = \wdat~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat),
	.cin(gnd),
	.combout(\Reg[21][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[21][1]~feeder .lut_mask = 16'hFF00;
defparam \Reg[21][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N26
cycloneive_lcell_comb \Decoder0~0 (
// Equation(s):
// \Decoder0~0_combout  = (\rwWB~4_combout  & (\rwWB~1_combout  & memwb_ifregWEN_o))

	.dataa(rwWB4),
	.datab(rwWB1),
	.datac(memwb_ifregWEN_o),
	.datad(gnd),
	.cin(gnd),
	.combout(\Decoder0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~0 .lut_mask = 16'h8080;
defparam \Decoder0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N22
cycloneive_lcell_comb \Decoder0~1 (
// Equation(s):
// \Decoder0~1_combout  = (!\rwWB~0_combout  & (\rwWB~3_combout  & (!\rwWB~2_combout  & \Decoder0~0_combout )))

	.dataa(rwWB),
	.datab(rwWB3),
	.datac(rwWB2),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~1 .lut_mask = 16'h0400;
defparam \Decoder0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N11
dffeas \Reg[21][1] (
	.clk(!CLK),
	.d(\Reg[21][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][1] .is_wysiwyg = "true";
defparam \Reg[21][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N4
cycloneive_lcell_comb \Reg[29][1]~feeder (
// Equation(s):
// \Reg[29][1]~feeder_combout  = \wdat~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat),
	.cin(gnd),
	.combout(\Reg[29][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[29][1]~feeder .lut_mask = 16'hFF00;
defparam \Reg[29][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N0
cycloneive_lcell_comb \Decoder0~4 (
// Equation(s):
// \Decoder0~4_combout  = (!\rwWB~0_combout  & (\rwWB~3_combout  & (\rwWB~2_combout  & \Decoder0~0_combout )))

	.dataa(rwWB),
	.datab(rwWB3),
	.datac(rwWB2),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~4 .lut_mask = 16'h4000;
defparam \Decoder0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N5
dffeas \Reg[29][1] (
	.clk(!CLK),
	.d(\Reg[29][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][1] .is_wysiwyg = "true";
defparam \Reg[29][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N20
cycloneive_lcell_comb \Decoder0~2 (
// Equation(s):
// \Decoder0~2_combout  = (!\rwWB~0_combout  & (!\rwWB~3_combout  & (\rwWB~2_combout  & \Decoder0~0_combout )))

	.dataa(rwWB),
	.datab(rwWB3),
	.datac(rwWB2),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~2 .lut_mask = 16'h1000;
defparam \Decoder0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N9
dffeas \Reg[25][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][1] .is_wysiwyg = "true";
defparam \Reg[25][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N26
cycloneive_lcell_comb \Decoder0~3 (
// Equation(s):
// \Decoder0~3_combout  = (!\rwWB~0_combout  & (!\rwWB~3_combout  & (!\rwWB~2_combout  & \Decoder0~0_combout )))

	.dataa(rwWB),
	.datab(rwWB3),
	.datac(rwWB2),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~3 .lut_mask = 16'h0100;
defparam \Decoder0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N31
dffeas \Reg[17][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][1] .is_wysiwyg = "true";
defparam \Reg[17][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N8
cycloneive_lcell_comb \Mux62~0 (
// Equation(s):
// \Mux62~0_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Reg[25][1]~q )) # (!ifid_ifinstr_o_19 & ((\Reg[17][1]~q )))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[25][1]~q ),
	.datad(\Reg[17][1]~q ),
	.cin(gnd),
	.combout(\Mux62~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~0 .lut_mask = 16'hD9C8;
defparam \Mux62~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N20
cycloneive_lcell_comb \Mux62~1 (
// Equation(s):
// \Mux62~1_combout  = (\Mux62~0_combout  & (((\Reg[29][1]~q ) # (!ifid_ifinstr_o_18)))) # (!\Mux62~0_combout  & (\Reg[21][1]~q  & ((ifid_ifinstr_o_18))))

	.dataa(\Reg[21][1]~q ),
	.datab(\Reg[29][1]~q ),
	.datac(\Mux62~0_combout ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux62~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~1 .lut_mask = 16'hCAF0;
defparam \Mux62~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N8
cycloneive_lcell_comb \Decoder0~5 (
// Equation(s):
// \Decoder0~5_combout  = (\rwWB~4_combout  & (!\rwWB~1_combout  & memwb_ifregWEN_o))

	.dataa(rwWB4),
	.datab(rwWB1),
	.datac(memwb_ifregWEN_o),
	.datad(gnd),
	.cin(gnd),
	.combout(\Decoder0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~5 .lut_mask = 16'h2020;
defparam \Decoder0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N18
cycloneive_lcell_comb \Decoder0~6 (
// Equation(s):
// \Decoder0~6_combout  = (!\rwWB~3_combout  & (\rwWB~2_combout  & (\rwWB~0_combout  & \Decoder0~5_combout )))

	.dataa(rwWB3),
	.datab(rwWB2),
	.datac(rwWB),
	.datad(\Decoder0~5_combout ),
	.cin(gnd),
	.combout(\Decoder0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~6 .lut_mask = 16'h4000;
defparam \Decoder0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N17
dffeas \Reg[26][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][1] .is_wysiwyg = "true";
defparam \Reg[26][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N0
cycloneive_lcell_comb \Decoder0~7 (
// Equation(s):
// \Decoder0~7_combout  = (\rwWB~3_combout  & (!\rwWB~2_combout  & (\rwWB~0_combout  & \Decoder0~5_combout )))

	.dataa(rwWB3),
	.datab(rwWB2),
	.datac(rwWB),
	.datad(\Decoder0~5_combout ),
	.cin(gnd),
	.combout(\Decoder0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~7 .lut_mask = 16'h2000;
defparam \Decoder0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N17
dffeas \Reg[22][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][1] .is_wysiwyg = "true";
defparam \Reg[22][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N2
cycloneive_lcell_comb \Decoder0~8 (
// Equation(s):
// \Decoder0~8_combout  = (!\rwWB~2_combout  & (\rwWB~0_combout  & (!\rwWB~3_combout  & \Decoder0~5_combout )))

	.dataa(rwWB2),
	.datab(rwWB),
	.datac(rwWB3),
	.datad(\Decoder0~5_combout ),
	.cin(gnd),
	.combout(\Decoder0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~8 .lut_mask = 16'h0400;
defparam \Decoder0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N5
dffeas \Reg[18][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][1] .is_wysiwyg = "true";
defparam \Reg[18][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N16
cycloneive_lcell_comb \Mux62~2 (
// Equation(s):
// \Mux62~2_combout  = (ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19) # ((\Reg[22][1]~q )))) # (!ifid_ifinstr_o_18 & (!ifid_ifinstr_o_19 & ((\Reg[18][1]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[22][1]~q ),
	.datad(\Reg[18][1]~q ),
	.cin(gnd),
	.combout(\Mux62~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~2 .lut_mask = 16'hB9A8;
defparam \Mux62~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N16
cycloneive_lcell_comb \Mux62~3 (
// Equation(s):
// \Mux62~3_combout  = (ifid_ifinstr_o_19 & ((\Mux62~2_combout  & (\Reg[30][1]~q )) # (!\Mux62~2_combout  & ((\Reg[26][1]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux62~2_combout ))))

	.dataa(\Reg[30][1]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[26][1]~q ),
	.datad(\Mux62~2_combout ),
	.cin(gnd),
	.combout(\Mux62~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~3 .lut_mask = 16'hBBC0;
defparam \Mux62~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N8
cycloneive_lcell_comb \Decoder0~11 (
// Equation(s):
// \Decoder0~11_combout  = (\rwWB~3_combout  & (!\rwWB~2_combout  & (!\rwWB~0_combout  & \Decoder0~5_combout )))

	.dataa(rwWB3),
	.datab(rwWB2),
	.datac(rwWB),
	.datad(\Decoder0~5_combout ),
	.cin(gnd),
	.combout(\Decoder0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~11 .lut_mask = 16'h0200;
defparam \Decoder0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N25
dffeas \Reg[20][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][1] .is_wysiwyg = "true";
defparam \Reg[20][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N26
cycloneive_lcell_comb \Decoder0~12 (
// Equation(s):
// \Decoder0~12_combout  = (!\rwWB~2_combout  & (!\rwWB~0_combout  & (!\rwWB~3_combout  & \Decoder0~5_combout )))

	.dataa(rwWB2),
	.datab(rwWB),
	.datac(rwWB3),
	.datad(\Decoder0~5_combout ),
	.cin(gnd),
	.combout(\Decoder0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~12 .lut_mask = 16'h0100;
defparam \Decoder0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N27
dffeas \Reg[16][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][1] .is_wysiwyg = "true";
defparam \Reg[16][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N24
cycloneive_lcell_comb \Mux62~4 (
// Equation(s):
// \Mux62~4_combout  = (ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19) # ((\Reg[20][1]~q )))) # (!ifid_ifinstr_o_18 & (!ifid_ifinstr_o_19 & ((\Reg[16][1]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[20][1]~q ),
	.datad(\Reg[16][1]~q ),
	.cin(gnd),
	.combout(\Mux62~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~4 .lut_mask = 16'hB9A8;
defparam \Mux62~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N26
cycloneive_lcell_comb \Decoder0~13 (
// Equation(s):
// \Decoder0~13_combout  = (\rwWB~3_combout  & (\rwWB~2_combout  & (!\rwWB~0_combout  & \Decoder0~5_combout )))

	.dataa(rwWB3),
	.datab(rwWB2),
	.datac(rwWB),
	.datad(\Decoder0~5_combout ),
	.cin(gnd),
	.combout(\Decoder0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~13 .lut_mask = 16'h0800;
defparam \Decoder0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N7
dffeas \Reg[28][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][1] .is_wysiwyg = "true";
defparam \Reg[28][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N4
cycloneive_lcell_comb \Reg[24][1]~feeder (
// Equation(s):
// \Reg[24][1]~feeder_combout  = \wdat~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat),
	.cin(gnd),
	.combout(\Reg[24][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[24][1]~feeder .lut_mask = 16'hFF00;
defparam \Reg[24][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N28
cycloneive_lcell_comb \Decoder0~10 (
// Equation(s):
// \Decoder0~10_combout  = (\rwWB~2_combout  & (!\rwWB~0_combout  & (!\rwWB~3_combout  & \Decoder0~5_combout )))

	.dataa(rwWB2),
	.datab(rwWB),
	.datac(rwWB3),
	.datad(\Decoder0~5_combout ),
	.cin(gnd),
	.combout(\Decoder0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~10 .lut_mask = 16'h0200;
defparam \Decoder0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N5
dffeas \Reg[24][1] (
	.clk(!CLK),
	.d(\Reg[24][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][1] .is_wysiwyg = "true";
defparam \Reg[24][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N6
cycloneive_lcell_comb \Mux62~5 (
// Equation(s):
// \Mux62~5_combout  = (ifid_ifinstr_o_19 & ((\Mux62~4_combout  & (\Reg[28][1]~q )) # (!\Mux62~4_combout  & ((\Reg[24][1]~q ))))) # (!ifid_ifinstr_o_19 & (\Mux62~4_combout ))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Mux62~4_combout ),
	.datac(\Reg[28][1]~q ),
	.datad(\Reg[24][1]~q ),
	.cin(gnd),
	.combout(\Mux62~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~5 .lut_mask = 16'hE6C4;
defparam \Mux62~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N14
cycloneive_lcell_comb \Mux62~6 (
// Equation(s):
// \Mux62~6_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Mux62~3_combout )) # (!ifid_ifinstr_o_17 & ((\Mux62~5_combout )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux62~3_combout ),
	.datad(\Mux62~5_combout ),
	.cin(gnd),
	.combout(\Mux62~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~6 .lut_mask = 16'hD9C8;
defparam \Mux62~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N10
cycloneive_lcell_comb \Decoder0~14 (
// Equation(s):
// \Decoder0~14_combout  = (\rwWB~0_combout  & (\rwWB~3_combout  & (!\rwWB~2_combout  & \Decoder0~0_combout )))

	.dataa(rwWB),
	.datab(rwWB3),
	.datac(rwWB2),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~14 .lut_mask = 16'h0800;
defparam \Decoder0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N1
dffeas \Reg[23][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][1] .is_wysiwyg = "true";
defparam \Reg[23][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N2
cycloneive_lcell_comb \Decoder0~16 (
// Equation(s):
// \Decoder0~16_combout  = (\rwWB~0_combout  & (!\rwWB~3_combout  & (!\rwWB~2_combout  & \Decoder0~0_combout )))

	.dataa(rwWB),
	.datab(rwWB3),
	.datac(rwWB2),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~16 .lut_mask = 16'h0200;
defparam \Decoder0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N11
dffeas \Reg[19][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][1] .is_wysiwyg = "true";
defparam \Reg[19][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N16
cycloneive_lcell_comb \Decoder0~15 (
// Equation(s):
// \Decoder0~15_combout  = (\rwWB~0_combout  & (!\rwWB~3_combout  & (\rwWB~2_combout  & \Decoder0~0_combout )))

	.dataa(rwWB),
	.datab(rwWB3),
	.datac(rwWB2),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~15 .lut_mask = 16'h2000;
defparam \Decoder0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N21
dffeas \Reg[27][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][1] .is_wysiwyg = "true";
defparam \Reg[27][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N10
cycloneive_lcell_comb \Mux62~7 (
// Equation(s):
// \Mux62~7_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[27][1]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[19][1]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[19][1]~q ),
	.datad(\Reg[27][1]~q ),
	.cin(gnd),
	.combout(\Mux62~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~7 .lut_mask = 16'hDC98;
defparam \Mux62~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N28
cycloneive_lcell_comb \Decoder0~17 (
// Equation(s):
// \Decoder0~17_combout  = (\rwWB~0_combout  & (\rwWB~3_combout  & (\rwWB~2_combout  & \Decoder0~0_combout )))

	.dataa(rwWB),
	.datab(rwWB3),
	.datac(rwWB2),
	.datad(\Decoder0~0_combout ),
	.cin(gnd),
	.combout(\Decoder0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~17 .lut_mask = 16'h8000;
defparam \Decoder0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N19
dffeas \Reg[31][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][1] .is_wysiwyg = "true";
defparam \Reg[31][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N18
cycloneive_lcell_comb \Mux62~8 (
// Equation(s):
// \Mux62~8_combout  = (\Mux62~7_combout  & (((\Reg[31][1]~q ) # (!ifid_ifinstr_o_18)))) # (!\Mux62~7_combout  & (\Reg[23][1]~q  & ((ifid_ifinstr_o_18))))

	.dataa(\Reg[23][1]~q ),
	.datab(\Mux62~7_combout ),
	.datac(\Reg[31][1]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux62~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~8 .lut_mask = 16'hE2CC;
defparam \Mux62~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N0
cycloneive_lcell_comb \Decoder0~36 (
// Equation(s):
// \Decoder0~36_combout  = (\Decoder0~20_combout  & (\rwWB~0_combout  & \rwWB~2_combout ))

	.dataa(\Decoder0~20_combout ),
	.datab(rwWB),
	.datac(gnd),
	.datad(rwWB2),
	.cin(gnd),
	.combout(\Decoder0~36_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~36 .lut_mask = 16'h8800;
defparam \Decoder0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N7
dffeas \Reg[15][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][1] .is_wysiwyg = "true";
defparam \Reg[15][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N30
cycloneive_lcell_comb \Decoder0~18 (
// Equation(s):
// \Decoder0~18_combout  = (!\rwWB~4_combout  & (memwb_ifregWEN_o & (!\rwWB~1_combout  & \rwWB~3_combout )))

	.dataa(rwWB4),
	.datab(memwb_ifregWEN_o),
	.datac(rwWB1),
	.datad(rwWB3),
	.cin(gnd),
	.combout(\Decoder0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~18 .lut_mask = 16'h0400;
defparam \Decoder0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N18
cycloneive_lcell_comb \Decoder0~33 (
// Equation(s):
// \Decoder0~33_combout  = (\rwWB~0_combout  & (\rwWB~2_combout  & \Decoder0~18_combout ))

	.dataa(rwWB),
	.datab(gnd),
	.datac(rwWB2),
	.datad(\Decoder0~18_combout ),
	.cin(gnd),
	.combout(\Decoder0~33_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~33 .lut_mask = 16'hA000;
defparam \Decoder0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N13
dffeas \Reg[14][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][1] .is_wysiwyg = "true";
defparam \Reg[14][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N30
cycloneive_lcell_comb \Decoder0~35 (
// Equation(s):
// \Decoder0~35_combout  = (!\rwWB~0_combout  & (\rwWB~2_combout  & \Decoder0~18_combout ))

	.dataa(rwWB),
	.datab(gnd),
	.datac(rwWB2),
	.datad(\Decoder0~18_combout ),
	.cin(gnd),
	.combout(\Decoder0~35_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~35 .lut_mask = 16'h5000;
defparam \Decoder0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y34_N5
dffeas \Reg[12][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][1] .is_wysiwyg = "true";
defparam \Reg[12][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N30
cycloneive_lcell_comb \Decoder0~20 (
// Equation(s):
// \Decoder0~20_combout  = (\rwWB~3_combout  & (memwb_ifregWEN_o & (!\rwWB~4_combout  & \rwWB~1_combout )))

	.dataa(rwWB3),
	.datab(memwb_ifregWEN_o),
	.datac(rwWB4),
	.datad(rwWB1),
	.cin(gnd),
	.combout(\Decoder0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~20 .lut_mask = 16'h0800;
defparam \Decoder0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N8
cycloneive_lcell_comb \Decoder0~34 (
// Equation(s):
// \Decoder0~34_combout  = (!\rwWB~0_combout  & (\rwWB~2_combout  & \Decoder0~20_combout ))

	.dataa(rwWB),
	.datab(gnd),
	.datac(rwWB2),
	.datad(\Decoder0~20_combout ),
	.cin(gnd),
	.combout(\Decoder0~34_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~34 .lut_mask = 16'h5000;
defparam \Decoder0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N25
dffeas \Reg[13][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][1] .is_wysiwyg = "true";
defparam \Reg[13][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N4
cycloneive_lcell_comb \Mux62~17 (
// Equation(s):
// \Mux62~17_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17) # ((\Reg[13][1]~q )))) # (!ifid_ifinstr_o_16 & (!ifid_ifinstr_o_17 & (\Reg[12][1]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[12][1]~q ),
	.datad(\Reg[13][1]~q ),
	.cin(gnd),
	.combout(\Mux62~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~17 .lut_mask = 16'hBA98;
defparam \Mux62~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N12
cycloneive_lcell_comb \Mux62~18 (
// Equation(s):
// \Mux62~18_combout  = (ifid_ifinstr_o_17 & ((\Mux62~17_combout  & (\Reg[15][1]~q )) # (!\Mux62~17_combout  & ((\Reg[14][1]~q ))))) # (!ifid_ifinstr_o_17 & (((\Mux62~17_combout ))))

	.dataa(\Reg[15][1]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[14][1]~q ),
	.datad(\Mux62~17_combout ),
	.cin(gnd),
	.combout(\Mux62~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~18 .lut_mask = 16'hBBC0;
defparam \Mux62~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N28
cycloneive_lcell_comb \Decoder0~21 (
// Equation(s):
// \Decoder0~21_combout  = (\Decoder0~20_combout  & (!\rwWB~0_combout  & !\rwWB~2_combout ))

	.dataa(\Decoder0~20_combout ),
	.datab(rwWB),
	.datac(gnd),
	.datad(rwWB2),
	.cin(gnd),
	.combout(\Decoder0~21_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~21 .lut_mask = 16'h0022;
defparam \Decoder0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N13
dffeas \Reg[5][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][1] .is_wysiwyg = "true";
defparam \Reg[5][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N12
cycloneive_lcell_comb \Mux62~10 (
// Equation(s):
// \Mux62~10_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[5][1]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[4][1]~q ))))

	.dataa(\Reg[4][1]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[5][1]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux62~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~10 .lut_mask = 16'hFC22;
defparam \Mux62~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N28
cycloneive_lcell_comb \Reg[7][1]~feeder (
// Equation(s):
// \Reg[7][1]~feeder_combout  = \wdat~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat),
	.cin(gnd),
	.combout(\Reg[7][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[7][1]~feeder .lut_mask = 16'hFF00;
defparam \Reg[7][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N12
cycloneive_lcell_comb \Decoder0~23 (
// Equation(s):
// \Decoder0~23_combout  = (\rwWB~0_combout  & (!\rwWB~2_combout  & \Decoder0~20_combout ))

	.dataa(rwWB),
	.datab(rwWB2),
	.datac(gnd),
	.datad(\Decoder0~20_combout ),
	.cin(gnd),
	.combout(\Decoder0~23_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~23 .lut_mask = 16'h2200;
defparam \Decoder0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N29
dffeas \Reg[7][1] (
	.clk(!CLK),
	.d(\Reg[7][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][1] .is_wysiwyg = "true";
defparam \Reg[7][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N10
cycloneive_lcell_comb \Reg[6][1]~feeder (
// Equation(s):
// \Reg[6][1]~feeder_combout  = \wdat~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat),
	.cin(gnd),
	.combout(\Reg[6][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[6][1]~feeder .lut_mask = 16'hFF00;
defparam \Reg[6][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N14
cycloneive_lcell_comb \Decoder0~19 (
// Equation(s):
// \Decoder0~19_combout  = (\rwWB~0_combout  & (!\rwWB~2_combout  & \Decoder0~18_combout ))

	.dataa(rwWB),
	.datab(gnd),
	.datac(rwWB2),
	.datad(\Decoder0~18_combout ),
	.cin(gnd),
	.combout(\Decoder0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~19 .lut_mask = 16'h0A00;
defparam \Decoder0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N11
dffeas \Reg[6][1] (
	.clk(!CLK),
	.d(\Reg[6][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][1] .is_wysiwyg = "true";
defparam \Reg[6][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N16
cycloneive_lcell_comb \Mux62~11 (
// Equation(s):
// \Mux62~11_combout  = (\Mux62~10_combout  & (((\Reg[7][1]~q )) # (!ifid_ifinstr_o_17))) # (!\Mux62~10_combout  & (ifid_ifinstr_o_17 & ((\Reg[6][1]~q ))))

	.dataa(\Mux62~10_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[7][1]~q ),
	.datad(\Reg[6][1]~q ),
	.cin(gnd),
	.combout(\Mux62~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~11 .lut_mask = 16'hE6A2;
defparam \Mux62~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N18
cycloneive_lcell_comb \Reg[2][1]~feeder (
// Equation(s):
// \Reg[2][1]~feeder_combout  = \wdat~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat),
	.cin(gnd),
	.combout(\Reg[2][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[2][1]~feeder .lut_mask = 16'hFF00;
defparam \Reg[2][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N26
cycloneive_lcell_comb \Decoder0~26 (
// Equation(s):
// \Decoder0~26_combout  = (!\rwWB~3_combout  & (memwb_ifregWEN_o & (!\rwWB~4_combout  & !\rwWB~1_combout )))

	.dataa(rwWB3),
	.datab(memwb_ifregWEN_o),
	.datac(rwWB4),
	.datad(rwWB1),
	.cin(gnd),
	.combout(\Decoder0~26_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~26 .lut_mask = 16'h0004;
defparam \Decoder0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N10
cycloneive_lcell_comb \Decoder0~32 (
// Equation(s):
// \Decoder0~32_combout  = (!\rwWB~2_combout  & (\Decoder0~26_combout  & \rwWB~0_combout ))

	.dataa(rwWB2),
	.datab(gnd),
	.datac(\Decoder0~26_combout ),
	.datad(rwWB),
	.cin(gnd),
	.combout(\Decoder0~32_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~32 .lut_mask = 16'h5000;
defparam \Decoder0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N19
dffeas \Reg[2][1] (
	.clk(!CLK),
	.d(\Reg[2][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][1] .is_wysiwyg = "true";
defparam \Reg[2][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N22
cycloneive_lcell_comb \Mux62~15 (
// Equation(s):
// \Mux62~15_combout  = (\Mux62~14_combout ) # ((ifid_ifinstr_o_17 & (\Reg[2][1]~q  & !ifid_ifinstr_o_16)))

	.dataa(\Mux62~14_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[2][1]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux62~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~15 .lut_mask = 16'hAAEA;
defparam \Mux62~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N18
cycloneive_lcell_comb \Decoder0~24 (
// Equation(s):
// \Decoder0~24_combout  = (!\rwWB~3_combout  & (memwb_ifregWEN_o & (!\rwWB~4_combout  & \rwWB~1_combout )))

	.dataa(rwWB3),
	.datab(memwb_ifregWEN_o),
	.datac(rwWB4),
	.datad(rwWB1),
	.cin(gnd),
	.combout(\Decoder0~24_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~24 .lut_mask = 16'h0400;
defparam \Decoder0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N16
cycloneive_lcell_comb \Decoder0~25 (
// Equation(s):
// \Decoder0~25_combout  = (\rwWB~2_combout  & (\Decoder0~24_combout  & !\rwWB~0_combout ))

	.dataa(rwWB2),
	.datab(\Decoder0~24_combout ),
	.datac(gnd),
	.datad(rwWB),
	.cin(gnd),
	.combout(\Decoder0~25_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~25 .lut_mask = 16'h0088;
defparam \Decoder0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N21
dffeas \Reg[9][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][1] .is_wysiwyg = "true";
defparam \Reg[9][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N4
cycloneive_lcell_comb \Decoder0~29 (
// Equation(s):
// \Decoder0~29_combout  = (\rwWB~2_combout  & (\Decoder0~24_combout  & \rwWB~0_combout ))

	.dataa(rwWB2),
	.datab(\Decoder0~24_combout ),
	.datac(gnd),
	.datad(rwWB),
	.cin(gnd),
	.combout(\Decoder0~29_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~29 .lut_mask = 16'h8800;
defparam \Decoder0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N15
dffeas \Reg[11][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][1] .is_wysiwyg = "true";
defparam \Reg[11][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N2
cycloneive_lcell_comb \Decoder0~28 (
// Equation(s):
// \Decoder0~28_combout  = (\rwWB~2_combout  & (\Decoder0~26_combout  & !\rwWB~0_combout ))

	.dataa(rwWB2),
	.datab(gnd),
	.datac(\Decoder0~26_combout ),
	.datad(rwWB),
	.cin(gnd),
	.combout(\Decoder0~28_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~28 .lut_mask = 16'h00A0;
defparam \Decoder0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N7
dffeas \Reg[8][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][1] .is_wysiwyg = "true";
defparam \Reg[8][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N24
cycloneive_lcell_comb \Decoder0~27 (
// Equation(s):
// \Decoder0~27_combout  = (\rwWB~2_combout  & (\Decoder0~26_combout  & \rwWB~0_combout ))

	.dataa(rwWB2),
	.datab(gnd),
	.datac(\Decoder0~26_combout ),
	.datad(rwWB),
	.cin(gnd),
	.combout(\Decoder0~27_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~27 .lut_mask = 16'hA000;
defparam \Decoder0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N17
dffeas \Reg[10][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][1] .is_wysiwyg = "true";
defparam \Reg[10][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N6
cycloneive_lcell_comb \Mux62~12 (
// Equation(s):
// \Mux62~12_combout  = (ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16) # ((\Reg[10][1]~q )))) # (!ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & (\Reg[8][1]~q )))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[8][1]~q ),
	.datad(\Reg[10][1]~q ),
	.cin(gnd),
	.combout(\Mux62~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~12 .lut_mask = 16'hBA98;
defparam \Mux62~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N14
cycloneive_lcell_comb \Mux62~13 (
// Equation(s):
// \Mux62~13_combout  = (ifid_ifinstr_o_16 & ((\Mux62~12_combout  & ((\Reg[11][1]~q ))) # (!\Mux62~12_combout  & (\Reg[9][1]~q )))) # (!ifid_ifinstr_o_16 & (((\Mux62~12_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[9][1]~q ),
	.datac(\Reg[11][1]~q ),
	.datad(\Mux62~12_combout ),
	.cin(gnd),
	.combout(\Mux62~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~13 .lut_mask = 16'hF588;
defparam \Mux62~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N24
cycloneive_lcell_comb \Mux62~16 (
// Equation(s):
// \Mux62~16_combout  = (ifid_ifinstr_o_19 & (((ifid_ifinstr_o_18) # (\Mux62~13_combout )))) # (!ifid_ifinstr_o_19 & (\Mux62~15_combout  & (!ifid_ifinstr_o_18)))

	.dataa(\Mux62~15_combout ),
	.datab(ifid_ifinstr_o_19),
	.datac(ifid_ifinstr_o_18),
	.datad(\Mux62~13_combout ),
	.cin(gnd),
	.combout(\Mux62~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~16 .lut_mask = 16'hCEC2;
defparam \Mux62~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N30
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// \Mux30~0_combout  = (ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24) # ((\Reg[21][1]~q )))) # (!ifid_ifinstr_o_23 & (!ifid_ifinstr_o_24 & (\Reg[17][1]~q )))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[17][1]~q ),
	.datad(\Reg[21][1]~q ),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'hBA98;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N4
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// \Mux30~1_combout  = (\Mux30~0_combout  & (((\Reg[29][1]~q ) # (!ifid_ifinstr_o_24)))) # (!\Mux30~0_combout  & (\Reg[25][1]~q  & (ifid_ifinstr_o_24)))

	.dataa(\Mux30~0_combout ),
	.datab(\Reg[25][1]~q ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Reg[29][1]~q ),
	.cin(gnd),
	.combout(\Mux30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'hEA4A;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N4
cycloneive_lcell_comb \Mux30~2 (
// Equation(s):
// \Mux30~2_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[26][1]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & (\Reg[18][1]~q )))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[18][1]~q ),
	.datad(\Reg[26][1]~q ),
	.cin(gnd),
	.combout(\Mux30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~2 .lut_mask = 16'hBA98;
defparam \Mux30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N22
cycloneive_lcell_comb \Decoder0~9 (
// Equation(s):
// \Decoder0~9_combout  = (\rwWB~3_combout  & (\rwWB~2_combout  & (\rwWB~0_combout  & \Decoder0~5_combout )))

	.dataa(rwWB3),
	.datab(rwWB2),
	.datac(rwWB),
	.datad(\Decoder0~5_combout ),
	.cin(gnd),
	.combout(\Decoder0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~9 .lut_mask = 16'h8000;
defparam \Decoder0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N5
dffeas \Reg[30][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][1] .is_wysiwyg = "true";
defparam \Reg[30][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N4
cycloneive_lcell_comb \Mux30~3 (
// Equation(s):
// \Mux30~3_combout  = (ifid_ifinstr_o_23 & ((\Mux30~2_combout  & (\Reg[30][1]~q )) # (!\Mux30~2_combout  & ((\Reg[22][1]~q ))))) # (!ifid_ifinstr_o_23 & (\Mux30~2_combout ))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux30~2_combout ),
	.datac(\Reg[30][1]~q ),
	.datad(\Reg[22][1]~q ),
	.cin(gnd),
	.combout(\Mux30~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~3 .lut_mask = 16'hE6C4;
defparam \Mux30~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N26
cycloneive_lcell_comb \Mux30~4 (
// Equation(s):
// \Mux30~4_combout  = (ifid_ifinstr_o_24 & ((\Reg[24][1]~q ) # ((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & (((\Reg[16][1]~q  & !ifid_ifinstr_o_23))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[24][1]~q ),
	.datac(\Reg[16][1]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux30~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~4 .lut_mask = 16'hAAD8;
defparam \Mux30~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N0
cycloneive_lcell_comb \Mux30~5 (
// Equation(s):
// \Mux30~5_combout  = (ifid_ifinstr_o_23 & ((\Mux30~4_combout  & (\Reg[28][1]~q )) # (!\Mux30~4_combout  & ((\Reg[20][1]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux30~4_combout ))))

	.dataa(\Reg[28][1]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[20][1]~q ),
	.datad(\Mux30~4_combout ),
	.cin(gnd),
	.combout(\Mux30~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~5 .lut_mask = 16'hBBC0;
defparam \Mux30~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N6
cycloneive_lcell_comb \Mux30~6 (
// Equation(s):
// \Mux30~6_combout  = (ifid_ifinstr_o_22 & ((\Mux30~3_combout ) # ((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & (((\Mux30~5_combout  & !ifid_ifinstr_o_21))))

	.dataa(\Mux30~3_combout ),
	.datab(\Mux30~5_combout ),
	.datac(ifid_ifinstr_o_22),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux30~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~6 .lut_mask = 16'hF0AC;
defparam \Mux30~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N0
cycloneive_lcell_comb \Mux30~7 (
// Equation(s):
// \Mux30~7_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & (\Reg[23][1]~q )) # (!ifid_ifinstr_o_23 & ((\Reg[19][1]~q )))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[23][1]~q ),
	.datad(\Reg[19][1]~q ),
	.cin(gnd),
	.combout(\Mux30~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~7 .lut_mask = 16'hD9C8;
defparam \Mux30~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N20
cycloneive_lcell_comb \Mux30~8 (
// Equation(s):
// \Mux30~8_combout  = (ifid_ifinstr_o_24 & ((\Mux30~7_combout  & ((\Reg[31][1]~q ))) # (!\Mux30~7_combout  & (\Reg[27][1]~q )))) # (!ifid_ifinstr_o_24 & (\Mux30~7_combout ))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux30~7_combout ),
	.datac(\Reg[27][1]~q ),
	.datad(\Reg[31][1]~q ),
	.cin(gnd),
	.combout(\Mux30~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~8 .lut_mask = 16'hEC64;
defparam \Mux30~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N16
cycloneive_lcell_comb \Mux30~10 (
// Equation(s):
// \Mux30~10_combout  = (ifid_ifinstr_o_21 & (ifid_ifinstr_o_22)) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[10][1]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[8][1]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[10][1]~q ),
	.datad(\Reg[8][1]~q ),
	.cin(gnd),
	.combout(\Mux30~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~10 .lut_mask = 16'hD9C8;
defparam \Mux30~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N20
cycloneive_lcell_comb \Mux30~11 (
// Equation(s):
// \Mux30~11_combout  = (ifid_ifinstr_o_21 & ((\Mux30~10_combout  & (\Reg[11][1]~q )) # (!\Mux30~10_combout  & ((\Reg[9][1]~q ))))) # (!ifid_ifinstr_o_21 & (((\Mux30~10_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[11][1]~q ),
	.datac(\Reg[9][1]~q ),
	.datad(\Mux30~10_combout ),
	.cin(gnd),
	.combout(\Mux30~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~11 .lut_mask = 16'hDDA0;
defparam \Mux30~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N24
cycloneive_lcell_comb \Decoder0~22 (
// Equation(s):
// \Decoder0~22_combout  = (!\rwWB~0_combout  & (!\rwWB~2_combout  & \Decoder0~18_combout ))

	.dataa(rwWB),
	.datab(gnd),
	.datac(rwWB2),
	.datad(\Decoder0~18_combout ),
	.cin(gnd),
	.combout(\Decoder0~22_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~22 .lut_mask = 16'h0500;
defparam \Decoder0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N31
dffeas \Reg[4][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][1] .is_wysiwyg = "true";
defparam \Reg[4][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N30
cycloneive_lcell_comb \Mux30~12 (
// Equation(s):
// \Mux30~12_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22) # ((\Reg[5][1]~q )))) # (!ifid_ifinstr_o_21 & (!ifid_ifinstr_o_22 & (\Reg[4][1]~q )))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[4][1]~q ),
	.datad(\Reg[5][1]~q ),
	.cin(gnd),
	.combout(\Mux30~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~12 .lut_mask = 16'hBA98;
defparam \Mux30~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N0
cycloneive_lcell_comb \Mux30~13 (
// Equation(s):
// \Mux30~13_combout  = (ifid_ifinstr_o_22 & ((\Mux30~12_combout  & (\Reg[7][1]~q )) # (!\Mux30~12_combout  & ((\Reg[6][1]~q ))))) # (!ifid_ifinstr_o_22 & (((\Mux30~12_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[7][1]~q ),
	.datac(\Mux30~12_combout ),
	.datad(\Reg[6][1]~q ),
	.cin(gnd),
	.combout(\Mux30~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~13 .lut_mask = 16'hDAD0;
defparam \Mux30~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N8
cycloneive_lcell_comb \Decoder0~31 (
// Equation(s):
// \Decoder0~31_combout  = (!\rwWB~2_combout  & (!\rwWB~0_combout  & \Decoder0~24_combout ))

	.dataa(rwWB2),
	.datab(rwWB),
	.datac(gnd),
	.datad(\Decoder0~24_combout ),
	.cin(gnd),
	.combout(\Decoder0~31_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~31 .lut_mask = 16'h1100;
defparam \Decoder0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N11
dffeas \Reg[1][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][1] .is_wysiwyg = "true";
defparam \Reg[1][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N14
cycloneive_lcell_comb \Decoder0~30 (
// Equation(s):
// \Decoder0~30_combout  = (!\rwWB~2_combout  & (\Decoder0~24_combout  & \rwWB~0_combout ))

	.dataa(rwWB2),
	.datab(\Decoder0~24_combout ),
	.datac(gnd),
	.datad(rwWB),
	.cin(gnd),
	.combout(\Decoder0~30_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~30 .lut_mask = 16'h4400;
defparam \Decoder0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N25
dffeas \Reg[3][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][1] .is_wysiwyg = "true";
defparam \Reg[3][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N10
cycloneive_lcell_comb \Mux30~14 (
// Equation(s):
// \Mux30~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][1]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][1]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[1][1]~q ),
	.datad(\Reg[3][1]~q ),
	.cin(gnd),
	.combout(\Mux30~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~14 .lut_mask = 16'hA820;
defparam \Mux30~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N6
cycloneive_lcell_comb \Mux30~15 (
// Equation(s):
// \Mux30~15_combout  = (\Mux30~14_combout ) # ((ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & \Reg[2][1]~q )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux30~14_combout ),
	.datad(\Reg[2][1]~q ),
	.cin(gnd),
	.combout(\Mux30~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~15 .lut_mask = 16'hF2F0;
defparam \Mux30~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N4
cycloneive_lcell_comb \Mux30~16 (
// Equation(s):
// \Mux30~16_combout  = (ifid_ifinstr_o_23 & ((\Mux30~13_combout ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((!ifid_ifinstr_o_24 & \Mux30~15_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux30~13_combout ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Mux30~15_combout ),
	.cin(gnd),
	.combout(\Mux30~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~16 .lut_mask = 16'hADA8;
defparam \Mux30~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N24
cycloneive_lcell_comb \Mux30~17 (
// Equation(s):
// \Mux30~17_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[13][1]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[12][1]~q ))))

	.dataa(\Reg[12][1]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[13][1]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux30~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~17 .lut_mask = 16'hFC22;
defparam \Mux30~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N6
cycloneive_lcell_comb \Mux30~18 (
// Equation(s):
// \Mux30~18_combout  = (ifid_ifinstr_o_22 & ((\Mux30~17_combout  & ((\Reg[15][1]~q ))) # (!\Mux30~17_combout  & (\Reg[14][1]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux30~17_combout ))))

	.dataa(\Reg[14][1]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[15][1]~q ),
	.datad(\Mux30~17_combout ),
	.cin(gnd),
	.combout(\Mux30~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~18 .lut_mask = 16'hF388;
defparam \Mux30~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N10
cycloneive_lcell_comb \Reg[25][0]~feeder (
// Equation(s):
// \Reg[25][0]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\Reg[25][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][0]~feeder .lut_mask = 16'hFF00;
defparam \Reg[25][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N11
dffeas \Reg[25][0] (
	.clk(!CLK),
	.d(\Reg[25][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][0] .is_wysiwyg = "true";
defparam \Reg[25][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N20
cycloneive_lcell_comb \Reg[29][0]~feeder (
// Equation(s):
// \Reg[29][0]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\Reg[29][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[29][0]~feeder .lut_mask = 16'hFF00;
defparam \Reg[29][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N21
dffeas \Reg[29][0] (
	.clk(!CLK),
	.d(\Reg[29][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][0] .is_wysiwyg = "true";
defparam \Reg[29][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N24
cycloneive_lcell_comb \Reg[21][0]~feeder (
// Equation(s):
// \Reg[21][0]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat1),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[21][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[21][0]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[21][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N25
dffeas \Reg[21][0] (
	.clk(!CLK),
	.d(\Reg[21][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][0] .is_wysiwyg = "true";
defparam \Reg[21][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N2
cycloneive_lcell_comb \Reg[17][0]~feeder (
// Equation(s):
// \Reg[17][0]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\Reg[17][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[17][0]~feeder .lut_mask = 16'hFF00;
defparam \Reg[17][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N3
dffeas \Reg[17][0] (
	.clk(!CLK),
	.d(\Reg[17][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][0] .is_wysiwyg = "true";
defparam \Reg[17][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N14
cycloneive_lcell_comb \Mux63~0 (
// Equation(s):
// \Mux63~0_combout  = (ifid_ifinstr_o_18 & ((\Reg[21][0]~q ) # ((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (((\Reg[17][0]~q  & !ifid_ifinstr_o_19))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[21][0]~q ),
	.datac(\Reg[17][0]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux63~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~0 .lut_mask = 16'hAAD8;
defparam \Mux63~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N26
cycloneive_lcell_comb \Mux63~1 (
// Equation(s):
// \Mux63~1_combout  = (\Mux63~0_combout  & (((\Reg[29][0]~q ) # (!ifid_ifinstr_o_19)))) # (!\Mux63~0_combout  & (\Reg[25][0]~q  & ((ifid_ifinstr_o_19))))

	.dataa(\Reg[25][0]~q ),
	.datab(\Reg[29][0]~q ),
	.datac(\Mux63~0_combout ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux63~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~1 .lut_mask = 16'hCAF0;
defparam \Mux63~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N27
dffeas \Reg[19][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][0] .is_wysiwyg = "true";
defparam \Reg[19][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N1
dffeas \Reg[23][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][0] .is_wysiwyg = "true";
defparam \Reg[23][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N26
cycloneive_lcell_comb \Mux63~7 (
// Equation(s):
// \Mux63~7_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Reg[23][0]~q ))) # (!ifid_ifinstr_o_18 & (\Reg[19][0]~q ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[19][0]~q ),
	.datad(\Reg[23][0]~q ),
	.cin(gnd),
	.combout(\Mux63~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~7 .lut_mask = 16'hDC98;
defparam \Mux63~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N1
dffeas \Reg[27][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][0] .is_wysiwyg = "true";
defparam \Reg[27][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N19
dffeas \Reg[31][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][0] .is_wysiwyg = "true";
defparam \Reg[31][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N18
cycloneive_lcell_comb \Mux63~8 (
// Equation(s):
// \Mux63~8_combout  = (\Mux63~7_combout  & (((\Reg[31][0]~q ) # (!ifid_ifinstr_o_19)))) # (!\Mux63~7_combout  & (\Reg[27][0]~q  & ((ifid_ifinstr_o_19))))

	.dataa(\Mux63~7_combout ),
	.datab(\Reg[27][0]~q ),
	.datac(\Reg[31][0]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux63~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~8 .lut_mask = 16'hE4AA;
defparam \Mux63~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N10
cycloneive_lcell_comb \Reg[28][0]~feeder (
// Equation(s):
// \Reg[28][0]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\Reg[28][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[28][0]~feeder .lut_mask = 16'hFF00;
defparam \Reg[28][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N11
dffeas \Reg[28][0] (
	.clk(!CLK),
	.d(\Reg[28][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][0] .is_wysiwyg = "true";
defparam \Reg[28][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y34_N17
dffeas \Reg[24][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][0] .is_wysiwyg = "true";
defparam \Reg[24][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N18
cycloneive_lcell_comb \Reg[16][0]~feeder (
// Equation(s):
// \Reg[16][0]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat1),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[16][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[16][0]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[16][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y34_N19
dffeas \Reg[16][0] (
	.clk(!CLK),
	.d(\Reg[16][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][0] .is_wysiwyg = "true";
defparam \Reg[16][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N16
cycloneive_lcell_comb \Mux63~4 (
// Equation(s):
// \Mux63~4_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Reg[24][0]~q )) # (!ifid_ifinstr_o_19 & ((\Reg[16][0]~q )))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[24][0]~q ),
	.datad(\Reg[16][0]~q ),
	.cin(gnd),
	.combout(\Mux63~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~4 .lut_mask = 16'hD9C8;
defparam \Mux63~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N0
cycloneive_lcell_comb \Mux63~5 (
// Equation(s):
// \Mux63~5_combout  = (\Mux63~4_combout  & (((\Reg[28][0]~q ) # (!ifid_ifinstr_o_18)))) # (!\Mux63~4_combout  & (\Reg[20][0]~q  & ((ifid_ifinstr_o_18))))

	.dataa(\Reg[20][0]~q ),
	.datab(\Reg[28][0]~q ),
	.datac(\Mux63~4_combout ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux63~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~5 .lut_mask = 16'hCAF0;
defparam \Mux63~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N26
cycloneive_lcell_comb \Reg[30][0]~feeder (
// Equation(s):
// \Reg[30][0]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat1),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[30][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[30][0]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[30][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N27
dffeas \Reg[30][0] (
	.clk(!CLK),
	.d(\Reg[30][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][0] .is_wysiwyg = "true";
defparam \Reg[30][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N15
dffeas \Reg[18][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][0] .is_wysiwyg = "true";
defparam \Reg[18][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N13
dffeas \Reg[26][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][0] .is_wysiwyg = "true";
defparam \Reg[26][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N8
cycloneive_lcell_comb \Mux63~2 (
// Equation(s):
// \Mux63~2_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[26][0]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[18][0]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[18][0]~q ),
	.datad(\Reg[26][0]~q ),
	.cin(gnd),
	.combout(\Mux63~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~2 .lut_mask = 16'hDC98;
defparam \Mux63~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N16
cycloneive_lcell_comb \Reg[22][0]~feeder (
// Equation(s):
// \Reg[22][0]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\Reg[22][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[22][0]~feeder .lut_mask = 16'hFF00;
defparam \Reg[22][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N17
dffeas \Reg[22][0] (
	.clk(!CLK),
	.d(\Reg[22][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][0] .is_wysiwyg = "true";
defparam \Reg[22][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N26
cycloneive_lcell_comb \Mux63~3 (
// Equation(s):
// \Mux63~3_combout  = (ifid_ifinstr_o_18 & ((\Mux63~2_combout  & (\Reg[30][0]~q )) # (!\Mux63~2_combout  & ((\Reg[22][0]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux63~2_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[30][0]~q ),
	.datac(\Mux63~2_combout ),
	.datad(\Reg[22][0]~q ),
	.cin(gnd),
	.combout(\Mux63~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~3 .lut_mask = 16'hDAD0;
defparam \Mux63~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N28
cycloneive_lcell_comb \Mux63~6 (
// Equation(s):
// \Mux63~6_combout  = (ifid_ifinstr_o_16 & (((ifid_ifinstr_o_17)))) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Mux63~3_combout ))) # (!ifid_ifinstr_o_17 & (\Mux63~5_combout ))))

	.dataa(\Mux63~5_combout ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux63~3_combout ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux63~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~6 .lut_mask = 16'hFC22;
defparam \Mux63~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N10
cycloneive_lcell_comb \Reg[15][0]~feeder (
// Equation(s):
// \Reg[15][0]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat1),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[15][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[15][0]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[15][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N11
dffeas \Reg[15][0] (
	.clk(!CLK),
	.d(\Reg[15][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][0] .is_wysiwyg = "true";
defparam \Reg[15][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N20
cycloneive_lcell_comb \Reg[14][0]~feeder (
// Equation(s):
// \Reg[14][0]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat1),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[14][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[14][0]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[14][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N21
dffeas \Reg[14][0] (
	.clk(!CLK),
	.d(\Reg[14][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][0] .is_wysiwyg = "true";
defparam \Reg[14][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N13
dffeas \Reg[13][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][0] .is_wysiwyg = "true";
defparam \Reg[13][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N12
cycloneive_lcell_comb \Mux63~17 (
// Equation(s):
// \Mux63~17_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[13][0]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[12][0]~q ))))

	.dataa(\Reg[12][0]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[13][0]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux63~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~17 .lut_mask = 16'hFC22;
defparam \Mux63~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N28
cycloneive_lcell_comb \Mux63~18 (
// Equation(s):
// \Mux63~18_combout  = (ifid_ifinstr_o_17 & ((\Mux63~17_combout  & (\Reg[15][0]~q )) # (!\Mux63~17_combout  & ((\Reg[14][0]~q ))))) # (!ifid_ifinstr_o_17 & (((\Mux63~17_combout ))))

	.dataa(\Reg[15][0]~q ),
	.datab(\Reg[14][0]~q ),
	.datac(ifid_ifinstr_o_17),
	.datad(\Mux63~17_combout ),
	.cin(gnd),
	.combout(\Mux63~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~18 .lut_mask = 16'hAFC0;
defparam \Mux63~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N15
dffeas \Reg[1][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][0] .is_wysiwyg = "true";
defparam \Reg[1][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N16
cycloneive_lcell_comb \Reg[3][0]~feeder (
// Equation(s):
// \Reg[3][0]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat1),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[3][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[3][0]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[3][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N17
dffeas \Reg[3][0] (
	.clk(!CLK),
	.d(\Reg[3][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][0] .is_wysiwyg = "true";
defparam \Reg[3][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N4
cycloneive_lcell_comb \Mux63~14 (
// Equation(s):
// \Mux63~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[3][0]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[1][0]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[1][0]~q ),
	.datad(\Reg[3][0]~q ),
	.cin(gnd),
	.combout(\Mux63~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~14 .lut_mask = 16'hA820;
defparam \Mux63~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N14
cycloneive_lcell_comb \Reg[2][0]~feeder (
// Equation(s):
// \Reg[2][0]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\Reg[2][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[2][0]~feeder .lut_mask = 16'hFF00;
defparam \Reg[2][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N15
dffeas \Reg[2][0] (
	.clk(!CLK),
	.d(\Reg[2][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][0] .is_wysiwyg = "true";
defparam \Reg[2][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N22
cycloneive_lcell_comb \Mux63~15 (
// Equation(s):
// \Mux63~15_combout  = (\Mux63~14_combout ) # ((!ifid_ifinstr_o_16 & (ifid_ifinstr_o_17 & \Reg[2][0]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux63~14_combout ),
	.datad(\Reg[2][0]~q ),
	.cin(gnd),
	.combout(\Mux63~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~15 .lut_mask = 16'hF4F0;
defparam \Mux63~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N23
dffeas \Reg[4][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][0] .is_wysiwyg = "true";
defparam \Reg[4][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N25
dffeas \Reg[5][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][0] .is_wysiwyg = "true";
defparam \Reg[5][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N22
cycloneive_lcell_comb \Mux63~12 (
// Equation(s):
// \Mux63~12_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17) # ((\Reg[5][0]~q )))) # (!ifid_ifinstr_o_16 & (!ifid_ifinstr_o_17 & (\Reg[4][0]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[4][0]~q ),
	.datad(\Reg[5][0]~q ),
	.cin(gnd),
	.combout(\Mux63~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~12 .lut_mask = 16'hBA98;
defparam \Mux63~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N3
dffeas \Reg[7][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][0] .is_wysiwyg = "true";
defparam \Reg[7][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y39_N1
dffeas \Reg[6][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][0] .is_wysiwyg = "true";
defparam \Reg[6][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N2
cycloneive_lcell_comb \Mux63~13 (
// Equation(s):
// \Mux63~13_combout  = (ifid_ifinstr_o_17 & ((\Mux63~12_combout  & (\Reg[7][0]~q )) # (!\Mux63~12_combout  & ((\Reg[6][0]~q ))))) # (!ifid_ifinstr_o_17 & (\Mux63~12_combout ))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux63~12_combout ),
	.datac(\Reg[7][0]~q ),
	.datad(\Reg[6][0]~q ),
	.cin(gnd),
	.combout(\Mux63~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~13 .lut_mask = 16'hE6C4;
defparam \Mux63~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N0
cycloneive_lcell_comb \Mux63~16 (
// Equation(s):
// \Mux63~16_combout  = (ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19) # ((\Mux63~13_combout )))) # (!ifid_ifinstr_o_18 & (!ifid_ifinstr_o_19 & (\Mux63~15_combout )))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Mux63~15_combout ),
	.datad(\Mux63~13_combout ),
	.cin(gnd),
	.combout(\Mux63~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~16 .lut_mask = 16'hBA98;
defparam \Mux63~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N23
dffeas \Reg[11][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][0] .is_wysiwyg = "true";
defparam \Reg[11][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N1
dffeas \Reg[10][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][0] .is_wysiwyg = "true";
defparam \Reg[10][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N19
dffeas \Reg[8][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][0] .is_wysiwyg = "true";
defparam \Reg[8][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N0
cycloneive_lcell_comb \Mux63~10 (
// Equation(s):
// \Mux63~10_combout  = (ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16) # ((\Reg[10][0]~q )))) # (!ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & ((\Reg[8][0]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[10][0]~q ),
	.datad(\Reg[8][0]~q ),
	.cin(gnd),
	.combout(\Mux63~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~10 .lut_mask = 16'hB9A8;
defparam \Mux63~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N5
dffeas \Reg[9][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][0] .is_wysiwyg = "true";
defparam \Reg[9][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N4
cycloneive_lcell_comb \Mux63~11 (
// Equation(s):
// \Mux63~11_combout  = (\Mux63~10_combout  & ((\Reg[11][0]~q ) # ((!ifid_ifinstr_o_16)))) # (!\Mux63~10_combout  & (((\Reg[9][0]~q  & ifid_ifinstr_o_16))))

	.dataa(\Reg[11][0]~q ),
	.datab(\Mux63~10_combout ),
	.datac(\Reg[9][0]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux63~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~11 .lut_mask = 16'hB8CC;
defparam \Mux63~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N12
cycloneive_lcell_comb \Mux31~0 (
// Equation(s):
// \Mux31~0_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[25][0]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[17][0]~q )))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[25][0]~q ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Reg[17][0]~q ),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~0 .lut_mask = 16'hE5E0;
defparam \Mux31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N16
cycloneive_lcell_comb \Mux31~1 (
// Equation(s):
// \Mux31~1_combout  = (\Mux31~0_combout  & (((\Reg[29][0]~q ) # (!ifid_ifinstr_o_23)))) # (!\Mux31~0_combout  & (\Reg[21][0]~q  & (ifid_ifinstr_o_23)))

	.dataa(\Mux31~0_combout ),
	.datab(\Reg[21][0]~q ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Reg[29][0]~q ),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~1 .lut_mask = 16'hEA4A;
defparam \Mux31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N0
cycloneive_lcell_comb \Mux31~7 (
// Equation(s):
// \Mux31~7_combout  = (ifid_ifinstr_o_24 & (((\Reg[27][0]~q ) # (ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & (\Reg[19][0]~q  & ((!ifid_ifinstr_o_23))))

	.dataa(\Reg[19][0]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[27][0]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux31~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~7 .lut_mask = 16'hCCE2;
defparam \Mux31~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N0
cycloneive_lcell_comb \Mux31~8 (
// Equation(s):
// \Mux31~8_combout  = (ifid_ifinstr_o_23 & ((\Mux31~7_combout  & ((\Reg[31][0]~q ))) # (!\Mux31~7_combout  & (\Reg[23][0]~q )))) # (!ifid_ifinstr_o_23 & (\Mux31~7_combout ))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux31~7_combout ),
	.datac(\Reg[23][0]~q ),
	.datad(\Reg[31][0]~q ),
	.cin(gnd),
	.combout(\Mux31~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~8 .lut_mask = 16'hEC64;
defparam \Mux31~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N12
cycloneive_lcell_comb \Reg[20][0]~feeder (
// Equation(s):
// \Reg[20][0]~feeder_combout  = \wdat~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat1),
	.cin(gnd),
	.combout(\Reg[20][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[20][0]~feeder .lut_mask = 16'hFF00;
defparam \Reg[20][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N13
dffeas \Reg[20][0] (
	.clk(!CLK),
	.d(\Reg[20][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][0] .is_wysiwyg = "true";
defparam \Reg[20][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N8
cycloneive_lcell_comb \Mux31~4 (
// Equation(s):
// \Mux31~4_combout  = (ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24) # ((\Reg[20][0]~q )))) # (!ifid_ifinstr_o_23 & (!ifid_ifinstr_o_24 & ((\Reg[16][0]~q ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[20][0]~q ),
	.datad(\Reg[16][0]~q ),
	.cin(gnd),
	.combout(\Mux31~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~4 .lut_mask = 16'hB9A8;
defparam \Mux31~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N22
cycloneive_lcell_comb \Mux31~5 (
// Equation(s):
// \Mux31~5_combout  = (ifid_ifinstr_o_24 & ((\Mux31~4_combout  & (\Reg[28][0]~q )) # (!\Mux31~4_combout  & ((\Reg[24][0]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux31~4_combout ))))

	.dataa(\Reg[28][0]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Mux31~4_combout ),
	.datad(\Reg[24][0]~q ),
	.cin(gnd),
	.combout(\Mux31~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~5 .lut_mask = 16'hBCB0;
defparam \Mux31~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N14
cycloneive_lcell_comb \Mux31~2 (
// Equation(s):
// \Mux31~2_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[22][0]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[18][0]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[18][0]~q ),
	.datad(\Reg[22][0]~q ),
	.cin(gnd),
	.combout(\Mux31~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~2 .lut_mask = 16'hDC98;
defparam \Mux31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N20
cycloneive_lcell_comb \Mux31~3 (
// Equation(s):
// \Mux31~3_combout  = (\Mux31~2_combout  & (((\Reg[30][0]~q ) # (!ifid_ifinstr_o_24)))) # (!\Mux31~2_combout  & (\Reg[26][0]~q  & ((ifid_ifinstr_o_24))))

	.dataa(\Reg[26][0]~q ),
	.datab(\Mux31~2_combout ),
	.datac(\Reg[30][0]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux31~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~3 .lut_mask = 16'hE2CC;
defparam \Mux31~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N16
cycloneive_lcell_comb \Mux31~6 (
// Equation(s):
// \Mux31~6_combout  = (ifid_ifinstr_o_21 & (ifid_ifinstr_o_22)) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Mux31~3_combout ))) # (!ifid_ifinstr_o_22 & (\Mux31~5_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Mux31~5_combout ),
	.datad(\Mux31~3_combout ),
	.cin(gnd),
	.combout(\Mux31~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~6 .lut_mask = 16'hDC98;
defparam \Mux31~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N31
dffeas \Reg[12][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat1),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][0] .is_wysiwyg = "true";
defparam \Reg[12][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N30
cycloneive_lcell_comb \Mux31~17 (
// Equation(s):
// \Mux31~17_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22) # ((\Reg[13][0]~q )))) # (!ifid_ifinstr_o_21 & (!ifid_ifinstr_o_22 & (\Reg[12][0]~q )))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[12][0]~q ),
	.datad(\Reg[13][0]~q ),
	.cin(gnd),
	.combout(\Mux31~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~17 .lut_mask = 16'hBA98;
defparam \Mux31~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N20
cycloneive_lcell_comb \Mux31~18 (
// Equation(s):
// \Mux31~18_combout  = (\Mux31~17_combout  & (((\Reg[15][0]~q ) # (!ifid_ifinstr_o_22)))) # (!\Mux31~17_combout  & (\Reg[14][0]~q  & ((ifid_ifinstr_o_22))))

	.dataa(\Reg[14][0]~q ),
	.datab(\Reg[15][0]~q ),
	.datac(\Mux31~17_combout ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux31~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~18 .lut_mask = 16'hCAF0;
defparam \Mux31~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N14
cycloneive_lcell_comb \Mux31~14 (
// Equation(s):
// \Mux31~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][0]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][0]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[1][0]~q ),
	.datad(\Reg[3][0]~q ),
	.cin(gnd),
	.combout(\Mux31~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~14 .lut_mask = 16'hA820;
defparam \Mux31~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N8
cycloneive_lcell_comb \Mux31~15 (
// Equation(s):
// \Mux31~15_combout  = (\Mux31~14_combout ) # ((\Reg[2][0]~q  & (!ifid_ifinstr_o_21 & ifid_ifinstr_o_22)))

	.dataa(\Reg[2][0]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux31~14_combout ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux31~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~15 .lut_mask = 16'hF2F0;
defparam \Mux31~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N18
cycloneive_lcell_comb \Mux31~12 (
// Equation(s):
// \Mux31~12_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[10][0]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[8][0]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[10][0]~q ),
	.datac(\Reg[8][0]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux31~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~12 .lut_mask = 16'hEE50;
defparam \Mux31~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N22
cycloneive_lcell_comb \Mux31~13 (
// Equation(s):
// \Mux31~13_combout  = (ifid_ifinstr_o_21 & ((\Mux31~12_combout  & ((\Reg[11][0]~q ))) # (!\Mux31~12_combout  & (\Reg[9][0]~q )))) # (!ifid_ifinstr_o_21 & (((\Mux31~12_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[9][0]~q ),
	.datac(\Reg[11][0]~q ),
	.datad(\Mux31~12_combout ),
	.cin(gnd),
	.combout(\Mux31~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~13 .lut_mask = 16'hF588;
defparam \Mux31~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N22
cycloneive_lcell_comb \Mux31~16 (
// Equation(s):
// \Mux31~16_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Mux31~13_combout ))) # (!ifid_ifinstr_o_24 & (\Mux31~15_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux31~15_combout ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Mux31~13_combout ),
	.cin(gnd),
	.combout(\Mux31~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~16 .lut_mask = 16'hF4A4;
defparam \Mux31~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N24
cycloneive_lcell_comb \Mux31~10 (
// Equation(s):
// \Mux31~10_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[5][0]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[4][0]~q ))))

	.dataa(\Reg[4][0]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[5][0]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux31~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~10 .lut_mask = 16'hFC22;
defparam \Mux31~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N0
cycloneive_lcell_comb \Mux31~11 (
// Equation(s):
// \Mux31~11_combout  = (\Mux31~10_combout  & (((\Reg[7][0]~q )) # (!ifid_ifinstr_o_22))) # (!\Mux31~10_combout  & (ifid_ifinstr_o_22 & (\Reg[6][0]~q )))

	.dataa(\Mux31~10_combout ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[6][0]~q ),
	.datad(\Reg[7][0]~q ),
	.cin(gnd),
	.combout(\Mux31~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~11 .lut_mask = 16'hEA62;
defparam \Mux31~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N24
cycloneive_lcell_comb \Reg[21][2]~feeder (
// Equation(s):
// \Reg[21][2]~feeder_combout  = \wdat~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat2),
	.cin(gnd),
	.combout(\Reg[21][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[21][2]~feeder .lut_mask = 16'hFF00;
defparam \Reg[21][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N25
dffeas \Reg[21][2] (
	.clk(!CLK),
	.d(\Reg[21][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][2] .is_wysiwyg = "true";
defparam \Reg[21][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N2
cycloneive_lcell_comb \Reg[29][2]~feeder (
// Equation(s):
// \Reg[29][2]~feeder_combout  = \wdat~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat2),
	.cin(gnd),
	.combout(\Reg[29][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[29][2]~feeder .lut_mask = 16'hFF00;
defparam \Reg[29][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N3
dffeas \Reg[29][2] (
	.clk(!CLK),
	.d(\Reg[29][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][2] .is_wysiwyg = "true";
defparam \Reg[29][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N0
cycloneive_lcell_comb \Reg[17][2]~feeder (
// Equation(s):
// \Reg[17][2]~feeder_combout  = \wdat~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat2),
	.cin(gnd),
	.combout(\Reg[17][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[17][2]~feeder .lut_mask = 16'hFF00;
defparam \Reg[17][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N1
dffeas \Reg[17][2] (
	.clk(!CLK),
	.d(\Reg[17][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][2] .is_wysiwyg = "true";
defparam \Reg[17][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N22
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[25][2]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[17][2]~q )))))

	.dataa(\Reg[25][2]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(ifid_ifinstr_o_24),
	.datad(\Reg[17][2]~q ),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'hE3E0;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N0
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// \Mux29~1_combout  = (ifid_ifinstr_o_23 & ((\Mux29~0_combout  & ((\Reg[29][2]~q ))) # (!\Mux29~0_combout  & (\Reg[21][2]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux29~0_combout ))))

	.dataa(\Reg[21][2]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[29][2]~q ),
	.datad(\Mux29~0_combout ),
	.cin(gnd),
	.combout(\Mux29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'hF388;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N5
dffeas \Reg[27][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][2] .is_wysiwyg = "true";
defparam \Reg[27][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N23
dffeas \Reg[19][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][2] .is_wysiwyg = "true";
defparam \Reg[19][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N4
cycloneive_lcell_comb \Mux29~7 (
// Equation(s):
// \Mux29~7_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[27][2]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[19][2]~q )))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[27][2]~q ),
	.datad(\Reg[19][2]~q ),
	.cin(gnd),
	.combout(\Mux29~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~7 .lut_mask = 16'hD9C8;
defparam \Mux29~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N7
dffeas \Reg[31][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][2] .is_wysiwyg = "true";
defparam \Reg[31][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N24
cycloneive_lcell_comb \Reg[23][2]~feeder (
// Equation(s):
// \Reg[23][2]~feeder_combout  = \wdat~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat2),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[23][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[23][2]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[23][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N25
dffeas \Reg[23][2] (
	.clk(!CLK),
	.d(\Reg[23][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][2] .is_wysiwyg = "true";
defparam \Reg[23][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N6
cycloneive_lcell_comb \Mux29~8 (
// Equation(s):
// \Mux29~8_combout  = (ifid_ifinstr_o_23 & ((\Mux29~7_combout  & (\Reg[31][2]~q )) # (!\Mux29~7_combout  & ((\Reg[23][2]~q ))))) # (!ifid_ifinstr_o_23 & (\Mux29~7_combout ))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux29~7_combout ),
	.datac(\Reg[31][2]~q ),
	.datad(\Reg[23][2]~q ),
	.cin(gnd),
	.combout(\Mux29~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~8 .lut_mask = 16'hE6C4;
defparam \Mux29~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y30_N25
dffeas \Reg[26][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][2] .is_wysiwyg = "true";
defparam \Reg[26][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N27
dffeas \Reg[18][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][2] .is_wysiwyg = "true";
defparam \Reg[18][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y30_N13
dffeas \Reg[22][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][2] .is_wysiwyg = "true";
defparam \Reg[22][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N12
cycloneive_lcell_comb \Mux29~2 (
// Equation(s):
// \Mux29~2_combout  = (ifid_ifinstr_o_23 & (((\Reg[22][2]~q ) # (ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (\Reg[18][2]~q  & ((!ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[18][2]~q ),
	.datac(\Reg[22][2]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux29~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~2 .lut_mask = 16'hAAE4;
defparam \Mux29~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N24
cycloneive_lcell_comb \Mux29~3 (
// Equation(s):
// \Mux29~3_combout  = (ifid_ifinstr_o_24 & ((\Mux29~2_combout  & (\Reg[30][2]~q )) # (!\Mux29~2_combout  & ((\Reg[26][2]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux29~2_combout ))))

	.dataa(\Reg[30][2]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[26][2]~q ),
	.datad(\Mux29~2_combout ),
	.cin(gnd),
	.combout(\Mux29~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~3 .lut_mask = 16'hBBC0;
defparam \Mux29~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y34_N13
dffeas \Reg[24][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][2] .is_wysiwyg = "true";
defparam \Reg[24][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y34_N23
dffeas \Reg[28][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][2] .is_wysiwyg = "true";
defparam \Reg[28][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y34_N15
dffeas \Reg[16][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][2] .is_wysiwyg = "true";
defparam \Reg[16][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y34_N1
dffeas \Reg[20][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][2] .is_wysiwyg = "true";
defparam \Reg[20][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N14
cycloneive_lcell_comb \Mux29~4 (
// Equation(s):
// \Mux29~4_combout  = (ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24) # ((\Reg[20][2]~q )))) # (!ifid_ifinstr_o_23 & (!ifid_ifinstr_o_24 & (\Reg[16][2]~q )))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[16][2]~q ),
	.datad(\Reg[20][2]~q ),
	.cin(gnd),
	.combout(\Mux29~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~4 .lut_mask = 16'hBA98;
defparam \Mux29~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N22
cycloneive_lcell_comb \Mux29~5 (
// Equation(s):
// \Mux29~5_combout  = (ifid_ifinstr_o_24 & ((\Mux29~4_combout  & ((\Reg[28][2]~q ))) # (!\Mux29~4_combout  & (\Reg[24][2]~q )))) # (!ifid_ifinstr_o_24 & (((\Mux29~4_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[24][2]~q ),
	.datac(\Reg[28][2]~q ),
	.datad(\Mux29~4_combout ),
	.cin(gnd),
	.combout(\Mux29~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~5 .lut_mask = 16'hF588;
defparam \Mux29~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N30
cycloneive_lcell_comb \Mux29~6 (
// Equation(s):
// \Mux29~6_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Mux29~3_combout )) # (!ifid_ifinstr_o_22 & ((\Mux29~5_combout )))))

	.dataa(\Mux29~3_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(ifid_ifinstr_o_22),
	.datad(\Mux29~5_combout ),
	.cin(gnd),
	.combout(\Mux29~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~6 .lut_mask = 16'hE3E0;
defparam \Mux29~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N15
dffeas \Reg[4][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][2] .is_wysiwyg = "true";
defparam \Reg[4][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N29
dffeas \Reg[5][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][2] .is_wysiwyg = "true";
defparam \Reg[5][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N28
cycloneive_lcell_comb \Mux29~10 (
// Equation(s):
// \Mux29~10_combout  = (ifid_ifinstr_o_21 & (((\Reg[5][2]~q ) # (ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & (\Reg[4][2]~q  & ((!ifid_ifinstr_o_22))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[4][2]~q ),
	.datac(\Reg[5][2]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux29~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~10 .lut_mask = 16'hAAE4;
defparam \Mux29~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N16
cycloneive_lcell_comb \Reg[6][2]~feeder (
// Equation(s):
// \Reg[6][2]~feeder_combout  = \wdat~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat2),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[6][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[6][2]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[6][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N17
dffeas \Reg[6][2] (
	.clk(!CLK),
	.d(\Reg[6][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][2] .is_wysiwyg = "true";
defparam \Reg[6][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y39_N23
dffeas \Reg[7][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][2] .is_wysiwyg = "true";
defparam \Reg[7][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N24
cycloneive_lcell_comb \Mux29~11 (
// Equation(s):
// \Mux29~11_combout  = (\Mux29~10_combout  & (((\Reg[7][2]~q ) # (!ifid_ifinstr_o_22)))) # (!\Mux29~10_combout  & (\Reg[6][2]~q  & ((ifid_ifinstr_o_22))))

	.dataa(\Mux29~10_combout ),
	.datab(\Reg[6][2]~q ),
	.datac(\Reg[7][2]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux29~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~11 .lut_mask = 16'hE4AA;
defparam \Mux29~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y34_N21
dffeas \Reg[12][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][2] .is_wysiwyg = "true";
defparam \Reg[12][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N3
dffeas \Reg[13][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][2] .is_wysiwyg = "true";
defparam \Reg[13][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N20
cycloneive_lcell_comb \Mux29~17 (
// Equation(s):
// \Mux29~17_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[13][2]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[12][2]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[12][2]~q ),
	.datad(\Reg[13][2]~q ),
	.cin(gnd),
	.combout(\Mux29~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~17 .lut_mask = 16'hDC98;
defparam \Mux29~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y37_N3
dffeas \Reg[15][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][2] .is_wysiwyg = "true";
defparam \Reg[15][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y37_N13
dffeas \Reg[14][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][2] .is_wysiwyg = "true";
defparam \Reg[14][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N2
cycloneive_lcell_comb \Mux29~18 (
// Equation(s):
// \Mux29~18_combout  = (ifid_ifinstr_o_22 & ((\Mux29~17_combout  & (\Reg[15][2]~q )) # (!\Mux29~17_combout  & ((\Reg[14][2]~q ))))) # (!ifid_ifinstr_o_22 & (\Mux29~17_combout ))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Mux29~17_combout ),
	.datac(\Reg[15][2]~q ),
	.datad(\Reg[14][2]~q ),
	.cin(gnd),
	.combout(\Mux29~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~18 .lut_mask = 16'hE6C4;
defparam \Mux29~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N13
dffeas \Reg[2][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][2] .is_wysiwyg = "true";
defparam \Reg[2][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N1
dffeas \Reg[3][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][2] .is_wysiwyg = "true";
defparam \Reg[3][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N0
cycloneive_lcell_comb \Mux29~14 (
// Equation(s):
// \Mux29~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][2]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][2]~q ))))

	.dataa(\Reg[1][2]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[3][2]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux29~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~14 .lut_mask = 16'hC088;
defparam \Mux29~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N12
cycloneive_lcell_comb \Mux29~15 (
// Equation(s):
// \Mux29~15_combout  = (\Mux29~14_combout ) # ((ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & \Reg[2][2]~q )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[2][2]~q ),
	.datad(\Mux29~14_combout ),
	.cin(gnd),
	.combout(\Mux29~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~15 .lut_mask = 16'hFF20;
defparam \Mux29~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N25
dffeas \Reg[9][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][2] .is_wysiwyg = "true";
defparam \Reg[9][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N7
dffeas \Reg[11][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][2] .is_wysiwyg = "true";
defparam \Reg[11][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N25
dffeas \Reg[10][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][2] .is_wysiwyg = "true";
defparam \Reg[10][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N31
dffeas \Reg[8][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][2] .is_wysiwyg = "true";
defparam \Reg[8][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N30
cycloneive_lcell_comb \Mux29~12 (
// Equation(s):
// \Mux29~12_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[10][2]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[8][2]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[10][2]~q ),
	.datac(\Reg[8][2]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux29~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~12 .lut_mask = 16'hEE50;
defparam \Mux29~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N6
cycloneive_lcell_comb \Mux29~13 (
// Equation(s):
// \Mux29~13_combout  = (ifid_ifinstr_o_21 & ((\Mux29~12_combout  & ((\Reg[11][2]~q ))) # (!\Mux29~12_combout  & (\Reg[9][2]~q )))) # (!ifid_ifinstr_o_21 & (((\Mux29~12_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[9][2]~q ),
	.datac(\Reg[11][2]~q ),
	.datad(\Mux29~12_combout ),
	.cin(gnd),
	.combout(\Mux29~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~13 .lut_mask = 16'hF588;
defparam \Mux29~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N12
cycloneive_lcell_comb \Mux29~16 (
// Equation(s):
// \Mux29~16_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23) # (\Mux29~13_combout )))) # (!ifid_ifinstr_o_24 & (\Mux29~15_combout  & (!ifid_ifinstr_o_23)))

	.dataa(\Mux29~15_combout ),
	.datab(ifid_ifinstr_o_24),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux29~13_combout ),
	.cin(gnd),
	.combout(\Mux29~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~16 .lut_mask = 16'hCEC2;
defparam \Mux29~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N22
cycloneive_lcell_comb \Reg[29][4]~feeder (
// Equation(s):
// \Reg[29][4]~feeder_combout  = \wdat~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat3),
	.cin(gnd),
	.combout(\Reg[29][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[29][4]~feeder .lut_mask = 16'hFF00;
defparam \Reg[29][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N23
dffeas \Reg[29][4] (
	.clk(!CLK),
	.d(\Reg[29][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][4] .is_wysiwyg = "true";
defparam \Reg[29][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N21
dffeas \Reg[17][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][4] .is_wysiwyg = "true";
defparam \Reg[17][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N14
cycloneive_lcell_comb \Reg[25][4]~feeder (
// Equation(s):
// \Reg[25][4]~feeder_combout  = \wdat~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat3),
	.cin(gnd),
	.combout(\Reg[25][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][4]~feeder .lut_mask = 16'hFF00;
defparam \Reg[25][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N15
dffeas \Reg[25][4] (
	.clk(!CLK),
	.d(\Reg[25][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][4] .is_wysiwyg = "true";
defparam \Reg[25][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N20
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Reg[25][4]~q ))) # (!ifid_ifinstr_o_24 & (\Reg[17][4]~q ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[17][4]~q ),
	.datad(\Reg[25][4]~q ),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'hDC98;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N13
dffeas \Reg[21][4] (
	.clk(!CLK),
	.d(wdat3),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][4] .is_wysiwyg = "true";
defparam \Reg[21][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N0
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// \Mux27~1_combout  = (\Mux27~0_combout  & ((\Reg[29][4]~q ) # ((!ifid_ifinstr_o_23)))) # (!\Mux27~0_combout  & (((ifid_ifinstr_o_23 & \Reg[21][4]~q ))))

	.dataa(\Reg[29][4]~q ),
	.datab(\Mux27~0_combout ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Reg[21][4]~q ),
	.cin(gnd),
	.combout(\Mux27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hBC8C;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y34_N31
dffeas \Reg[16][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][4] .is_wysiwyg = "true";
defparam \Reg[16][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N4
cycloneive_lcell_comb \Reg[20][4]~feeder (
// Equation(s):
// \Reg[20][4]~feeder_combout  = \wdat~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat3),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[20][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[20][4]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[20][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N5
dffeas \Reg[20][4] (
	.clk(!CLK),
	.d(\Reg[20][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][4] .is_wysiwyg = "true";
defparam \Reg[20][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N30
cycloneive_lcell_comb \Mux27~4 (
// Equation(s):
// \Mux27~4_combout  = (ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24) # ((\Reg[20][4]~q )))) # (!ifid_ifinstr_o_23 & (!ifid_ifinstr_o_24 & (\Reg[16][4]~q )))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[16][4]~q ),
	.datad(\Reg[20][4]~q ),
	.cin(gnd),
	.combout(\Mux27~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~4 .lut_mask = 16'hBA98;
defparam \Mux27~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y34_N25
dffeas \Reg[24][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][4] .is_wysiwyg = "true";
defparam \Reg[24][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N7
dffeas \Reg[28][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][4] .is_wysiwyg = "true";
defparam \Reg[28][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N24
cycloneive_lcell_comb \Mux27~5 (
// Equation(s):
// \Mux27~5_combout  = (ifid_ifinstr_o_24 & ((\Mux27~4_combout  & ((\Reg[28][4]~q ))) # (!\Mux27~4_combout  & (\Reg[24][4]~q )))) # (!ifid_ifinstr_o_24 & (\Mux27~4_combout ))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux27~4_combout ),
	.datac(\Reg[24][4]~q ),
	.datad(\Reg[28][4]~q ),
	.cin(gnd),
	.combout(\Mux27~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~5 .lut_mask = 16'hEC64;
defparam \Mux27~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N16
cycloneive_lcell_comb \Reg[22][4]~feeder (
// Equation(s):
// \Reg[22][4]~feeder_combout  = \wdat~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat3),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[22][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[22][4]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[22][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N17
dffeas \Reg[22][4] (
	.clk(!CLK),
	.d(\Reg[22][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][4] .is_wysiwyg = "true";
defparam \Reg[22][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N24
cycloneive_lcell_comb \Mux27~2 (
// Equation(s):
// \Mux27~2_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24) # (\Reg[22][4]~q )))) # (!ifid_ifinstr_o_23 & (\Reg[18][4]~q  & (!ifid_ifinstr_o_24)))

	.dataa(\Reg[18][4]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(ifid_ifinstr_o_24),
	.datad(\Reg[22][4]~q ),
	.cin(gnd),
	.combout(\Mux27~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~2 .lut_mask = 16'hCEC2;
defparam \Mux27~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N23
dffeas \Reg[30][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][4] .is_wysiwyg = "true";
defparam \Reg[30][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N22
cycloneive_lcell_comb \Mux27~3 (
// Equation(s):
// \Mux27~3_combout  = (\Mux27~2_combout  & (((\Reg[30][4]~q ) # (!ifid_ifinstr_o_24)))) # (!\Mux27~2_combout  & (\Reg[26][4]~q  & ((ifid_ifinstr_o_24))))

	.dataa(\Reg[26][4]~q ),
	.datab(\Mux27~2_combout ),
	.datac(\Reg[30][4]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux27~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~3 .lut_mask = 16'hE2CC;
defparam \Mux27~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N0
cycloneive_lcell_comb \Mux27~6 (
// Equation(s):
// \Mux27~6_combout  = (ifid_ifinstr_o_22 & (((\Mux27~3_combout ) # (ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & (\Mux27~5_combout  & ((!ifid_ifinstr_o_21))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Mux27~5_combout ),
	.datac(\Mux27~3_combout ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux27~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~6 .lut_mask = 16'hAAE4;
defparam \Mux27~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N12
cycloneive_lcell_comb \Reg[23][4]~feeder (
// Equation(s):
// \Reg[23][4]~feeder_combout  = \wdat~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat3),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[23][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[23][4]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[23][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N13
dffeas \Reg[23][4] (
	.clk(!CLK),
	.d(\Reg[23][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][4] .is_wysiwyg = "true";
defparam \Reg[23][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N21
dffeas \Reg[27][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][4] .is_wysiwyg = "true";
defparam \Reg[27][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N19
dffeas \Reg[19][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][4] .is_wysiwyg = "true";
defparam \Reg[19][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N20
cycloneive_lcell_comb \Mux27~7 (
// Equation(s):
// \Mux27~7_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[27][4]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[19][4]~q )))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[27][4]~q ),
	.datad(\Reg[19][4]~q ),
	.cin(gnd),
	.combout(\Mux27~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~7 .lut_mask = 16'hD9C8;
defparam \Mux27~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N3
dffeas \Reg[31][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][4] .is_wysiwyg = "true";
defparam \Reg[31][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N2
cycloneive_lcell_comb \Mux27~8 (
// Equation(s):
// \Mux27~8_combout  = (\Mux27~7_combout  & (((\Reg[31][4]~q ) # (!ifid_ifinstr_o_23)))) # (!\Mux27~7_combout  & (\Reg[23][4]~q  & ((ifid_ifinstr_o_23))))

	.dataa(\Reg[23][4]~q ),
	.datab(\Mux27~7_combout ),
	.datac(\Reg[31][4]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux27~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~8 .lut_mask = 16'hE2CC;
defparam \Mux27~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N3
dffeas \Reg[2][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][4] .is_wysiwyg = "true";
defparam \Reg[2][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N8
cycloneive_lcell_comb \Mux27~15 (
// Equation(s):
// \Mux27~15_combout  = (\Mux27~14_combout ) # ((\Reg[2][4]~q  & (ifid_ifinstr_o_22 & !ifid_ifinstr_o_21)))

	.dataa(\Mux27~14_combout ),
	.datab(\Reg[2][4]~q ),
	.datac(ifid_ifinstr_o_22),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux27~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~15 .lut_mask = 16'hAAEA;
defparam \Mux27~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N9
dffeas \Reg[10][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][4] .is_wysiwyg = "true";
defparam \Reg[10][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N15
dffeas \Reg[8][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][4] .is_wysiwyg = "true";
defparam \Reg[8][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N14
cycloneive_lcell_comb \Mux27~12 (
// Equation(s):
// \Mux27~12_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[10][4]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[8][4]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[10][4]~q ),
	.datac(\Reg[8][4]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux27~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~12 .lut_mask = 16'hEE50;
defparam \Mux27~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N3
dffeas \Reg[11][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][4] .is_wysiwyg = "true";
defparam \Reg[11][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N13
dffeas \Reg[9][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][4] .is_wysiwyg = "true";
defparam \Reg[9][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N2
cycloneive_lcell_comb \Mux27~13 (
// Equation(s):
// \Mux27~13_combout  = (ifid_ifinstr_o_21 & ((\Mux27~12_combout  & (\Reg[11][4]~q )) # (!\Mux27~12_combout  & ((\Reg[9][4]~q ))))) # (!ifid_ifinstr_o_21 & (\Mux27~12_combout ))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux27~12_combout ),
	.datac(\Reg[11][4]~q ),
	.datad(\Reg[9][4]~q ),
	.cin(gnd),
	.combout(\Mux27~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~13 .lut_mask = 16'hE6C4;
defparam \Mux27~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N26
cycloneive_lcell_comb \Mux27~16 (
// Equation(s):
// \Mux27~16_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23) # (\Mux27~13_combout )))) # (!ifid_ifinstr_o_24 & (\Mux27~15_combout  & (!ifid_ifinstr_o_23)))

	.dataa(\Mux27~15_combout ),
	.datab(ifid_ifinstr_o_24),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux27~13_combout ),
	.cin(gnd),
	.combout(\Mux27~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~16 .lut_mask = 16'hCEC2;
defparam \Mux27~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N21
dffeas \Reg[5][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][4] .is_wysiwyg = "true";
defparam \Reg[5][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N19
dffeas \Reg[4][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][4] .is_wysiwyg = "true";
defparam \Reg[4][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N20
cycloneive_lcell_comb \Mux27~10 (
// Equation(s):
// \Mux27~10_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22) # ((\Reg[5][4]~q )))) # (!ifid_ifinstr_o_21 & (!ifid_ifinstr_o_22 & ((\Reg[4][4]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[5][4]~q ),
	.datad(\Reg[4][4]~q ),
	.cin(gnd),
	.combout(\Mux27~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~10 .lut_mask = 16'hB9A8;
defparam \Mux27~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N7
dffeas \Reg[6][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][4] .is_wysiwyg = "true";
defparam \Reg[6][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y39_N21
dffeas \Reg[7][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][4] .is_wysiwyg = "true";
defparam \Reg[7][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N6
cycloneive_lcell_comb \Mux27~11 (
// Equation(s):
// \Mux27~11_combout  = (\Mux27~10_combout  & (((\Reg[7][4]~q )) # (!ifid_ifinstr_o_22))) # (!\Mux27~10_combout  & (ifid_ifinstr_o_22 & (\Reg[6][4]~q )))

	.dataa(\Mux27~10_combout ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[6][4]~q ),
	.datad(\Reg[7][4]~q ),
	.cin(gnd),
	.combout(\Mux27~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~11 .lut_mask = 16'hEA62;
defparam \Mux27~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y37_N1
dffeas \Reg[14][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][4] .is_wysiwyg = "true";
defparam \Reg[14][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y37_N23
dffeas \Reg[15][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][4] .is_wysiwyg = "true";
defparam \Reg[15][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N17
dffeas \Reg[12][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][4] .is_wysiwyg = "true";
defparam \Reg[12][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N19
dffeas \Reg[13][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][4] .is_wysiwyg = "true";
defparam \Reg[13][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N18
cycloneive_lcell_comb \Mux27~17 (
// Equation(s):
// \Mux27~17_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[13][4]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[12][4]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[12][4]~q ),
	.datac(\Reg[13][4]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux27~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~17 .lut_mask = 16'hFA44;
defparam \Mux27~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N22
cycloneive_lcell_comb \Mux27~18 (
// Equation(s):
// \Mux27~18_combout  = (ifid_ifinstr_o_22 & ((\Mux27~17_combout  & ((\Reg[15][4]~q ))) # (!\Mux27~17_combout  & (\Reg[14][4]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux27~17_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[14][4]~q ),
	.datac(\Reg[15][4]~q ),
	.datad(\Mux27~17_combout ),
	.cin(gnd),
	.combout(\Mux27~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~18 .lut_mask = 16'hF588;
defparam \Mux27~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N15
dffeas \Reg[19][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][3] .is_wysiwyg = "true";
defparam \Reg[19][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N5
dffeas \Reg[23][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][3] .is_wysiwyg = "true";
defparam \Reg[23][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N4
cycloneive_lcell_comb \Mux28~7 (
// Equation(s):
// \Mux28~7_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[23][3]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[19][3]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[19][3]~q ),
	.datac(\Reg[23][3]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux28~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~7 .lut_mask = 16'hFA44;
defparam \Mux28~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N31
dffeas \Reg[31][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][3] .is_wysiwyg = "true";
defparam \Reg[31][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N24
cycloneive_lcell_comb \Reg[27][3]~feeder (
// Equation(s):
// \Reg[27][3]~feeder_combout  = \wdat~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat4),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[27][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[27][3]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[27][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N25
dffeas \Reg[27][3] (
	.clk(!CLK),
	.d(\Reg[27][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][3] .is_wysiwyg = "true";
defparam \Reg[27][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N30
cycloneive_lcell_comb \Mux28~8 (
// Equation(s):
// \Mux28~8_combout  = (\Mux28~7_combout  & (((\Reg[31][3]~q )) # (!ifid_ifinstr_o_24))) # (!\Mux28~7_combout  & (ifid_ifinstr_o_24 & ((\Reg[27][3]~q ))))

	.dataa(\Mux28~7_combout ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[31][3]~q ),
	.datad(\Reg[27][3]~q ),
	.cin(gnd),
	.combout(\Mux28~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~8 .lut_mask = 16'hE6A2;
defparam \Mux28~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N3
dffeas \Reg[25][3] (
	.clk(!CLK),
	.d(wdat4),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][3] .is_wysiwyg = "true";
defparam \Reg[25][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N18
cycloneive_lcell_comb \Reg[29][3]~feeder (
// Equation(s):
// \Reg[29][3]~feeder_combout  = \wdat~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat4),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[29][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[29][3]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[29][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N19
dffeas \Reg[29][3] (
	.clk(!CLK),
	.d(\Reg[29][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][3] .is_wysiwyg = "true";
defparam \Reg[29][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y38_N21
dffeas \Reg[21][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][3] .is_wysiwyg = "true";
defparam \Reg[21][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N27
dffeas \Reg[17][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][3] .is_wysiwyg = "true";
defparam \Reg[17][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N20
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & (\Reg[21][3]~q )) # (!ifid_ifinstr_o_23 & ((\Reg[17][3]~q )))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[21][3]~q ),
	.datad(\Reg[17][3]~q ),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'hD9C8;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N8
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// \Mux28~1_combout  = (\Mux28~0_combout  & (((\Reg[29][3]~q ) # (!ifid_ifinstr_o_24)))) # (!\Mux28~0_combout  & (\Reg[25][3]~q  & ((ifid_ifinstr_o_24))))

	.dataa(\Reg[25][3]~q ),
	.datab(\Reg[29][3]~q ),
	.datac(\Mux28~0_combout ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hCAF0;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N12
cycloneive_lcell_comb \Reg[30][3]~feeder (
// Equation(s):
// \Reg[30][3]~feeder_combout  = \wdat~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat4),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[30][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[30][3]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[30][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N13
dffeas \Reg[30][3] (
	.clk(!CLK),
	.d(\Reg[30][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][3] .is_wysiwyg = "true";
defparam \Reg[30][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N7
dffeas \Reg[22][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][3] .is_wysiwyg = "true";
defparam \Reg[22][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N4
cycloneive_lcell_comb \Reg[26][3]~feeder (
// Equation(s):
// \Reg[26][3]~feeder_combout  = \wdat~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat4),
	.cin(gnd),
	.combout(\Reg[26][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[26][3]~feeder .lut_mask = 16'hFF00;
defparam \Reg[26][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N5
dffeas \Reg[26][3] (
	.clk(!CLK),
	.d(\Reg[26][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][3] .is_wysiwyg = "true";
defparam \Reg[26][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N2
cycloneive_lcell_comb \Reg[18][3]~feeder (
// Equation(s):
// \Reg[18][3]~feeder_combout  = \wdat~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat4),
	.cin(gnd),
	.combout(\Reg[18][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[18][3]~feeder .lut_mask = 16'hFF00;
defparam \Reg[18][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N3
dffeas \Reg[18][3] (
	.clk(!CLK),
	.d(\Reg[18][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][3] .is_wysiwyg = "true";
defparam \Reg[18][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N24
cycloneive_lcell_comb \Mux28~2 (
// Equation(s):
// \Mux28~2_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[26][3]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & ((\Reg[18][3]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[26][3]~q ),
	.datad(\Reg[18][3]~q ),
	.cin(gnd),
	.combout(\Mux28~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~2 .lut_mask = 16'hB9A8;
defparam \Mux28~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N6
cycloneive_lcell_comb \Mux28~3 (
// Equation(s):
// \Mux28~3_combout  = (ifid_ifinstr_o_23 & ((\Mux28~2_combout  & (\Reg[30][3]~q )) # (!\Mux28~2_combout  & ((\Reg[22][3]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux28~2_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[30][3]~q ),
	.datac(\Reg[22][3]~q ),
	.datad(\Mux28~2_combout ),
	.cin(gnd),
	.combout(\Mux28~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~3 .lut_mask = 16'hDDA0;
defparam \Mux28~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N7
dffeas \Reg[16][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][3] .is_wysiwyg = "true";
defparam \Reg[16][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N28
cycloneive_lcell_comb \Reg[24][3]~feeder (
// Equation(s):
// \Reg[24][3]~feeder_combout  = \wdat~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat4),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[24][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[24][3]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[24][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N29
dffeas \Reg[24][3] (
	.clk(!CLK),
	.d(\Reg[24][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][3] .is_wysiwyg = "true";
defparam \Reg[24][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N6
cycloneive_lcell_comb \Mux28~4 (
// Equation(s):
// \Mux28~4_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Reg[24][3]~q ))) # (!ifid_ifinstr_o_24 & (\Reg[16][3]~q ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[16][3]~q ),
	.datad(\Reg[24][3]~q ),
	.cin(gnd),
	.combout(\Mux28~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~4 .lut_mask = 16'hDC98;
defparam \Mux28~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N23
dffeas \Reg[20][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][3] .is_wysiwyg = "true";
defparam \Reg[20][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y33_N15
dffeas \Reg[28][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][3] .is_wysiwyg = "true";
defparam \Reg[28][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N30
cycloneive_lcell_comb \Mux28~5 (
// Equation(s):
// \Mux28~5_combout  = (ifid_ifinstr_o_23 & ((\Mux28~4_combout  & ((\Reg[28][3]~q ))) # (!\Mux28~4_combout  & (\Reg[20][3]~q )))) # (!ifid_ifinstr_o_23 & (\Mux28~4_combout ))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux28~4_combout ),
	.datac(\Reg[20][3]~q ),
	.datad(\Reg[28][3]~q ),
	.cin(gnd),
	.combout(\Mux28~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~5 .lut_mask = 16'hEC64;
defparam \Mux28~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N12
cycloneive_lcell_comb \Mux28~6 (
// Equation(s):
// \Mux28~6_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Mux28~3_combout )) # (!ifid_ifinstr_o_22 & ((\Mux28~5_combout )))))

	.dataa(\Mux28~3_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux28~5_combout ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux28~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~6 .lut_mask = 16'hEE30;
defparam \Mux28~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N9
dffeas \Reg[5][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][3] .is_wysiwyg = "true";
defparam \Reg[5][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N27
dffeas \Reg[4][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][3] .is_wysiwyg = "true";
defparam \Reg[4][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N26
cycloneive_lcell_comb \Mux28~12 (
// Equation(s):
// \Mux28~12_combout  = (ifid_ifinstr_o_21 & ((\Reg[5][3]~q ) # ((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & (((\Reg[4][3]~q  & !ifid_ifinstr_o_22))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[5][3]~q ),
	.datac(\Reg[4][3]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux28~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~12 .lut_mask = 16'hAAD8;
defparam \Mux28~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N25
dffeas \Reg[7][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][3] .is_wysiwyg = "true";
defparam \Reg[7][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N24
cycloneive_lcell_comb \Mux28~13 (
// Equation(s):
// \Mux28~13_combout  = (\Mux28~12_combout  & (((\Reg[7][3]~q ) # (!ifid_ifinstr_o_22)))) # (!\Mux28~12_combout  & (\Reg[6][3]~q  & ((ifid_ifinstr_o_22))))

	.dataa(\Reg[6][3]~q ),
	.datab(\Mux28~12_combout ),
	.datac(\Reg[7][3]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux28~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~13 .lut_mask = 16'hE2CC;
defparam \Mux28~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N3
dffeas \Reg[2][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][3] .is_wysiwyg = "true";
defparam \Reg[2][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N2
cycloneive_lcell_comb \Mux28~15 (
// Equation(s):
// \Mux28~15_combout  = (\Mux28~14_combout ) # ((!ifid_ifinstr_o_21 & (\Reg[2][3]~q  & ifid_ifinstr_o_22)))

	.dataa(\Mux28~14_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[2][3]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux28~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~15 .lut_mask = 16'hBAAA;
defparam \Mux28~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N16
cycloneive_lcell_comb \Mux28~16 (
// Equation(s):
// \Mux28~16_combout  = (ifid_ifinstr_o_23 & ((\Mux28~13_combout ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((!ifid_ifinstr_o_24 & \Mux28~15_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux28~13_combout ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Mux28~15_combout ),
	.cin(gnd),
	.combout(\Mux28~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~16 .lut_mask = 16'hADA8;
defparam \Mux28~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N21
dffeas \Reg[13][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][3] .is_wysiwyg = "true";
defparam \Reg[13][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N15
dffeas \Reg[12][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][3] .is_wysiwyg = "true";
defparam \Reg[12][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N14
cycloneive_lcell_comb \Mux28~17 (
// Equation(s):
// \Mux28~17_combout  = (ifid_ifinstr_o_21 & ((\Reg[13][3]~q ) # ((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & (((\Reg[12][3]~q  & !ifid_ifinstr_o_22))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[13][3]~q ),
	.datac(\Reg[12][3]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux28~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~17 .lut_mask = 16'hAAD8;
defparam \Mux28~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N17
dffeas \Reg[14][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][3] .is_wysiwyg = "true";
defparam \Reg[14][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N11
dffeas \Reg[15][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][3] .is_wysiwyg = "true";
defparam \Reg[15][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N10
cycloneive_lcell_comb \Mux28~18 (
// Equation(s):
// \Mux28~18_combout  = (\Mux28~17_combout  & (((\Reg[15][3]~q ) # (!ifid_ifinstr_o_22)))) # (!\Mux28~17_combout  & (\Reg[14][3]~q  & ((ifid_ifinstr_o_22))))

	.dataa(\Mux28~17_combout ),
	.datab(\Reg[14][3]~q ),
	.datac(\Reg[15][3]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux28~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~18 .lut_mask = 16'hE4AA;
defparam \Mux28~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N19
dffeas \Reg[11][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][3] .is_wysiwyg = "true";
defparam \Reg[11][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N9
dffeas \Reg[9][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][3] .is_wysiwyg = "true";
defparam \Reg[9][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N5
dffeas \Reg[10][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][3] .is_wysiwyg = "true";
defparam \Reg[10][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N4
cycloneive_lcell_comb \Mux28~10 (
// Equation(s):
// \Mux28~10_combout  = (ifid_ifinstr_o_22 & (((\Reg[10][3]~q ) # (ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & (\Reg[8][3]~q  & ((!ifid_ifinstr_o_21))))

	.dataa(\Reg[8][3]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[10][3]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux28~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~10 .lut_mask = 16'hCCE2;
defparam \Mux28~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N8
cycloneive_lcell_comb \Mux28~11 (
// Equation(s):
// \Mux28~11_combout  = (ifid_ifinstr_o_21 & ((\Mux28~10_combout  & (\Reg[11][3]~q )) # (!\Mux28~10_combout  & ((\Reg[9][3]~q ))))) # (!ifid_ifinstr_o_21 & (((\Mux28~10_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[11][3]~q ),
	.datac(\Reg[9][3]~q ),
	.datad(\Mux28~10_combout ),
	.cin(gnd),
	.combout(\Mux28~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~11 .lut_mask = 16'hDDA0;
defparam \Mux28~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N12
cycloneive_lcell_comb \Mux61~4 (
// Equation(s):
// \Mux61~4_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[24][2]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[16][2]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[16][2]~q ),
	.datac(\Reg[24][2]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux61~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~4 .lut_mask = 16'hFA44;
defparam \Mux61~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N0
cycloneive_lcell_comb \Mux61~5 (
// Equation(s):
// \Mux61~5_combout  = (ifid_ifinstr_o_18 & ((\Mux61~4_combout  & (\Reg[28][2]~q )) # (!\Mux61~4_combout  & ((\Reg[20][2]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux61~4_combout ))))

	.dataa(\Reg[28][2]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[20][2]~q ),
	.datad(\Mux61~4_combout ),
	.cin(gnd),
	.combout(\Mux61~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~5 .lut_mask = 16'hBBC0;
defparam \Mux61~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N11
dffeas \Reg[30][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat2),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][2] .is_wysiwyg = "true";
defparam \Reg[30][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N10
cycloneive_lcell_comb \Mux61~3 (
// Equation(s):
// \Mux61~3_combout  = (\Mux61~2_combout  & (((\Reg[30][2]~q )) # (!ifid_ifinstr_o_18))) # (!\Mux61~2_combout  & (ifid_ifinstr_o_18 & ((\Reg[22][2]~q ))))

	.dataa(\Mux61~2_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[30][2]~q ),
	.datad(\Reg[22][2]~q ),
	.cin(gnd),
	.combout(\Mux61~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~3 .lut_mask = 16'hE6A2;
defparam \Mux61~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N2
cycloneive_lcell_comb \Mux61~6 (
// Equation(s):
// \Mux61~6_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Mux61~3_combout ))) # (!ifid_ifinstr_o_17 & (\Mux61~5_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux61~5_combout ),
	.datad(\Mux61~3_combout ),
	.cin(gnd),
	.combout(\Mux61~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~6 .lut_mask = 16'hDC98;
defparam \Mux61~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N22
cycloneive_lcell_comb \Mux61~7 (
// Equation(s):
// \Mux61~7_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Reg[23][2]~q ))) # (!ifid_ifinstr_o_18 & (\Reg[19][2]~q ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[19][2]~q ),
	.datad(\Reg[23][2]~q ),
	.cin(gnd),
	.combout(\Mux61~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~7 .lut_mask = 16'hDC98;
defparam \Mux61~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N16
cycloneive_lcell_comb \Mux61~8 (
// Equation(s):
// \Mux61~8_combout  = (ifid_ifinstr_o_19 & ((\Mux61~7_combout  & (\Reg[31][2]~q )) # (!\Mux61~7_combout  & ((\Reg[27][2]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux61~7_combout ))))

	.dataa(\Reg[31][2]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[27][2]~q ),
	.datad(\Mux61~7_combout ),
	.cin(gnd),
	.combout(\Mux61~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~8 .lut_mask = 16'hBBC0;
defparam \Mux61~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N24
cycloneive_lcell_comb \Mux61~0 (
// Equation(s):
// \Mux61~0_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19) # (\Reg[21][2]~q )))) # (!ifid_ifinstr_o_18 & (\Reg[17][2]~q  & (!ifid_ifinstr_o_19)))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[17][2]~q ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Reg[21][2]~q ),
	.cin(gnd),
	.combout(\Mux61~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~0 .lut_mask = 16'hAEA4;
defparam \Mux61~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N10
cycloneive_lcell_comb \Reg[25][2]~feeder (
// Equation(s):
// \Reg[25][2]~feeder_combout  = \wdat~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat2),
	.cin(gnd),
	.combout(\Reg[25][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][2]~feeder .lut_mask = 16'hFF00;
defparam \Reg[25][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N11
dffeas \Reg[25][2] (
	.clk(!CLK),
	.d(\Reg[25][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][2] .is_wysiwyg = "true";
defparam \Reg[25][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N18
cycloneive_lcell_comb \Mux61~1 (
// Equation(s):
// \Mux61~1_combout  = (\Mux61~0_combout  & ((\Reg[29][2]~q ) # ((!ifid_ifinstr_o_19)))) # (!\Mux61~0_combout  & (((ifid_ifinstr_o_19 & \Reg[25][2]~q ))))

	.dataa(\Reg[29][2]~q ),
	.datab(\Mux61~0_combout ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Reg[25][2]~q ),
	.cin(gnd),
	.combout(\Mux61~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~1 .lut_mask = 16'hBC8C;
defparam \Mux61~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N24
cycloneive_lcell_comb \Mux61~10 (
// Equation(s):
// \Mux61~10_combout  = (ifid_ifinstr_o_16 & (((ifid_ifinstr_o_17)))) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[10][2]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[8][2]~q ))))

	.dataa(\Reg[8][2]~q ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[10][2]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux61~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~10 .lut_mask = 16'hFC22;
defparam \Mux61~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N24
cycloneive_lcell_comb \Mux61~11 (
// Equation(s):
// \Mux61~11_combout  = (ifid_ifinstr_o_16 & ((\Mux61~10_combout  & ((\Reg[11][2]~q ))) # (!\Mux61~10_combout  & (\Reg[9][2]~q )))) # (!ifid_ifinstr_o_16 & (\Mux61~10_combout ))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux61~10_combout ),
	.datac(\Reg[9][2]~q ),
	.datad(\Reg[11][2]~q ),
	.cin(gnd),
	.combout(\Mux61~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~11 .lut_mask = 16'hEC64;
defparam \Mux61~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N2
cycloneive_lcell_comb \Mux61~17 (
// Equation(s):
// \Mux61~17_combout  = (ifid_ifinstr_o_16 & (((\Reg[13][2]~q ) # (ifid_ifinstr_o_17)))) # (!ifid_ifinstr_o_16 & (\Reg[12][2]~q  & ((!ifid_ifinstr_o_17))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[12][2]~q ),
	.datac(\Reg[13][2]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux61~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~17 .lut_mask = 16'hAAE4;
defparam \Mux61~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N12
cycloneive_lcell_comb \Mux61~18 (
// Equation(s):
// \Mux61~18_combout  = (\Mux61~17_combout  & (((\Reg[15][2]~q )) # (!ifid_ifinstr_o_17))) # (!\Mux61~17_combout  & (ifid_ifinstr_o_17 & (\Reg[14][2]~q )))

	.dataa(\Mux61~17_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[14][2]~q ),
	.datad(\Reg[15][2]~q ),
	.cin(gnd),
	.combout(\Mux61~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~18 .lut_mask = 16'hEA62;
defparam \Mux61~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N30
cycloneive_lcell_comb \Reg[1][2]~feeder (
// Equation(s):
// \Reg[1][2]~feeder_combout  = \wdat~5_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat2),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[1][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[1][2]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[1][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y36_N31
dffeas \Reg[1][2] (
	.clk(!CLK),
	.d(\Reg[1][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][2] .is_wysiwyg = "true";
defparam \Reg[1][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N20
cycloneive_lcell_comb \Mux61~14 (
// Equation(s):
// \Mux61~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[3][2]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[1][2]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[1][2]~q ),
	.datad(\Reg[3][2]~q ),
	.cin(gnd),
	.combout(\Mux61~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~14 .lut_mask = 16'hC840;
defparam \Mux61~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N30
cycloneive_lcell_comb \Mux61~15 (
// Equation(s):
// \Mux61~15_combout  = (\Mux61~14_combout ) # ((\Reg[2][2]~q  & (ifid_ifinstr_o_17 & !ifid_ifinstr_o_16)))

	.dataa(\Reg[2][2]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux61~14_combout ),
	.cin(gnd),
	.combout(\Mux61~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~15 .lut_mask = 16'hFF08;
defparam \Mux61~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N22
cycloneive_lcell_comb \Mux61~13 (
// Equation(s):
// \Mux61~13_combout  = (\Mux61~12_combout  & (((\Reg[7][2]~q )) # (!ifid_ifinstr_o_17))) # (!\Mux61~12_combout  & (ifid_ifinstr_o_17 & ((\Reg[6][2]~q ))))

	.dataa(\Mux61~12_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[7][2]~q ),
	.datad(\Reg[6][2]~q ),
	.cin(gnd),
	.combout(\Mux61~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~13 .lut_mask = 16'hE6A2;
defparam \Mux61~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N10
cycloneive_lcell_comb \Mux61~16 (
// Equation(s):
// \Mux61~16_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Mux61~13_combout ))) # (!ifid_ifinstr_o_18 & (\Mux61~15_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Mux61~15_combout ),
	.datad(\Mux61~13_combout ),
	.cin(gnd),
	.combout(\Mux61~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~16 .lut_mask = 16'hDC98;
defparam \Mux61~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N15
dffeas \Reg[30][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][8] .is_wysiwyg = "true";
defparam \Reg[30][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N9
dffeas \Reg[26][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][8] .is_wysiwyg = "true";
defparam \Reg[26][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N0
cycloneive_lcell_comb \Reg[18][8]~feeder (
// Equation(s):
// \Reg[18][8]~feeder_combout  = \wdat~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat5),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[18][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[18][8]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[18][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N1
dffeas \Reg[18][8] (
	.clk(!CLK),
	.d(\Reg[18][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][8] .is_wysiwyg = "true";
defparam \Reg[18][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y30_N21
dffeas \Reg[22][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][8] .is_wysiwyg = "true";
defparam \Reg[22][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N20
cycloneive_lcell_comb \Mux23~2 (
// Equation(s):
// \Mux23~2_combout  = (ifid_ifinstr_o_23 & (((\Reg[22][8]~q ) # (ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (\Reg[18][8]~q  & ((!ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[18][8]~q ),
	.datac(\Reg[22][8]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux23~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~2 .lut_mask = 16'hAAE4;
defparam \Mux23~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N8
cycloneive_lcell_comb \Mux23~3 (
// Equation(s):
// \Mux23~3_combout  = (ifid_ifinstr_o_24 & ((\Mux23~2_combout  & (\Reg[30][8]~q )) # (!\Mux23~2_combout  & ((\Reg[26][8]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux23~2_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[30][8]~q ),
	.datac(\Reg[26][8]~q ),
	.datad(\Mux23~2_combout ),
	.cin(gnd),
	.combout(\Mux23~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~3 .lut_mask = 16'hDDA0;
defparam \Mux23~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N29
dffeas \Reg[24][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][8] .is_wysiwyg = "true";
defparam \Reg[24][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y33_N19
dffeas \Reg[16][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][8] .is_wysiwyg = "true";
defparam \Reg[16][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N30
cycloneive_lcell_comb \Reg[20][8]~feeder (
// Equation(s):
// \Reg[20][8]~feeder_combout  = \wdat~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat5),
	.cin(gnd),
	.combout(\Reg[20][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[20][8]~feeder .lut_mask = 16'hFF00;
defparam \Reg[20][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N31
dffeas \Reg[20][8] (
	.clk(!CLK),
	.d(\Reg[20][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][8] .is_wysiwyg = "true";
defparam \Reg[20][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N18
cycloneive_lcell_comb \Mux23~4 (
// Equation(s):
// \Mux23~4_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[20][8]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[16][8]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[16][8]~q ),
	.datad(\Reg[20][8]~q ),
	.cin(gnd),
	.combout(\Mux23~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~4 .lut_mask = 16'hDC98;
defparam \Mux23~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N18
cycloneive_lcell_comb \Mux23~5 (
// Equation(s):
// \Mux23~5_combout  = (\Mux23~4_combout  & ((\Reg[28][8]~q ) # ((!ifid_ifinstr_o_24)))) # (!\Mux23~4_combout  & (((\Reg[24][8]~q  & ifid_ifinstr_o_24))))

	.dataa(\Reg[28][8]~q ),
	.datab(\Reg[24][8]~q ),
	.datac(\Mux23~4_combout ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux23~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~5 .lut_mask = 16'hACF0;
defparam \Mux23~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N28
cycloneive_lcell_comb \Mux23~6 (
// Equation(s):
// \Mux23~6_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Mux23~3_combout )) # (!ifid_ifinstr_o_22 & ((\Mux23~5_combout )))))

	.dataa(\Mux23~3_combout ),
	.datab(\Mux23~5_combout ),
	.datac(ifid_ifinstr_o_21),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux23~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~6 .lut_mask = 16'hFA0C;
defparam \Mux23~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N21
dffeas \Reg[23][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][8] .is_wysiwyg = "true";
defparam \Reg[23][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N27
dffeas \Reg[31][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][8] .is_wysiwyg = "true";
defparam \Reg[31][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N5
dffeas \Reg[27][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][8] .is_wysiwyg = "true";
defparam \Reg[27][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N4
cycloneive_lcell_comb \Mux23~7 (
// Equation(s):
// \Mux23~7_combout  = (ifid_ifinstr_o_24 & (((\Reg[27][8]~q ) # (ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & (\Reg[19][8]~q  & ((!ifid_ifinstr_o_23))))

	.dataa(\Reg[19][8]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[27][8]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux23~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~7 .lut_mask = 16'hCCE2;
defparam \Mux23~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N26
cycloneive_lcell_comb \Mux23~8 (
// Equation(s):
// \Mux23~8_combout  = (ifid_ifinstr_o_23 & ((\Mux23~7_combout  & ((\Reg[31][8]~q ))) # (!\Mux23~7_combout  & (\Reg[23][8]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux23~7_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[23][8]~q ),
	.datac(\Reg[31][8]~q ),
	.datad(\Mux23~7_combout ),
	.cin(gnd),
	.combout(\Mux23~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~8 .lut_mask = 16'hF588;
defparam \Mux23~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N2
cycloneive_lcell_comb \Reg[21][8]~feeder (
// Equation(s):
// \Reg[21][8]~feeder_combout  = \wdat~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat5),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[21][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[21][8]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[21][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y37_N3
dffeas \Reg[21][8] (
	.clk(!CLK),
	.d(\Reg[21][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][8] .is_wysiwyg = "true";
defparam \Reg[21][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N20
cycloneive_lcell_comb \Reg[25][8]~feeder (
// Equation(s):
// \Reg[25][8]~feeder_combout  = \wdat~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat5),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[25][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][8]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[25][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y30_N21
dffeas \Reg[25][8] (
	.clk(!CLK),
	.d(\Reg[25][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][8] .is_wysiwyg = "true";
defparam \Reg[25][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N20
cycloneive_lcell_comb \Reg[17][8]~feeder (
// Equation(s):
// \Reg[17][8]~feeder_combout  = \wdat~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat5),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[17][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[17][8]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[17][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N21
dffeas \Reg[17][8] (
	.clk(!CLK),
	.d(\Reg[17][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][8] .is_wysiwyg = "true";
defparam \Reg[17][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N14
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// \Mux23~0_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[25][8]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[17][8]~q )))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[25][8]~q ),
	.datac(\Reg[17][8]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hEE50;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N16
cycloneive_lcell_comb \Reg[29][8]~feeder (
// Equation(s):
// \Reg[29][8]~feeder_combout  = \wdat~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat5),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[29][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[29][8]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[29][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N17
dffeas \Reg[29][8] (
	.clk(!CLK),
	.d(\Reg[29][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][8] .is_wysiwyg = "true";
defparam \Reg[29][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N16
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// \Mux23~1_combout  = (ifid_ifinstr_o_23 & ((\Mux23~0_combout  & ((\Reg[29][8]~q ))) # (!\Mux23~0_combout  & (\Reg[21][8]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux23~0_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[21][8]~q ),
	.datac(\Mux23~0_combout ),
	.datad(\Reg[29][8]~q ),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'hF858;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N7
dffeas \Reg[7][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][8] .is_wysiwyg = "true";
defparam \Reg[7][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y39_N29
dffeas \Reg[6][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][8] .is_wysiwyg = "true";
defparam \Reg[6][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N29
dffeas \Reg[5][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][8] .is_wysiwyg = "true";
defparam \Reg[5][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N23
dffeas \Reg[4][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][8] .is_wysiwyg = "true";
defparam \Reg[4][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N28
cycloneive_lcell_comb \Mux23~10 (
// Equation(s):
// \Mux23~10_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[5][8]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[4][8]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[5][8]~q ),
	.datad(\Reg[4][8]~q ),
	.cin(gnd),
	.combout(\Mux23~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~10 .lut_mask = 16'hD9C8;
defparam \Mux23~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N28
cycloneive_lcell_comb \Mux23~11 (
// Equation(s):
// \Mux23~11_combout  = (ifid_ifinstr_o_22 & ((\Mux23~10_combout  & (\Reg[7][8]~q )) # (!\Mux23~10_combout  & ((\Reg[6][8]~q ))))) # (!ifid_ifinstr_o_22 & (((\Mux23~10_combout ))))

	.dataa(\Reg[7][8]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[6][8]~q ),
	.datad(\Mux23~10_combout ),
	.cin(gnd),
	.combout(\Mux23~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~11 .lut_mask = 16'hBBC0;
defparam \Mux23~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N23
dffeas \Reg[12][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][8] .is_wysiwyg = "true";
defparam \Reg[12][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N24
cycloneive_lcell_comb \Reg[13][8]~feeder (
// Equation(s):
// \Reg[13][8]~feeder_combout  = \wdat~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat5),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[13][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[13][8]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[13][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N25
dffeas \Reg[13][8] (
	.clk(!CLK),
	.d(\Reg[13][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][8] .is_wysiwyg = "true";
defparam \Reg[13][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N0
cycloneive_lcell_comb \Mux23~17 (
// Equation(s):
// \Mux23~17_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22) # ((\Reg[13][8]~q )))) # (!ifid_ifinstr_o_21 & (!ifid_ifinstr_o_22 & (\Reg[12][8]~q )))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[12][8]~q ),
	.datad(\Reg[13][8]~q ),
	.cin(gnd),
	.combout(\Mux23~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~17 .lut_mask = 16'hBA98;
defparam \Mux23~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y37_N27
dffeas \Reg[15][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][8] .is_wysiwyg = "true";
defparam \Reg[15][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y37_N29
dffeas \Reg[14][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][8] .is_wysiwyg = "true";
defparam \Reg[14][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N26
cycloneive_lcell_comb \Mux23~18 (
// Equation(s):
// \Mux23~18_combout  = (ifid_ifinstr_o_22 & ((\Mux23~17_combout  & (\Reg[15][8]~q )) # (!\Mux23~17_combout  & ((\Reg[14][8]~q ))))) # (!ifid_ifinstr_o_22 & (\Mux23~17_combout ))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Mux23~17_combout ),
	.datac(\Reg[15][8]~q ),
	.datad(\Reg[14][8]~q ),
	.cin(gnd),
	.combout(\Mux23~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~18 .lut_mask = 16'hE6C4;
defparam \Mux23~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y31_N29
dffeas \Reg[11][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][8] .is_wysiwyg = "true";
defparam \Reg[11][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N5
dffeas \Reg[10][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][8] .is_wysiwyg = "true";
defparam \Reg[10][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N27
dffeas \Reg[8][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][8] .is_wysiwyg = "true";
defparam \Reg[8][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N26
cycloneive_lcell_comb \Mux23~12 (
// Equation(s):
// \Mux23~12_combout  = (ifid_ifinstr_o_22 & ((\Reg[10][8]~q ) # ((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & (((\Reg[8][8]~q  & !ifid_ifinstr_o_21))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[10][8]~q ),
	.datac(\Reg[8][8]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux23~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~12 .lut_mask = 16'hAAD8;
defparam \Mux23~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N2
cycloneive_lcell_comb \Mux23~13 (
// Equation(s):
// \Mux23~13_combout  = (\Mux23~12_combout  & (((\Reg[11][8]~q ) # (!ifid_ifinstr_o_21)))) # (!\Mux23~12_combout  & (\Reg[9][8]~q  & ((ifid_ifinstr_o_21))))

	.dataa(\Reg[9][8]~q ),
	.datab(\Reg[11][8]~q ),
	.datac(\Mux23~12_combout ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux23~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~13 .lut_mask = 16'hCAF0;
defparam \Mux23~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y31_N1
dffeas \Reg[2][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][8] .is_wysiwyg = "true";
defparam \Reg[2][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N31
dffeas \Reg[1][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][8] .is_wysiwyg = "true";
defparam \Reg[1][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N5
dffeas \Reg[3][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][8] .is_wysiwyg = "true";
defparam \Reg[3][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N30
cycloneive_lcell_comb \Mux23~14 (
// Equation(s):
// \Mux23~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][8]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][8]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[1][8]~q ),
	.datad(\Reg[3][8]~q ),
	.cin(gnd),
	.combout(\Mux23~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~14 .lut_mask = 16'hC840;
defparam \Mux23~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N10
cycloneive_lcell_comb \Mux23~15 (
// Equation(s):
// \Mux23~15_combout  = (\Mux23~14_combout ) # ((ifid_ifinstr_o_22 & (\Reg[2][8]~q  & !ifid_ifinstr_o_21)))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[2][8]~q ),
	.datac(\Mux23~14_combout ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux23~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~15 .lut_mask = 16'hF0F8;
defparam \Mux23~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N28
cycloneive_lcell_comb \Mux23~16 (
// Equation(s):
// \Mux23~16_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Mux23~13_combout )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & ((\Mux23~15_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Mux23~13_combout ),
	.datad(\Mux23~15_combout ),
	.cin(gnd),
	.combout(\Mux23~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~16 .lut_mask = 16'hB9A8;
defparam \Mux23~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N14
cycloneive_lcell_comb \Reg[31][7]~feeder (
// Equation(s):
// \Reg[31][7]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat6),
	.cin(gnd),
	.combout(\Reg[31][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[31][7]~feeder .lut_mask = 16'hFF00;
defparam \Reg[31][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y29_N15
dffeas \Reg[31][7] (
	.clk(!CLK),
	.d(\Reg[31][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][7] .is_wysiwyg = "true";
defparam \Reg[31][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N13
dffeas \Reg[19][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][7] .is_wysiwyg = "true";
defparam \Reg[19][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N19
dffeas \Reg[23][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][7] .is_wysiwyg = "true";
defparam \Reg[23][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N12
cycloneive_lcell_comb \Mux24~7 (
// Equation(s):
// \Mux24~7_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[23][7]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[19][7]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[19][7]~q ),
	.datad(\Reg[23][7]~q ),
	.cin(gnd),
	.combout(\Mux24~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~7 .lut_mask = 16'hDC98;
defparam \Mux24~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N0
cycloneive_lcell_comb \Reg[27][7]~feeder (
// Equation(s):
// \Reg[27][7]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat6),
	.cin(gnd),
	.combout(\Reg[27][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[27][7]~feeder .lut_mask = 16'hFF00;
defparam \Reg[27][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y29_N1
dffeas \Reg[27][7] (
	.clk(!CLK),
	.d(\Reg[27][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][7] .is_wysiwyg = "true";
defparam \Reg[27][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N4
cycloneive_lcell_comb \Mux24~8 (
// Equation(s):
// \Mux24~8_combout  = (ifid_ifinstr_o_24 & ((\Mux24~7_combout  & (\Reg[31][7]~q )) # (!\Mux24~7_combout  & ((\Reg[27][7]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux24~7_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[31][7]~q ),
	.datac(\Mux24~7_combout ),
	.datad(\Reg[27][7]~q ),
	.cin(gnd),
	.combout(\Mux24~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~8 .lut_mask = 16'hDAD0;
defparam \Mux24~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y38_N1
dffeas \Reg[25][7] (
	.clk(!CLK),
	.d(wdat6),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][7] .is_wysiwyg = "true";
defparam \Reg[25][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N11
dffeas \Reg[17][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][7] .is_wysiwyg = "true";
defparam \Reg[17][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N26
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (ifid_ifinstr_o_23 & ((\Reg[21][7]~q ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((\Reg[17][7]~q  & !ifid_ifinstr_o_24))))

	.dataa(\Reg[21][7]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[17][7]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'hCCB8;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N16
cycloneive_lcell_comb \Reg[29][7]~feeder (
// Equation(s):
// \Reg[29][7]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat6),
	.cin(gnd),
	.combout(\Reg[29][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[29][7]~feeder .lut_mask = 16'hFF00;
defparam \Reg[29][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y38_N17
dffeas \Reg[29][7] (
	.clk(!CLK),
	.d(\Reg[29][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][7] .is_wysiwyg = "true";
defparam \Reg[29][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N18
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// \Mux24~1_combout  = (ifid_ifinstr_o_24 & ((\Mux24~0_combout  & ((\Reg[29][7]~q ))) # (!\Mux24~0_combout  & (\Reg[25][7]~q )))) # (!ifid_ifinstr_o_24 & (((\Mux24~0_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[25][7]~q ),
	.datac(\Mux24~0_combout ),
	.datad(\Reg[29][7]~q ),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'hF858;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N3
dffeas \Reg[28][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][7] .is_wysiwyg = "true";
defparam \Reg[28][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y33_N29
dffeas \Reg[20][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][7] .is_wysiwyg = "true";
defparam \Reg[20][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N2
cycloneive_lcell_comb \Mux24~5 (
// Equation(s):
// \Mux24~5_combout  = (\Mux24~4_combout  & (((\Reg[28][7]~q )) # (!ifid_ifinstr_o_23))) # (!\Mux24~4_combout  & (ifid_ifinstr_o_23 & ((\Reg[20][7]~q ))))

	.dataa(\Mux24~4_combout ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[28][7]~q ),
	.datad(\Reg[20][7]~q ),
	.cin(gnd),
	.combout(\Mux24~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~5 .lut_mask = 16'hE6A2;
defparam \Mux24~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N13
dffeas \Reg[18][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][7] .is_wysiwyg = "true";
defparam \Reg[18][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y30_N21
dffeas \Reg[26][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][7] .is_wysiwyg = "true";
defparam \Reg[26][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N20
cycloneive_lcell_comb \Mux24~2 (
// Equation(s):
// \Mux24~2_combout  = (ifid_ifinstr_o_24 & (((\Reg[26][7]~q ) # (ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & (\Reg[18][7]~q  & ((!ifid_ifinstr_o_23))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[18][7]~q ),
	.datac(\Reg[26][7]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux24~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~2 .lut_mask = 16'hAAE4;
defparam \Mux24~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N5
dffeas \Reg[22][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][7] .is_wysiwyg = "true";
defparam \Reg[22][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N4
cycloneive_lcell_comb \Mux24~3 (
// Equation(s):
// \Mux24~3_combout  = (\Mux24~2_combout  & ((\Reg[30][7]~q ) # ((!ifid_ifinstr_o_23)))) # (!\Mux24~2_combout  & (((\Reg[22][7]~q  & ifid_ifinstr_o_23))))

	.dataa(\Reg[30][7]~q ),
	.datab(\Mux24~2_combout ),
	.datac(\Reg[22][7]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux24~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~3 .lut_mask = 16'hB8CC;
defparam \Mux24~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N24
cycloneive_lcell_comb \Mux24~6 (
// Equation(s):
// \Mux24~6_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Mux24~3_combout ))) # (!ifid_ifinstr_o_22 & (\Mux24~5_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux24~5_combout ),
	.datac(\Mux24~3_combout ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux24~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~6 .lut_mask = 16'hFA44;
defparam \Mux24~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y31_N25
dffeas \Reg[2][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][7] .is_wysiwyg = "true";
defparam \Reg[2][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N19
dffeas \Reg[1][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][7] .is_wysiwyg = "true";
defparam \Reg[1][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N25
dffeas \Reg[3][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][7] .is_wysiwyg = "true";
defparam \Reg[3][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N18
cycloneive_lcell_comb \Mux24~14 (
// Equation(s):
// \Mux24~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][7]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][7]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[1][7]~q ),
	.datad(\Reg[3][7]~q ),
	.cin(gnd),
	.combout(\Mux24~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~14 .lut_mask = 16'hC840;
defparam \Mux24~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N4
cycloneive_lcell_comb \Mux24~15 (
// Equation(s):
// \Mux24~15_combout  = (\Mux24~14_combout ) # ((ifid_ifinstr_o_22 & (\Reg[2][7]~q  & !ifid_ifinstr_o_21)))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[2][7]~q ),
	.datac(ifid_ifinstr_o_21),
	.datad(\Mux24~14_combout ),
	.cin(gnd),
	.combout(\Mux24~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~15 .lut_mask = 16'hFF08;
defparam \Mux24~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N9
dffeas \Reg[6][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][7] .is_wysiwyg = "true";
defparam \Reg[6][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y39_N15
dffeas \Reg[7][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][7] .is_wysiwyg = "true";
defparam \Reg[7][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N14
cycloneive_lcell_comb \Mux24~13 (
// Equation(s):
// \Mux24~13_combout  = (\Mux24~12_combout  & (((\Reg[7][7]~q ) # (!ifid_ifinstr_o_22)))) # (!\Mux24~12_combout  & (\Reg[6][7]~q  & ((ifid_ifinstr_o_22))))

	.dataa(\Mux24~12_combout ),
	.datab(\Reg[6][7]~q ),
	.datac(\Reg[7][7]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux24~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~13 .lut_mask = 16'hE4AA;
defparam \Mux24~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N6
cycloneive_lcell_comb \Mux24~16 (
// Equation(s):
// \Mux24~16_combout  = (ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24) # ((\Mux24~13_combout )))) # (!ifid_ifinstr_o_23 & (!ifid_ifinstr_o_24 & (\Mux24~15_combout )))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Mux24~15_combout ),
	.datad(\Mux24~13_combout ),
	.cin(gnd),
	.combout(\Mux24~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~16 .lut_mask = 16'hBA98;
defparam \Mux24~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y37_N9
dffeas \Reg[14][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][7] .is_wysiwyg = "true";
defparam \Reg[14][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y37_N19
dffeas \Reg[15][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][7] .is_wysiwyg = "true";
defparam \Reg[15][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N5
dffeas \Reg[13][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][7] .is_wysiwyg = "true";
defparam \Reg[13][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N4
cycloneive_lcell_comb \Mux24~17 (
// Equation(s):
// \Mux24~17_combout  = (ifid_ifinstr_o_21 & (((\Reg[13][7]~q ) # (ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & (\Reg[12][7]~q  & ((!ifid_ifinstr_o_22))))

	.dataa(\Reg[12][7]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[13][7]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux24~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~17 .lut_mask = 16'hCCE2;
defparam \Mux24~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N18
cycloneive_lcell_comb \Mux24~18 (
// Equation(s):
// \Mux24~18_combout  = (ifid_ifinstr_o_22 & ((\Mux24~17_combout  & ((\Reg[15][7]~q ))) # (!\Mux24~17_combout  & (\Reg[14][7]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux24~17_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[14][7]~q ),
	.datac(\Reg[15][7]~q ),
	.datad(\Mux24~17_combout ),
	.cin(gnd),
	.combout(\Mux24~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~18 .lut_mask = 16'hF588;
defparam \Mux24~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N22
cycloneive_lcell_comb \Reg[9][7]~feeder (
// Equation(s):
// \Reg[9][7]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat6),
	.cin(gnd),
	.combout(\Reg[9][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[9][7]~feeder .lut_mask = 16'hFF00;
defparam \Reg[9][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N23
dffeas \Reg[9][7] (
	.clk(!CLK),
	.d(\Reg[9][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][7] .is_wysiwyg = "true";
defparam \Reg[9][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N4
cycloneive_lcell_comb \Reg[11][7]~feeder (
// Equation(s):
// \Reg[11][7]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat6),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[11][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[11][7]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[11][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y31_N5
dffeas \Reg[11][7] (
	.clk(!CLK),
	.d(\Reg[11][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][7] .is_wysiwyg = "true";
defparam \Reg[11][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N25
dffeas \Reg[10][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][7] .is_wysiwyg = "true";
defparam \Reg[10][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N24
cycloneive_lcell_comb \Mux24~10 (
// Equation(s):
// \Mux24~10_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[10][7]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[8][7]~q ))))

	.dataa(\Reg[8][7]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[10][7]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux24~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~10 .lut_mask = 16'hFC22;
defparam \Mux24~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N30
cycloneive_lcell_comb \Mux24~11 (
// Equation(s):
// \Mux24~11_combout  = (ifid_ifinstr_o_21 & ((\Mux24~10_combout  & ((\Reg[11][7]~q ))) # (!\Mux24~10_combout  & (\Reg[9][7]~q )))) # (!ifid_ifinstr_o_21 & (((\Mux24~10_combout ))))

	.dataa(\Reg[9][7]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[11][7]~q ),
	.datad(\Mux24~10_combout ),
	.cin(gnd),
	.combout(\Mux24~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~11 .lut_mask = 16'hF388;
defparam \Mux24~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N4
cycloneive_lcell_comb \Reg[24][6]~feeder (
// Equation(s):
// \Reg[24][6]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat7),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[24][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[24][6]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[24][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N5
dffeas \Reg[24][6] (
	.clk(!CLK),
	.d(\Reg[24][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][6] .is_wysiwyg = "true";
defparam \Reg[24][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N27
dffeas \Reg[28][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][6] .is_wysiwyg = "true";
defparam \Reg[28][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y33_N27
dffeas \Reg[20][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][6] .is_wysiwyg = "true";
defparam \Reg[20][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y33_N9
dffeas \Reg[16][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][6] .is_wysiwyg = "true";
defparam \Reg[16][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N26
cycloneive_lcell_comb \Mux25~4 (
// Equation(s):
// \Mux25~4_combout  = (ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24) # ((\Reg[20][6]~q )))) # (!ifid_ifinstr_o_23 & (!ifid_ifinstr_o_24 & ((\Reg[16][6]~q ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[20][6]~q ),
	.datad(\Reg[16][6]~q ),
	.cin(gnd),
	.combout(\Mux25~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~4 .lut_mask = 16'hB9A8;
defparam \Mux25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N26
cycloneive_lcell_comb \Mux25~5 (
// Equation(s):
// \Mux25~5_combout  = (ifid_ifinstr_o_24 & ((\Mux25~4_combout  & ((\Reg[28][6]~q ))) # (!\Mux25~4_combout  & (\Reg[24][6]~q )))) # (!ifid_ifinstr_o_24 & (((\Mux25~4_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[24][6]~q ),
	.datac(\Reg[28][6]~q ),
	.datad(\Mux25~4_combout ),
	.cin(gnd),
	.combout(\Mux25~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~5 .lut_mask = 16'hF588;
defparam \Mux25~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N3
dffeas \Reg[26][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][6] .is_wysiwyg = "true";
defparam \Reg[26][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y33_N21
dffeas \Reg[18][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][6] .is_wysiwyg = "true";
defparam \Reg[18][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N0
cycloneive_lcell_comb \Reg[22][6]~feeder (
// Equation(s):
// \Reg[22][6]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat7),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[22][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[22][6]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[22][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N1
dffeas \Reg[22][6] (
	.clk(!CLK),
	.d(\Reg[22][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][6] .is_wysiwyg = "true";
defparam \Reg[22][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N20
cycloneive_lcell_comb \Mux25~2 (
// Equation(s):
// \Mux25~2_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[22][6]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[18][6]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[18][6]~q ),
	.datad(\Reg[22][6]~q ),
	.cin(gnd),
	.combout(\Mux25~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~2 .lut_mask = 16'hDC98;
defparam \Mux25~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N24
cycloneive_lcell_comb \Mux25~3 (
// Equation(s):
// \Mux25~3_combout  = (ifid_ifinstr_o_24 & ((\Mux25~2_combout  & (\Reg[30][6]~q )) # (!\Mux25~2_combout  & ((\Reg[26][6]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux25~2_combout ))))

	.dataa(\Reg[30][6]~q ),
	.datab(\Reg[26][6]~q ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Mux25~2_combout ),
	.cin(gnd),
	.combout(\Mux25~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~3 .lut_mask = 16'hAFC0;
defparam \Mux25~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N26
cycloneive_lcell_comb \Mux25~6 (
// Equation(s):
// \Mux25~6_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Mux25~3_combout ))) # (!ifid_ifinstr_o_22 & (\Mux25~5_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux25~5_combout ),
	.datac(ifid_ifinstr_o_22),
	.datad(\Mux25~3_combout ),
	.cin(gnd),
	.combout(\Mux25~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~6 .lut_mask = 16'hF4A4;
defparam \Mux25~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N0
cycloneive_lcell_comb \Reg[21][6]~feeder (
// Equation(s):
// \Reg[21][6]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat7),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[21][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[21][6]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[21][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y36_N1
dffeas \Reg[21][6] (
	.clk(!CLK),
	.d(\Reg[21][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][6] .is_wysiwyg = "true";
defparam \Reg[21][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N0
cycloneive_lcell_comb \Reg[25][6]~feeder (
// Equation(s):
// \Reg[25][6]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat7),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[25][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][6]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[25][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N1
dffeas \Reg[25][6] (
	.clk(!CLK),
	.d(\Reg[25][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][6] .is_wysiwyg = "true";
defparam \Reg[25][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N26
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Reg[25][6]~q ))) # (!ifid_ifinstr_o_24 & (\Reg[17][6]~q ))))

	.dataa(\Reg[17][6]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(ifid_ifinstr_o_24),
	.datad(\Reg[25][6]~q ),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hF2C2;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N2
cycloneive_lcell_comb \Reg[29][6]~feeder (
// Equation(s):
// \Reg[29][6]~feeder_combout  = \wdat~15_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat7),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[29][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[29][6]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[29][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N3
dffeas \Reg[29][6] (
	.clk(!CLK),
	.d(\Reg[29][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][6] .is_wysiwyg = "true";
defparam \Reg[29][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N24
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// \Mux25~1_combout  = (\Mux25~0_combout  & (((\Reg[29][6]~q ) # (!ifid_ifinstr_o_23)))) # (!\Mux25~0_combout  & (\Reg[21][6]~q  & (ifid_ifinstr_o_23)))

	.dataa(\Reg[21][6]~q ),
	.datab(\Mux25~0_combout ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Reg[29][6]~q ),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hEC2C;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N3
dffeas \Reg[23][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][6] .is_wysiwyg = "true";
defparam \Reg[23][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N25
dffeas \Reg[19][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][6] .is_wysiwyg = "true";
defparam \Reg[19][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N9
dffeas \Reg[27][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][6] .is_wysiwyg = "true";
defparam \Reg[27][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N24
cycloneive_lcell_comb \Mux25~7 (
// Equation(s):
// \Mux25~7_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[27][6]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & (\Reg[19][6]~q )))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[19][6]~q ),
	.datad(\Reg[27][6]~q ),
	.cin(gnd),
	.combout(\Mux25~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~7 .lut_mask = 16'hBA98;
defparam \Mux25~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N23
dffeas \Reg[31][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][6] .is_wysiwyg = "true";
defparam \Reg[31][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N22
cycloneive_lcell_comb \Mux25~8 (
// Equation(s):
// \Mux25~8_combout  = (\Mux25~7_combout  & (((\Reg[31][6]~q ) # (!ifid_ifinstr_o_23)))) # (!\Mux25~7_combout  & (\Reg[23][6]~q  & ((ifid_ifinstr_o_23))))

	.dataa(\Reg[23][6]~q ),
	.datab(\Mux25~7_combout ),
	.datac(\Reg[31][6]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux25~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~8 .lut_mask = 16'hE2CC;
defparam \Mux25~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N5
dffeas \Reg[14][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][6] .is_wysiwyg = "true";
defparam \Reg[14][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N31
dffeas \Reg[15][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][6] .is_wysiwyg = "true";
defparam \Reg[15][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y37_N9
dffeas \Reg[13][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][6] .is_wysiwyg = "true";
defparam \Reg[13][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y37_N31
dffeas \Reg[12][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][6] .is_wysiwyg = "true";
defparam \Reg[12][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y37_N30
cycloneive_lcell_comb \Mux25~17 (
// Equation(s):
// \Mux25~17_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[13][6]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[12][6]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[13][6]~q ),
	.datac(\Reg[12][6]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux25~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~17 .lut_mask = 16'hEE50;
defparam \Mux25~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N30
cycloneive_lcell_comb \Mux25~18 (
// Equation(s):
// \Mux25~18_combout  = (ifid_ifinstr_o_22 & ((\Mux25~17_combout  & ((\Reg[15][6]~q ))) # (!\Mux25~17_combout  & (\Reg[14][6]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux25~17_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[14][6]~q ),
	.datac(\Reg[15][6]~q ),
	.datad(\Mux25~17_combout ),
	.cin(gnd),
	.combout(\Mux25~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~18 .lut_mask = 16'hF588;
defparam \Mux25~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N9
dffeas \Reg[5][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][6] .is_wysiwyg = "true";
defparam \Reg[5][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N19
dffeas \Reg[4][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][6] .is_wysiwyg = "true";
defparam \Reg[4][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N8
cycloneive_lcell_comb \Mux25~10 (
// Equation(s):
// \Mux25~10_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[5][6]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[4][6]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[5][6]~q ),
	.datad(\Reg[4][6]~q ),
	.cin(gnd),
	.combout(\Mux25~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~10 .lut_mask = 16'hD9C8;
defparam \Mux25~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N13
dffeas \Reg[6][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][6] .is_wysiwyg = "true";
defparam \Reg[6][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y39_N11
dffeas \Reg[7][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][6] .is_wysiwyg = "true";
defparam \Reg[7][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N12
cycloneive_lcell_comb \Mux25~11 (
// Equation(s):
// \Mux25~11_combout  = (\Mux25~10_combout  & (((\Reg[7][6]~q )) # (!ifid_ifinstr_o_22))) # (!\Mux25~10_combout  & (ifid_ifinstr_o_22 & (\Reg[6][6]~q )))

	.dataa(\Mux25~10_combout ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[6][6]~q ),
	.datad(\Reg[7][6]~q ),
	.cin(gnd),
	.combout(\Mux25~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~11 .lut_mask = 16'hEA62;
defparam \Mux25~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N11
dffeas \Reg[2][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][6] .is_wysiwyg = "true";
defparam \Reg[2][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N10
cycloneive_lcell_comb \Mux25~15 (
// Equation(s):
// \Mux25~15_combout  = (\Mux25~14_combout ) # ((!ifid_ifinstr_o_21 & (\Reg[2][6]~q  & ifid_ifinstr_o_22)))

	.dataa(\Mux25~14_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[2][6]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux25~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~15 .lut_mask = 16'hBAAA;
defparam \Mux25~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N17
dffeas \Reg[9][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][6] .is_wysiwyg = "true";
defparam \Reg[9][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N11
dffeas \Reg[11][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][6] .is_wysiwyg = "true";
defparam \Reg[11][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N19
dffeas \Reg[8][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][6] .is_wysiwyg = "true";
defparam \Reg[8][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N21
dffeas \Reg[10][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][6] .is_wysiwyg = "true";
defparam \Reg[10][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N18
cycloneive_lcell_comb \Mux25~12 (
// Equation(s):
// \Mux25~12_combout  = (ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21) # ((\Reg[10][6]~q )))) # (!ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & (\Reg[8][6]~q )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[8][6]~q ),
	.datad(\Reg[10][6]~q ),
	.cin(gnd),
	.combout(\Mux25~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~12 .lut_mask = 16'hBA98;
defparam \Mux25~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N10
cycloneive_lcell_comb \Mux25~13 (
// Equation(s):
// \Mux25~13_combout  = (ifid_ifinstr_o_21 & ((\Mux25~12_combout  & ((\Reg[11][6]~q ))) # (!\Mux25~12_combout  & (\Reg[9][6]~q )))) # (!ifid_ifinstr_o_21 & (((\Mux25~12_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[9][6]~q ),
	.datac(\Reg[11][6]~q ),
	.datad(\Mux25~12_combout ),
	.cin(gnd),
	.combout(\Mux25~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~13 .lut_mask = 16'hF588;
defparam \Mux25~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N10
cycloneive_lcell_comb \Mux25~16 (
// Equation(s):
// \Mux25~16_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Mux25~13_combout ))) # (!ifid_ifinstr_o_24 & (\Mux25~15_combout ))))

	.dataa(\Mux25~15_combout ),
	.datab(ifid_ifinstr_o_23),
	.datac(ifid_ifinstr_o_24),
	.datad(\Mux25~13_combout ),
	.cin(gnd),
	.combout(\Mux25~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~16 .lut_mask = 16'hF2C2;
defparam \Mux25~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N20
cycloneive_lcell_comb \Reg[27][5]~feeder (
// Equation(s):
// \Reg[27][5]~feeder_combout  = \wdat~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat8),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[27][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[27][5]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[27][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N21
dffeas \Reg[27][5] (
	.clk(!CLK),
	.d(\Reg[27][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][5] .is_wysiwyg = "true";
defparam \Reg[27][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y29_N11
dffeas \Reg[31][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][5] .is_wysiwyg = "true";
defparam \Reg[31][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N7
dffeas \Reg[23][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][5] .is_wysiwyg = "true";
defparam \Reg[23][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N6
cycloneive_lcell_comb \Mux26~7 (
// Equation(s):
// \Mux26~7_combout  = (ifid_ifinstr_o_23 & (((\Reg[23][5]~q ) # (ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (\Reg[19][5]~q  & ((!ifid_ifinstr_o_24))))

	.dataa(\Reg[19][5]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[23][5]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux26~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~7 .lut_mask = 16'hCCE2;
defparam \Mux26~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N10
cycloneive_lcell_comb \Mux26~8 (
// Equation(s):
// \Mux26~8_combout  = (ifid_ifinstr_o_24 & ((\Mux26~7_combout  & ((\Reg[31][5]~q ))) # (!\Mux26~7_combout  & (\Reg[27][5]~q )))) # (!ifid_ifinstr_o_24 & (((\Mux26~7_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[27][5]~q ),
	.datac(\Reg[31][5]~q ),
	.datad(\Mux26~7_combout ),
	.cin(gnd),
	.combout(\Mux26~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~8 .lut_mask = 16'hF588;
defparam \Mux26~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N28
cycloneive_lcell_comb \Reg[21][5]~feeder (
// Equation(s):
// \Reg[21][5]~feeder_combout  = \wdat~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat8),
	.cin(gnd),
	.combout(\Reg[21][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[21][5]~feeder .lut_mask = 16'hFF00;
defparam \Reg[21][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N29
dffeas \Reg[21][5] (
	.clk(!CLK),
	.d(\Reg[21][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][5] .is_wysiwyg = "true";
defparam \Reg[21][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N5
dffeas \Reg[17][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][5] .is_wysiwyg = "true";
defparam \Reg[17][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N4
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (ifid_ifinstr_o_23 & ((\Reg[21][5]~q ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((\Reg[17][5]~q  & !ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[21][5]~q ),
	.datac(\Reg[17][5]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hAAD8;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N31
dffeas \Reg[29][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][5] .is_wysiwyg = "true";
defparam \Reg[29][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y38_N27
dffeas \Reg[25][5] (
	.clk(!CLK),
	.d(wdat8),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][5] .is_wysiwyg = "true";
defparam \Reg[25][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N30
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// \Mux26~1_combout  = (ifid_ifinstr_o_24 & ((\Mux26~0_combout  & (\Reg[29][5]~q )) # (!\Mux26~0_combout  & ((\Reg[25][5]~q ))))) # (!ifid_ifinstr_o_24 & (\Mux26~0_combout ))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux26~0_combout ),
	.datac(\Reg[29][5]~q ),
	.datad(\Reg[25][5]~q ),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hE6C4;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y33_N13
dffeas \Reg[16][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][5] .is_wysiwyg = "true";
defparam \Reg[16][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y33_N13
dffeas \Reg[24][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][5] .is_wysiwyg = "true";
defparam \Reg[24][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N12
cycloneive_lcell_comb \Mux26~4 (
// Equation(s):
// \Mux26~4_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Reg[24][5]~q ))) # (!ifid_ifinstr_o_24 & (\Reg[16][5]~q ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[16][5]~q ),
	.datad(\Reg[24][5]~q ),
	.cin(gnd),
	.combout(\Mux26~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~4 .lut_mask = 16'hDC98;
defparam \Mux26~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N31
dffeas \Reg[28][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][5] .is_wysiwyg = "true";
defparam \Reg[28][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y33_N19
dffeas \Reg[20][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][5] .is_wysiwyg = "true";
defparam \Reg[20][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N30
cycloneive_lcell_comb \Mux26~5 (
// Equation(s):
// \Mux26~5_combout  = (ifid_ifinstr_o_23 & ((\Mux26~4_combout  & (\Reg[28][5]~q )) # (!\Mux26~4_combout  & ((\Reg[20][5]~q ))))) # (!ifid_ifinstr_o_23 & (\Mux26~4_combout ))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux26~4_combout ),
	.datac(\Reg[28][5]~q ),
	.datad(\Reg[20][5]~q ),
	.cin(gnd),
	.combout(\Mux26~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~5 .lut_mask = 16'hE6C4;
defparam \Mux26~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N15
dffeas \Reg[18][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][5] .is_wysiwyg = "true";
defparam \Reg[18][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N6
cycloneive_lcell_comb \Reg[26][5]~feeder (
// Equation(s):
// \Reg[26][5]~feeder_combout  = \wdat~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat8),
	.cin(gnd),
	.combout(\Reg[26][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[26][5]~feeder .lut_mask = 16'hFF00;
defparam \Reg[26][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N7
dffeas \Reg[26][5] (
	.clk(!CLK),
	.d(\Reg[26][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][5] .is_wysiwyg = "true";
defparam \Reg[26][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N14
cycloneive_lcell_comb \Mux26~2 (
// Equation(s):
// \Mux26~2_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[26][5]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & (\Reg[18][5]~q )))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[18][5]~q ),
	.datad(\Reg[26][5]~q ),
	.cin(gnd),
	.combout(\Mux26~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~2 .lut_mask = 16'hBA98;
defparam \Mux26~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N5
dffeas \Reg[22][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][5] .is_wysiwyg = "true";
defparam \Reg[22][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N28
cycloneive_lcell_comb \Reg[30][5]~feeder (
// Equation(s):
// \Reg[30][5]~feeder_combout  = \wdat~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat8),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[30][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[30][5]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[30][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N29
dffeas \Reg[30][5] (
	.clk(!CLK),
	.d(\Reg[30][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][5] .is_wysiwyg = "true";
defparam \Reg[30][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N4
cycloneive_lcell_comb \Mux26~3 (
// Equation(s):
// \Mux26~3_combout  = (ifid_ifinstr_o_23 & ((\Mux26~2_combout  & ((\Reg[30][5]~q ))) # (!\Mux26~2_combout  & (\Reg[22][5]~q )))) # (!ifid_ifinstr_o_23 & (\Mux26~2_combout ))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux26~2_combout ),
	.datac(\Reg[22][5]~q ),
	.datad(\Reg[30][5]~q ),
	.cin(gnd),
	.combout(\Mux26~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~3 .lut_mask = 16'hEC64;
defparam \Mux26~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N22
cycloneive_lcell_comb \Mux26~6 (
// Equation(s):
// \Mux26~6_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Mux26~3_combout ))) # (!ifid_ifinstr_o_22 & (\Mux26~5_combout ))))

	.dataa(\Mux26~5_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(ifid_ifinstr_o_22),
	.datad(\Mux26~3_combout ),
	.cin(gnd),
	.combout(\Mux26~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~6 .lut_mask = 16'hF2C2;
defparam \Mux26~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N7
dffeas \Reg[7][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][5] .is_wysiwyg = "true";
defparam \Reg[7][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N3
dffeas \Reg[4][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][5] .is_wysiwyg = "true";
defparam \Reg[4][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N21
dffeas \Reg[5][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][5] .is_wysiwyg = "true";
defparam \Reg[5][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N2
cycloneive_lcell_comb \Mux26~12 (
// Equation(s):
// \Mux26~12_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[5][5]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[4][5]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[4][5]~q ),
	.datad(\Reg[5][5]~q ),
	.cin(gnd),
	.combout(\Mux26~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~12 .lut_mask = 16'hDC98;
defparam \Mux26~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N6
cycloneive_lcell_comb \Mux26~13 (
// Equation(s):
// \Mux26~13_combout  = (ifid_ifinstr_o_22 & ((\Mux26~12_combout  & ((\Reg[7][5]~q ))) # (!\Mux26~12_combout  & (\Reg[6][5]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux26~12_combout ))))

	.dataa(\Reg[6][5]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[7][5]~q ),
	.datad(\Mux26~12_combout ),
	.cin(gnd),
	.combout(\Mux26~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~13 .lut_mask = 16'hF388;
defparam \Mux26~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y31_N15
dffeas \Reg[2][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][5] .is_wysiwyg = "true";
defparam \Reg[2][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y35_N23
dffeas \Reg[1][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][5] .is_wysiwyg = "true";
defparam \Reg[1][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N12
cycloneive_lcell_comb \Reg[3][5]~feeder (
// Equation(s):
// \Reg[3][5]~feeder_combout  = \wdat~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat8),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[3][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[3][5]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[3][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y35_N13
dffeas \Reg[3][5] (
	.clk(!CLK),
	.d(\Reg[3][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][5] .is_wysiwyg = "true";
defparam \Reg[3][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N22
cycloneive_lcell_comb \Mux26~14 (
// Equation(s):
// \Mux26~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][5]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][5]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[1][5]~q ),
	.datad(\Reg[3][5]~q ),
	.cin(gnd),
	.combout(\Mux26~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~14 .lut_mask = 16'hA820;
defparam \Mux26~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N12
cycloneive_lcell_comb \Mux26~15 (
// Equation(s):
// \Mux26~15_combout  = (\Mux26~14_combout ) # ((ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & \Reg[2][5]~q )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[2][5]~q ),
	.datad(\Mux26~14_combout ),
	.cin(gnd),
	.combout(\Mux26~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~15 .lut_mask = 16'hFF20;
defparam \Mux26~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N20
cycloneive_lcell_comb \Mux26~16 (
// Equation(s):
// \Mux26~16_combout  = (ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24) # ((\Mux26~13_combout )))) # (!ifid_ifinstr_o_23 & (!ifid_ifinstr_o_24 & ((\Mux26~15_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Mux26~13_combout ),
	.datad(\Mux26~15_combout ),
	.cin(gnd),
	.combout(\Mux26~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~16 .lut_mask = 16'hB9A8;
defparam \Mux26~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y31_N29
dffeas \Reg[10][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][5] .is_wysiwyg = "true";
defparam \Reg[10][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N28
cycloneive_lcell_comb \Mux26~10 (
// Equation(s):
// \Mux26~10_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[10][5]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[8][5]~q ))))

	.dataa(\Reg[8][5]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[10][5]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux26~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~10 .lut_mask = 16'hFC22;
defparam \Mux26~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N27
dffeas \Reg[11][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][5] .is_wysiwyg = "true";
defparam \Reg[11][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N12
cycloneive_lcell_comb \Reg[9][5]~feeder (
// Equation(s):
// \Reg[9][5]~feeder_combout  = \wdat~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat8),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[9][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[9][5]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[9][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N13
dffeas \Reg[9][5] (
	.clk(!CLK),
	.d(\Reg[9][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][5] .is_wysiwyg = "true";
defparam \Reg[9][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N24
cycloneive_lcell_comb \Mux26~11 (
// Equation(s):
// \Mux26~11_combout  = (ifid_ifinstr_o_21 & ((\Mux26~10_combout  & (\Reg[11][5]~q )) # (!\Mux26~10_combout  & ((\Reg[9][5]~q ))))) # (!ifid_ifinstr_o_21 & (\Mux26~10_combout ))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux26~10_combout ),
	.datac(\Reg[11][5]~q ),
	.datad(\Reg[9][5]~q ),
	.cin(gnd),
	.combout(\Mux26~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~11 .lut_mask = 16'hE6C4;
defparam \Mux26~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N27
dffeas \Reg[15][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][5] .is_wysiwyg = "true";
defparam \Reg[15][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N25
dffeas \Reg[14][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][5] .is_wysiwyg = "true";
defparam \Reg[14][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N28
cycloneive_lcell_comb \Reg[13][5]~feeder (
// Equation(s):
// \Reg[13][5]~feeder_combout  = \wdat~17_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat8),
	.cin(gnd),
	.combout(\Reg[13][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[13][5]~feeder .lut_mask = 16'hFF00;
defparam \Reg[13][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N29
dffeas \Reg[13][5] (
	.clk(!CLK),
	.d(\Reg[13][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][5] .is_wysiwyg = "true";
defparam \Reg[13][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N30
cycloneive_lcell_comb \Mux26~17 (
// Equation(s):
// \Mux26~17_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[13][5]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[12][5]~q ))))

	.dataa(\Reg[12][5]~q ),
	.datab(\Reg[13][5]~q ),
	.datac(ifid_ifinstr_o_22),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux26~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~17 .lut_mask = 16'hFC0A;
defparam \Mux26~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N24
cycloneive_lcell_comb \Mux26~18 (
// Equation(s):
// \Mux26~18_combout  = (ifid_ifinstr_o_22 & ((\Mux26~17_combout  & (\Reg[15][5]~q )) # (!\Mux26~17_combout  & ((\Reg[14][5]~q ))))) # (!ifid_ifinstr_o_22 & (((\Mux26~17_combout ))))

	.dataa(\Reg[15][5]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[14][5]~q ),
	.datad(\Mux26~17_combout ),
	.cin(gnd),
	.combout(\Mux26~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~18 .lut_mask = 16'hBBC0;
defparam \Mux26~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N14
cycloneive_lcell_comb \Mux60~7 (
// Equation(s):
// \Mux60~7_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[27][3]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[19][3]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[19][3]~q ),
	.datad(\Reg[27][3]~q ),
	.cin(gnd),
	.combout(\Mux60~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~7 .lut_mask = 16'hDC98;
defparam \Mux60~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N8
cycloneive_lcell_comb \Mux60~8 (
// Equation(s):
// \Mux60~8_combout  = (\Mux60~7_combout  & (((\Reg[31][3]~q ) # (!ifid_ifinstr_o_18)))) # (!\Mux60~7_combout  & (\Reg[23][3]~q  & ((ifid_ifinstr_o_18))))

	.dataa(\Mux60~7_combout ),
	.datab(\Reg[23][3]~q ),
	.datac(\Reg[31][3]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux60~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~8 .lut_mask = 16'hE4AA;
defparam \Mux60~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N26
cycloneive_lcell_comb \Mux60~0 (
// Equation(s):
// \Mux60~0_combout  = (ifid_ifinstr_o_19 & ((\Reg[25][3]~q ) # ((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & (((\Reg[17][3]~q  & !ifid_ifinstr_o_18))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[25][3]~q ),
	.datac(\Reg[17][3]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux60~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~0 .lut_mask = 16'hAAD8;
defparam \Mux60~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N4
cycloneive_lcell_comb \Mux60~1 (
// Equation(s):
// \Mux60~1_combout  = (\Mux60~0_combout  & (((\Reg[29][3]~q ) # (!ifid_ifinstr_o_18)))) # (!\Mux60~0_combout  & (\Reg[21][3]~q  & ((ifid_ifinstr_o_18))))

	.dataa(\Mux60~0_combout ),
	.datab(\Reg[21][3]~q ),
	.datac(\Reg[29][3]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux60~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~1 .lut_mask = 16'hE4AA;
defparam \Mux60~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N20
cycloneive_lcell_comb \Mux60~3 (
// Equation(s):
// \Mux60~3_combout  = (\Mux60~2_combout  & ((\Reg[30][3]~q ) # ((!ifid_ifinstr_o_19)))) # (!\Mux60~2_combout  & (((ifid_ifinstr_o_19 & \Reg[26][3]~q ))))

	.dataa(\Mux60~2_combout ),
	.datab(\Reg[30][3]~q ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Reg[26][3]~q ),
	.cin(gnd),
	.combout(\Mux60~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~3 .lut_mask = 16'hDA8A;
defparam \Mux60~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N22
cycloneive_lcell_comb \Mux60~4 (
// Equation(s):
// \Mux60~4_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[20][3]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[16][3]~q )))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[20][3]~q ),
	.datad(\Reg[16][3]~q ),
	.cin(gnd),
	.combout(\Mux60~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~4 .lut_mask = 16'hD9C8;
defparam \Mux60~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N14
cycloneive_lcell_comb \Mux60~5 (
// Equation(s):
// \Mux60~5_combout  = (ifid_ifinstr_o_19 & ((\Mux60~4_combout  & ((\Reg[28][3]~q ))) # (!\Mux60~4_combout  & (\Reg[24][3]~q )))) # (!ifid_ifinstr_o_19 & (((\Mux60~4_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[24][3]~q ),
	.datac(\Reg[28][3]~q ),
	.datad(\Mux60~4_combout ),
	.cin(gnd),
	.combout(\Mux60~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~5 .lut_mask = 16'hF588;
defparam \Mux60~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N30
cycloneive_lcell_comb \Mux60~6 (
// Equation(s):
// \Mux60~6_combout  = (ifid_ifinstr_o_17 & ((\Mux60~3_combout ) # ((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & (((\Mux60~5_combout  & !ifid_ifinstr_o_16))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux60~3_combout ),
	.datac(\Mux60~5_combout ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux60~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~6 .lut_mask = 16'hAAD8;
defparam \Mux60~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N6
cycloneive_lcell_comb \Reg[6][3]~feeder (
// Equation(s):
// \Reg[6][3]~feeder_combout  = \wdat~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat4),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[6][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[6][3]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[6][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N7
dffeas \Reg[6][3] (
	.clk(!CLK),
	.d(\Reg[6][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][3] .is_wysiwyg = "true";
defparam \Reg[6][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N8
cycloneive_lcell_comb \Mux60~10 (
// Equation(s):
// \Mux60~10_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[5][3]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[4][3]~q ))))

	.dataa(\Reg[4][3]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[5][3]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux60~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~10 .lut_mask = 16'hFC22;
defparam \Mux60~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N24
cycloneive_lcell_comb \Mux60~11 (
// Equation(s):
// \Mux60~11_combout  = (ifid_ifinstr_o_17 & ((\Mux60~10_combout  & ((\Reg[7][3]~q ))) # (!\Mux60~10_combout  & (\Reg[6][3]~q )))) # (!ifid_ifinstr_o_17 & (((\Mux60~10_combout ))))

	.dataa(\Reg[6][3]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[7][3]~q ),
	.datad(\Mux60~10_combout ),
	.cin(gnd),
	.combout(\Mux60~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~11 .lut_mask = 16'hF388;
defparam \Mux60~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N20
cycloneive_lcell_comb \Mux60~17 (
// Equation(s):
// \Mux60~17_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[13][3]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[12][3]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[12][3]~q ),
	.datac(\Reg[13][3]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux60~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~17 .lut_mask = 16'hFA44;
defparam \Mux60~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N16
cycloneive_lcell_comb \Mux60~18 (
// Equation(s):
// \Mux60~18_combout  = (ifid_ifinstr_o_17 & ((\Mux60~17_combout  & ((\Reg[15][3]~q ))) # (!\Mux60~17_combout  & (\Reg[14][3]~q )))) # (!ifid_ifinstr_o_17 & (\Mux60~17_combout ))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux60~17_combout ),
	.datac(\Reg[14][3]~q ),
	.datad(\Reg[15][3]~q ),
	.cin(gnd),
	.combout(\Mux60~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~18 .lut_mask = 16'hEC64;
defparam \Mux60~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N23
dffeas \Reg[8][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][3] .is_wysiwyg = "true";
defparam \Reg[8][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N22
cycloneive_lcell_comb \Mux60~12 (
// Equation(s):
// \Mux60~12_combout  = (ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16) # ((\Reg[10][3]~q )))) # (!ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & (\Reg[8][3]~q )))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[8][3]~q ),
	.datad(\Reg[10][3]~q ),
	.cin(gnd),
	.combout(\Mux60~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~12 .lut_mask = 16'hBA98;
defparam \Mux60~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N18
cycloneive_lcell_comb \Mux60~13 (
// Equation(s):
// \Mux60~13_combout  = (ifid_ifinstr_o_16 & ((\Mux60~12_combout  & ((\Reg[11][3]~q ))) # (!\Mux60~12_combout  & (\Reg[9][3]~q )))) # (!ifid_ifinstr_o_16 & (((\Mux60~12_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[9][3]~q ),
	.datac(\Reg[11][3]~q ),
	.datad(\Mux60~12_combout ),
	.cin(gnd),
	.combout(\Mux60~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~13 .lut_mask = 16'hF588;
defparam \Mux60~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N29
dffeas \Reg[3][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat4),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][3] .is_wysiwyg = "true";
defparam \Reg[3][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N28
cycloneive_lcell_comb \Mux60~14 (
// Equation(s):
// \Mux60~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[3][3]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[1][3]~q ))))

	.dataa(\Reg[1][3]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[3][3]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux60~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~14 .lut_mask = 16'hE200;
defparam \Mux60~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N0
cycloneive_lcell_comb \Mux60~15 (
// Equation(s):
// \Mux60~15_combout  = (\Mux60~14_combout ) # ((ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & \Reg[2][3]~q )))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux60~14_combout ),
	.datad(\Reg[2][3]~q ),
	.cin(gnd),
	.combout(\Mux60~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~15 .lut_mask = 16'hF2F0;
defparam \Mux60~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N18
cycloneive_lcell_comb \Mux60~16 (
// Equation(s):
// \Mux60~16_combout  = (ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18) # ((\Mux60~13_combout )))) # (!ifid_ifinstr_o_19 & (!ifid_ifinstr_o_18 & ((\Mux60~15_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Mux60~13_combout ),
	.datad(\Mux60~15_combout ),
	.cin(gnd),
	.combout(\Mux60~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~16 .lut_mask = 16'hB9A8;
defparam \Mux60~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N15
dffeas \Reg[31][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][16] .is_wysiwyg = "true";
defparam \Reg[31][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N13
dffeas \Reg[27][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][16] .is_wysiwyg = "true";
defparam \Reg[27][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N31
dffeas \Reg[19][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][16] .is_wysiwyg = "true";
defparam \Reg[19][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N12
cycloneive_lcell_comb \Mux15~7 (
// Equation(s):
// \Mux15~7_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[27][16]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[19][16]~q )))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[27][16]~q ),
	.datad(\Reg[19][16]~q ),
	.cin(gnd),
	.combout(\Mux15~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~7 .lut_mask = 16'hD9C8;
defparam \Mux15~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N17
dffeas \Reg[23][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][16] .is_wysiwyg = "true";
defparam \Reg[23][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N16
cycloneive_lcell_comb \Mux15~8 (
// Equation(s):
// \Mux15~8_combout  = (\Mux15~7_combout  & ((\Reg[31][16]~q ) # ((!ifid_ifinstr_o_23)))) # (!\Mux15~7_combout  & (((\Reg[23][16]~q  & ifid_ifinstr_o_23))))

	.dataa(\Reg[31][16]~q ),
	.datab(\Mux15~7_combout ),
	.datac(\Reg[23][16]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux15~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~8 .lut_mask = 16'hB8CC;
defparam \Mux15~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N15
dffeas \Reg[17][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][16] .is_wysiwyg = "true";
defparam \Reg[17][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N16
cycloneive_lcell_comb \Reg[25][16]~feeder (
// Equation(s):
// \Reg[25][16]~feeder_combout  = \wdat~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat9),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[25][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][16]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[25][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N17
dffeas \Reg[25][16] (
	.clk(!CLK),
	.d(\Reg[25][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][16] .is_wysiwyg = "true";
defparam \Reg[25][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N14
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// \Mux15~0_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Reg[25][16]~q ))) # (!ifid_ifinstr_o_24 & (\Reg[17][16]~q ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[17][16]~q ),
	.datad(\Reg[25][16]~q ),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hDC98;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N24
cycloneive_lcell_comb \Reg[29][16]~feeder (
// Equation(s):
// \Reg[29][16]~feeder_combout  = \wdat~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat9),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[29][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[29][16]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[29][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y38_N25
dffeas \Reg[29][16] (
	.clk(!CLK),
	.d(\Reg[29][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][16] .is_wysiwyg = "true";
defparam \Reg[29][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y37_N27
dffeas \Reg[21][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][16] .is_wysiwyg = "true";
defparam \Reg[21][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N12
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// \Mux15~1_combout  = (\Mux15~0_combout  & ((\Reg[29][16]~q ) # ((!ifid_ifinstr_o_23)))) # (!\Mux15~0_combout  & (((\Reg[21][16]~q  & ifid_ifinstr_o_23))))

	.dataa(\Mux15~0_combout ),
	.datab(\Reg[29][16]~q ),
	.datac(\Reg[21][16]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'hD8AA;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y32_N5
dffeas \Reg[24][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][16] .is_wysiwyg = "true";
defparam \Reg[24][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y32_N23
dffeas \Reg[16][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][16] .is_wysiwyg = "true";
defparam \Reg[16][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N22
cycloneive_lcell_comb \Mux15~4 (
// Equation(s):
// \Mux15~4_combout  = (ifid_ifinstr_o_23 & ((\Reg[20][16]~q ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((\Reg[16][16]~q  & !ifid_ifinstr_o_24))))

	.dataa(\Reg[20][16]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[16][16]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux15~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~4 .lut_mask = 16'hCCB8;
defparam \Mux15~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N28
cycloneive_lcell_comb \Mux15~5 (
// Equation(s):
// \Mux15~5_combout  = (ifid_ifinstr_o_24 & ((\Mux15~4_combout  & (\Reg[28][16]~q )) # (!\Mux15~4_combout  & ((\Reg[24][16]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux15~4_combout ))))

	.dataa(\Reg[28][16]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[24][16]~q ),
	.datad(\Mux15~4_combout ),
	.cin(gnd),
	.combout(\Mux15~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~5 .lut_mask = 16'hBBC0;
defparam \Mux15~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N25
dffeas \Reg[30][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][16] .is_wysiwyg = "true";
defparam \Reg[30][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N21
dffeas \Reg[26][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][16] .is_wysiwyg = "true";
defparam \Reg[26][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N20
cycloneive_lcell_comb \Mux15~3 (
// Equation(s):
// \Mux15~3_combout  = (\Mux15~2_combout  & ((\Reg[30][16]~q ) # ((!ifid_ifinstr_o_24)))) # (!\Mux15~2_combout  & (((\Reg[26][16]~q  & ifid_ifinstr_o_24))))

	.dataa(\Mux15~2_combout ),
	.datab(\Reg[30][16]~q ),
	.datac(\Reg[26][16]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux15~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~3 .lut_mask = 16'hD8AA;
defparam \Mux15~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N10
cycloneive_lcell_comb \Mux15~6 (
// Equation(s):
// \Mux15~6_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Mux15~3_combout ))) # (!ifid_ifinstr_o_22 & (\Mux15~5_combout ))))

	.dataa(\Mux15~5_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux15~3_combout ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux15~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~6 .lut_mask = 16'hFC22;
defparam \Mux15~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N23
dffeas \Reg[15][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][16] .is_wysiwyg = "true";
defparam \Reg[15][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N29
dffeas \Reg[14][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][16] .is_wysiwyg = "true";
defparam \Reg[14][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N3
dffeas \Reg[13][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][16] .is_wysiwyg = "true";
defparam \Reg[13][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N29
dffeas \Reg[12][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][16] .is_wysiwyg = "true";
defparam \Reg[12][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N28
cycloneive_lcell_comb \Mux15~17 (
// Equation(s):
// \Mux15~17_combout  = (ifid_ifinstr_o_21 & ((\Reg[13][16]~q ) # ((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & (((\Reg[12][16]~q  & !ifid_ifinstr_o_22))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[13][16]~q ),
	.datac(\Reg[12][16]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux15~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~17 .lut_mask = 16'hAAD8;
defparam \Mux15~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N28
cycloneive_lcell_comb \Mux15~18 (
// Equation(s):
// \Mux15~18_combout  = (ifid_ifinstr_o_22 & ((\Mux15~17_combout  & (\Reg[15][16]~q )) # (!\Mux15~17_combout  & ((\Reg[14][16]~q ))))) # (!ifid_ifinstr_o_22 & (((\Mux15~17_combout ))))

	.dataa(\Reg[15][16]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[14][16]~q ),
	.datad(\Mux15~17_combout ),
	.cin(gnd),
	.combout(\Mux15~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~18 .lut_mask = 16'hBBC0;
defparam \Mux15~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N23
dffeas \Reg[7][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][16] .is_wysiwyg = "true";
defparam \Reg[7][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y39_N25
dffeas \Reg[6][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][16] .is_wysiwyg = "true";
defparam \Reg[6][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N17
dffeas \Reg[5][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][16] .is_wysiwyg = "true";
defparam \Reg[5][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N11
dffeas \Reg[4][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][16] .is_wysiwyg = "true";
defparam \Reg[4][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N16
cycloneive_lcell_comb \Mux15~10 (
// Equation(s):
// \Mux15~10_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22) # ((\Reg[5][16]~q )))) # (!ifid_ifinstr_o_21 & (!ifid_ifinstr_o_22 & ((\Reg[4][16]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[5][16]~q ),
	.datad(\Reg[4][16]~q ),
	.cin(gnd),
	.combout(\Mux15~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~10 .lut_mask = 16'hB9A8;
defparam \Mux15~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N24
cycloneive_lcell_comb \Mux15~11 (
// Equation(s):
// \Mux15~11_combout  = (ifid_ifinstr_o_22 & ((\Mux15~10_combout  & (\Reg[7][16]~q )) # (!\Mux15~10_combout  & ((\Reg[6][16]~q ))))) # (!ifid_ifinstr_o_22 & (((\Mux15~10_combout ))))

	.dataa(\Reg[7][16]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[6][16]~q ),
	.datad(\Mux15~10_combout ),
	.cin(gnd),
	.combout(\Mux15~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~11 .lut_mask = 16'hBBC0;
defparam \Mux15~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N19
dffeas \Reg[1][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][16] .is_wysiwyg = "true";
defparam \Reg[1][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N21
dffeas \Reg[3][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][16] .is_wysiwyg = "true";
defparam \Reg[3][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N18
cycloneive_lcell_comb \Mux15~14 (
// Equation(s):
// \Mux15~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][16]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][16]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[1][16]~q ),
	.datad(\Reg[3][16]~q ),
	.cin(gnd),
	.combout(\Mux15~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~14 .lut_mask = 16'hA820;
defparam \Mux15~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N12
cycloneive_lcell_comb \Reg[2][16]~feeder (
// Equation(s):
// \Reg[2][16]~feeder_combout  = \wdat~21_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat9),
	.cin(gnd),
	.combout(\Reg[2][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[2][16]~feeder .lut_mask = 16'hFF00;
defparam \Reg[2][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y36_N13
dffeas \Reg[2][16] (
	.clk(!CLK),
	.d(\Reg[2][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][16] .is_wysiwyg = "true";
defparam \Reg[2][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N26
cycloneive_lcell_comb \Mux15~15 (
// Equation(s):
// \Mux15~15_combout  = (\Mux15~14_combout ) # ((!ifid_ifinstr_o_21 & (ifid_ifinstr_o_22 & \Reg[2][16]~q )))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Mux15~14_combout ),
	.datad(\Reg[2][16]~q ),
	.cin(gnd),
	.combout(\Mux15~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~15 .lut_mask = 16'hF4F0;
defparam \Mux15~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N3
dffeas \Reg[9][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][16] .is_wysiwyg = "true";
defparam \Reg[9][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y35_N9
dffeas \Reg[11][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][16] .is_wysiwyg = "true";
defparam \Reg[11][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N11
dffeas \Reg[8][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][16] .is_wysiwyg = "true";
defparam \Reg[8][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N21
dffeas \Reg[10][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][16] .is_wysiwyg = "true";
defparam \Reg[10][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N10
cycloneive_lcell_comb \Mux15~12 (
// Equation(s):
// \Mux15~12_combout  = (ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21) # ((\Reg[10][16]~q )))) # (!ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & (\Reg[8][16]~q )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[8][16]~q ),
	.datad(\Reg[10][16]~q ),
	.cin(gnd),
	.combout(\Mux15~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~12 .lut_mask = 16'hBA98;
defparam \Mux15~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N8
cycloneive_lcell_comb \Mux15~13 (
// Equation(s):
// \Mux15~13_combout  = (ifid_ifinstr_o_21 & ((\Mux15~12_combout  & ((\Reg[11][16]~q ))) # (!\Mux15~12_combout  & (\Reg[9][16]~q )))) # (!ifid_ifinstr_o_21 & (((\Mux15~12_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[9][16]~q ),
	.datac(\Reg[11][16]~q ),
	.datad(\Mux15~12_combout ),
	.cin(gnd),
	.combout(\Mux15~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~13 .lut_mask = 16'hF588;
defparam \Mux15~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N24
cycloneive_lcell_comb \Mux15~16 (
// Equation(s):
// \Mux15~16_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Mux15~13_combout )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & (\Mux15~15_combout )))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Mux15~15_combout ),
	.datad(\Mux15~13_combout ),
	.cin(gnd),
	.combout(\Mux15~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~16 .lut_mask = 16'hBA98;
defparam \Mux15~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N12
cycloneive_lcell_comb \Reg[25][15]~feeder (
// Equation(s):
// \Reg[25][15]~feeder_combout  = \wdat~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat10),
	.cin(gnd),
	.combout(\Reg[25][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][15]~feeder .lut_mask = 16'hFF00;
defparam \Reg[25][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N13
dffeas \Reg[25][15] (
	.clk(!CLK),
	.d(\Reg[25][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][15] .is_wysiwyg = "true";
defparam \Reg[25][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y37_N27
dffeas \Reg[29][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][15] .is_wysiwyg = "true";
defparam \Reg[29][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y37_N25
dffeas \Reg[21][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][15] .is_wysiwyg = "true";
defparam \Reg[21][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N19
dffeas \Reg[17][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][15] .is_wysiwyg = "true";
defparam \Reg[17][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N18
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// \Mux16~0_combout  = (ifid_ifinstr_o_23 & ((\Reg[21][15]~q ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((\Reg[17][15]~q  & !ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[21][15]~q ),
	.datac(\Reg[17][15]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'hAAD8;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N26
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// \Mux16~1_combout  = (ifid_ifinstr_o_24 & ((\Mux16~0_combout  & ((\Reg[29][15]~q ))) # (!\Mux16~0_combout  & (\Reg[25][15]~q )))) # (!ifid_ifinstr_o_24 & (((\Mux16~0_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[25][15]~q ),
	.datac(\Reg[29][15]~q ),
	.datad(\Mux16~0_combout ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hF588;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N26
cycloneive_lcell_comb \Reg[31][15]~feeder (
// Equation(s):
// \Reg[31][15]~feeder_combout  = \wdat~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat10),
	.cin(gnd),
	.combout(\Reg[31][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[31][15]~feeder .lut_mask = 16'hFF00;
defparam \Reg[31][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N27
dffeas \Reg[31][15] (
	.clk(!CLK),
	.d(\Reg[31][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][15] .is_wysiwyg = "true";
defparam \Reg[31][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N29
dffeas \Reg[27][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][15] .is_wysiwyg = "true";
defparam \Reg[27][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N19
dffeas \Reg[23][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][15] .is_wysiwyg = "true";
defparam \Reg[23][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y36_N17
dffeas \Reg[19][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][15] .is_wysiwyg = "true";
defparam \Reg[19][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N16
cycloneive_lcell_comb \Mux16~7 (
// Equation(s):
// \Mux16~7_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & (\Reg[23][15]~q )) # (!ifid_ifinstr_o_23 & ((\Reg[19][15]~q )))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[23][15]~q ),
	.datac(\Reg[19][15]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux16~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~7 .lut_mask = 16'hEE50;
defparam \Mux16~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N30
cycloneive_lcell_comb \Mux16~8 (
// Equation(s):
// \Mux16~8_combout  = (ifid_ifinstr_o_24 & ((\Mux16~7_combout  & (\Reg[31][15]~q )) # (!\Mux16~7_combout  & ((\Reg[27][15]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux16~7_combout ))))

	.dataa(\Reg[31][15]~q ),
	.datab(\Reg[27][15]~q ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Mux16~7_combout ),
	.cin(gnd),
	.combout(\Mux16~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~8 .lut_mask = 16'hAFC0;
defparam \Mux16~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N29
dffeas \Reg[26][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][15] .is_wysiwyg = "true";
defparam \Reg[26][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N28
cycloneive_lcell_comb \Mux16~2 (
// Equation(s):
// \Mux16~2_combout  = (ifid_ifinstr_o_24 & (((\Reg[26][15]~q ) # (ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & (\Reg[18][15]~q  & ((!ifid_ifinstr_o_23))))

	.dataa(\Reg[18][15]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[26][15]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux16~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~2 .lut_mask = 16'hCCE2;
defparam \Mux16~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N27
dffeas \Reg[30][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][15] .is_wysiwyg = "true";
defparam \Reg[30][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N30
cycloneive_lcell_comb \Reg[22][15]~feeder (
// Equation(s):
// \Reg[22][15]~feeder_combout  = \wdat~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat10),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[22][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[22][15]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[22][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N31
dffeas \Reg[22][15] (
	.clk(!CLK),
	.d(\Reg[22][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][15] .is_wysiwyg = "true";
defparam \Reg[22][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N26
cycloneive_lcell_comb \Mux16~3 (
// Equation(s):
// \Mux16~3_combout  = (ifid_ifinstr_o_23 & ((\Mux16~2_combout  & (\Reg[30][15]~q )) # (!\Mux16~2_combout  & ((\Reg[22][15]~q ))))) # (!ifid_ifinstr_o_23 & (\Mux16~2_combout ))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux16~2_combout ),
	.datac(\Reg[30][15]~q ),
	.datad(\Reg[22][15]~q ),
	.cin(gnd),
	.combout(\Mux16~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~3 .lut_mask = 16'hE6C4;
defparam \Mux16~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y33_N23
dffeas \Reg[20][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][15] .is_wysiwyg = "true";
defparam \Reg[20][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y33_N19
dffeas \Reg[28][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][15] .is_wysiwyg = "true";
defparam \Reg[28][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y33_N9
dffeas \Reg[16][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][15] .is_wysiwyg = "true";
defparam \Reg[16][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y33_N21
dffeas \Reg[24][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][15] .is_wysiwyg = "true";
defparam \Reg[24][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N8
cycloneive_lcell_comb \Mux16~4 (
// Equation(s):
// \Mux16~4_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[24][15]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & (\Reg[16][15]~q )))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[16][15]~q ),
	.datad(\Reg[24][15]~q ),
	.cin(gnd),
	.combout(\Mux16~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~4 .lut_mask = 16'hBA98;
defparam \Mux16~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N18
cycloneive_lcell_comb \Mux16~5 (
// Equation(s):
// \Mux16~5_combout  = (ifid_ifinstr_o_23 & ((\Mux16~4_combout  & ((\Reg[28][15]~q ))) # (!\Mux16~4_combout  & (\Reg[20][15]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux16~4_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[20][15]~q ),
	.datac(\Reg[28][15]~q ),
	.datad(\Mux16~4_combout ),
	.cin(gnd),
	.combout(\Mux16~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~5 .lut_mask = 16'hF588;
defparam \Mux16~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N20
cycloneive_lcell_comb \Mux16~6 (
// Equation(s):
// \Mux16~6_combout  = (ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21) # ((\Mux16~3_combout )))) # (!ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & ((\Mux16~5_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux16~3_combout ),
	.datad(\Mux16~5_combout ),
	.cin(gnd),
	.combout(\Mux16~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~6 .lut_mask = 16'hB9A8;
defparam \Mux16~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y36_N17
dffeas \Reg[3][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][15] .is_wysiwyg = "true";
defparam \Reg[3][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N19
dffeas \Reg[1][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][15] .is_wysiwyg = "true";
defparam \Reg[1][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N16
cycloneive_lcell_comb \Mux16~14 (
// Equation(s):
// \Mux16~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[3][15]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[1][15]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[3][15]~q ),
	.datad(\Reg[1][15]~q ),
	.cin(gnd),
	.combout(\Mux16~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~14 .lut_mask = 16'hA280;
defparam \Mux16~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N4
cycloneive_lcell_comb \Reg[2][15]~feeder (
// Equation(s):
// \Reg[2][15]~feeder_combout  = \wdat~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat10),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[2][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[2][15]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[2][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N5
dffeas \Reg[2][15] (
	.clk(!CLK),
	.d(\Reg[2][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][15] .is_wysiwyg = "true";
defparam \Reg[2][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N26
cycloneive_lcell_comb \Mux16~15 (
// Equation(s):
// \Mux16~15_combout  = (\Mux16~14_combout ) # ((ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & \Reg[2][15]~q )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux16~14_combout ),
	.datad(\Reg[2][15]~q ),
	.cin(gnd),
	.combout(\Mux16~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~15 .lut_mask = 16'hF2F0;
defparam \Mux16~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N5
dffeas \Reg[6][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][15] .is_wysiwyg = "true";
defparam \Reg[6][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y39_N3
dffeas \Reg[7][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][15] .is_wysiwyg = "true";
defparam \Reg[7][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N2
cycloneive_lcell_comb \Mux16~13 (
// Equation(s):
// \Mux16~13_combout  = (\Mux16~12_combout  & (((\Reg[7][15]~q ) # (!ifid_ifinstr_o_22)))) # (!\Mux16~12_combout  & (\Reg[6][15]~q  & ((ifid_ifinstr_o_22))))

	.dataa(\Mux16~12_combout ),
	.datab(\Reg[6][15]~q ),
	.datac(\Reg[7][15]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux16~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~13 .lut_mask = 16'hE4AA;
defparam \Mux16~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N8
cycloneive_lcell_comb \Mux16~16 (
// Equation(s):
// \Mux16~16_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24) # (\Mux16~13_combout )))) # (!ifid_ifinstr_o_23 & (\Mux16~15_combout  & (!ifid_ifinstr_o_24)))

	.dataa(\Mux16~15_combout ),
	.datab(ifid_ifinstr_o_23),
	.datac(ifid_ifinstr_o_24),
	.datad(\Mux16~13_combout ),
	.cin(gnd),
	.combout(\Mux16~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~16 .lut_mask = 16'hCEC2;
defparam \Mux16~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N9
dffeas \Reg[12][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][15] .is_wysiwyg = "true";
defparam \Reg[12][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N11
dffeas \Reg[13][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][15] .is_wysiwyg = "true";
defparam \Reg[13][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N10
cycloneive_lcell_comb \Mux16~17 (
// Equation(s):
// \Mux16~17_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[13][15]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[12][15]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[12][15]~q ),
	.datac(\Reg[13][15]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux16~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~17 .lut_mask = 16'hFA44;
defparam \Mux16~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N21
dffeas \Reg[14][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][15] .is_wysiwyg = "true";
defparam \Reg[14][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N19
dffeas \Reg[15][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][15] .is_wysiwyg = "true";
defparam \Reg[15][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N20
cycloneive_lcell_comb \Mux16~18 (
// Equation(s):
// \Mux16~18_combout  = (\Mux16~17_combout  & (((\Reg[15][15]~q )) # (!ifid_ifinstr_o_22))) # (!\Mux16~17_combout  & (ifid_ifinstr_o_22 & (\Reg[14][15]~q )))

	.dataa(\Mux16~17_combout ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[14][15]~q ),
	.datad(\Reg[15][15]~q ),
	.cin(gnd),
	.combout(\Mux16~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~18 .lut_mask = 16'hEA62;
defparam \Mux16~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N31
dffeas \Reg[9][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][15] .is_wysiwyg = "true";
defparam \Reg[9][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N16
cycloneive_lcell_comb \Reg[11][15]~feeder (
// Equation(s):
// \Reg[11][15]~feeder_combout  = \wdat~23_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat10),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[11][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[11][15]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[11][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N17
dffeas \Reg[11][15] (
	.clk(!CLK),
	.d(\Reg[11][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][15] .is_wysiwyg = "true";
defparam \Reg[11][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N5
dffeas \Reg[10][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][15] .is_wysiwyg = "true";
defparam \Reg[10][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N4
cycloneive_lcell_comb \Mux16~10 (
// Equation(s):
// \Mux16~10_combout  = (ifid_ifinstr_o_22 & (((\Reg[10][15]~q ) # (ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & (\Reg[8][15]~q  & ((!ifid_ifinstr_o_21))))

	.dataa(\Reg[8][15]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[10][15]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux16~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~10 .lut_mask = 16'hCCE2;
defparam \Mux16~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N6
cycloneive_lcell_comb \Mux16~11 (
// Equation(s):
// \Mux16~11_combout  = (ifid_ifinstr_o_21 & ((\Mux16~10_combout  & ((\Reg[11][15]~q ))) # (!\Mux16~10_combout  & (\Reg[9][15]~q )))) # (!ifid_ifinstr_o_21 & (((\Mux16~10_combout ))))

	.dataa(\Reg[9][15]~q ),
	.datab(\Reg[11][15]~q ),
	.datac(ifid_ifinstr_o_21),
	.datad(\Mux16~10_combout ),
	.cin(gnd),
	.combout(\Mux16~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~11 .lut_mask = 16'hCFA0;
defparam \Mux16~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N18
cycloneive_lcell_comb \Reg[21][14]~feeder (
// Equation(s):
// \Reg[21][14]~feeder_combout  = \wdat~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat11),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[21][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[21][14]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[21][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N19
dffeas \Reg[21][14] (
	.clk(!CLK),
	.d(\Reg[21][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][14] .is_wysiwyg = "true";
defparam \Reg[21][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N13
dffeas \Reg[29][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][14] .is_wysiwyg = "true";
defparam \Reg[29][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N8
cycloneive_lcell_comb \Reg[17][14]~feeder (
// Equation(s):
// \Reg[17][14]~feeder_combout  = \wdat~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat11),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[17][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[17][14]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[17][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y37_N9
dffeas \Reg[17][14] (
	.clk(!CLK),
	.d(\Reg[17][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][14] .is_wysiwyg = "true";
defparam \Reg[17][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N2
cycloneive_lcell_comb \Reg[25][14]~feeder (
// Equation(s):
// \Reg[25][14]~feeder_combout  = \wdat~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat11),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[25][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][14]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[25][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N3
dffeas \Reg[25][14] (
	.clk(!CLK),
	.d(\Reg[25][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][14] .is_wysiwyg = "true";
defparam \Reg[25][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N22
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// \Mux17~0_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Reg[25][14]~q ))) # (!ifid_ifinstr_o_24 & (\Reg[17][14]~q ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[17][14]~q ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Reg[25][14]~q ),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'hF4A4;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N20
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// \Mux17~1_combout  = (ifid_ifinstr_o_23 & ((\Mux17~0_combout  & ((\Reg[29][14]~q ))) # (!\Mux17~0_combout  & (\Reg[21][14]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux17~0_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[21][14]~q ),
	.datac(\Reg[29][14]~q ),
	.datad(\Mux17~0_combout ),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hF588;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y34_N31
dffeas \Reg[28][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][14] .is_wysiwyg = "true";
defparam \Reg[28][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N28
cycloneive_lcell_comb \Reg[24][14]~feeder (
// Equation(s):
// \Reg[24][14]~feeder_combout  = \wdat~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat11),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[24][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[24][14]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[24][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N29
dffeas \Reg[24][14] (
	.clk(!CLK),
	.d(\Reg[24][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][14] .is_wysiwyg = "true";
defparam \Reg[24][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N30
cycloneive_lcell_comb \Mux17~5 (
// Equation(s):
// \Mux17~5_combout  = (\Mux17~4_combout  & (((\Reg[28][14]~q )) # (!ifid_ifinstr_o_24))) # (!\Mux17~4_combout  & (ifid_ifinstr_o_24 & ((\Reg[24][14]~q ))))

	.dataa(\Mux17~4_combout ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[28][14]~q ),
	.datad(\Reg[24][14]~q ),
	.cin(gnd),
	.combout(\Mux17~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~5 .lut_mask = 16'hE6A2;
defparam \Mux17~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N1
dffeas \Reg[26][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][14] .is_wysiwyg = "true";
defparam \Reg[26][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y33_N3
dffeas \Reg[18][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][14] .is_wysiwyg = "true";
defparam \Reg[18][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N28
cycloneive_lcell_comb \Reg[22][14]~feeder (
// Equation(s):
// \Reg[22][14]~feeder_combout  = \wdat~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat11),
	.cin(gnd),
	.combout(\Reg[22][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[22][14]~feeder .lut_mask = 16'hFF00;
defparam \Reg[22][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y36_N29
dffeas \Reg[22][14] (
	.clk(!CLK),
	.d(\Reg[22][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][14] .is_wysiwyg = "true";
defparam \Reg[22][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N2
cycloneive_lcell_comb \Mux17~2 (
// Equation(s):
// \Mux17~2_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[22][14]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[18][14]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[18][14]~q ),
	.datad(\Reg[22][14]~q ),
	.cin(gnd),
	.combout(\Mux17~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~2 .lut_mask = 16'hDC98;
defparam \Mux17~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N12
cycloneive_lcell_comb \Mux17~3 (
// Equation(s):
// \Mux17~3_combout  = (ifid_ifinstr_o_24 & ((\Mux17~2_combout  & (\Reg[30][14]~q )) # (!\Mux17~2_combout  & ((\Reg[26][14]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux17~2_combout ))))

	.dataa(\Reg[30][14]~q ),
	.datab(\Reg[26][14]~q ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Mux17~2_combout ),
	.cin(gnd),
	.combout(\Mux17~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~3 .lut_mask = 16'hAFC0;
defparam \Mux17~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N26
cycloneive_lcell_comb \Mux17~6 (
// Equation(s):
// \Mux17~6_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Mux17~3_combout ))) # (!ifid_ifinstr_o_22 & (\Mux17~5_combout ))))

	.dataa(\Mux17~5_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux17~3_combout ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux17~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~6 .lut_mask = 16'hFC22;
defparam \Mux17~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y29_N31
dffeas \Reg[31][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][14] .is_wysiwyg = "true";
defparam \Reg[31][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N29
dffeas \Reg[23][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][14] .is_wysiwyg = "true";
defparam \Reg[23][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N11
dffeas \Reg[19][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][14] .is_wysiwyg = "true";
defparam \Reg[19][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N24
cycloneive_lcell_comb \Reg[27][14]~feeder (
// Equation(s):
// \Reg[27][14]~feeder_combout  = \wdat~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat11),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[27][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[27][14]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[27][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y29_N25
dffeas \Reg[27][14] (
	.clk(!CLK),
	.d(\Reg[27][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][14] .is_wysiwyg = "true";
defparam \Reg[27][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N10
cycloneive_lcell_comb \Mux17~7 (
// Equation(s):
// \Mux17~7_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[27][14]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & (\Reg[19][14]~q )))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[19][14]~q ),
	.datad(\Reg[27][14]~q ),
	.cin(gnd),
	.combout(\Mux17~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~7 .lut_mask = 16'hBA98;
defparam \Mux17~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N28
cycloneive_lcell_comb \Mux17~8 (
// Equation(s):
// \Mux17~8_combout  = (ifid_ifinstr_o_23 & ((\Mux17~7_combout  & (\Reg[31][14]~q )) # (!\Mux17~7_combout  & ((\Reg[23][14]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux17~7_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[31][14]~q ),
	.datac(\Reg[23][14]~q ),
	.datad(\Mux17~7_combout ),
	.cin(gnd),
	.combout(\Mux17~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~8 .lut_mask = 16'hDDA0;
defparam \Mux17~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y38_N25
dffeas \Reg[15][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][14] .is_wysiwyg = "true";
defparam \Reg[15][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N1
dffeas \Reg[14][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][14] .is_wysiwyg = "true";
defparam \Reg[14][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N17
dffeas \Reg[13][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][14] .is_wysiwyg = "true";
defparam \Reg[13][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N7
dffeas \Reg[12][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][14] .is_wysiwyg = "true";
defparam \Reg[12][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N6
cycloneive_lcell_comb \Mux17~17 (
// Equation(s):
// \Mux17~17_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[13][14]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[12][14]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[13][14]~q ),
	.datac(\Reg[12][14]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux17~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~17 .lut_mask = 16'hEE50;
defparam \Mux17~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N0
cycloneive_lcell_comb \Mux17~18 (
// Equation(s):
// \Mux17~18_combout  = (ifid_ifinstr_o_22 & ((\Mux17~17_combout  & (\Reg[15][14]~q )) # (!\Mux17~17_combout  & ((\Reg[14][14]~q ))))) # (!ifid_ifinstr_o_22 & (((\Mux17~17_combout ))))

	.dataa(\Reg[15][14]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[14][14]~q ),
	.datad(\Mux17~17_combout ),
	.cin(gnd),
	.combout(\Mux17~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~18 .lut_mask = 16'hBBC0;
defparam \Mux17~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N31
dffeas \Reg[7][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][14] .is_wysiwyg = "true";
defparam \Reg[7][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y39_N17
dffeas \Reg[6][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][14] .is_wysiwyg = "true";
defparam \Reg[6][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y39_N9
dffeas \Reg[5][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][14] .is_wysiwyg = "true";
defparam \Reg[5][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y39_N11
dffeas \Reg[4][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][14] .is_wysiwyg = "true";
defparam \Reg[4][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N8
cycloneive_lcell_comb \Mux17~10 (
// Equation(s):
// \Mux17~10_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[5][14]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[4][14]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[5][14]~q ),
	.datad(\Reg[4][14]~q ),
	.cin(gnd),
	.combout(\Mux17~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~10 .lut_mask = 16'hD9C8;
defparam \Mux17~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N16
cycloneive_lcell_comb \Mux17~11 (
// Equation(s):
// \Mux17~11_combout  = (ifid_ifinstr_o_22 & ((\Mux17~10_combout  & (\Reg[7][14]~q )) # (!\Mux17~10_combout  & ((\Reg[6][14]~q ))))) # (!ifid_ifinstr_o_22 & (((\Mux17~10_combout ))))

	.dataa(\Reg[7][14]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[6][14]~q ),
	.datad(\Mux17~10_combout ),
	.cin(gnd),
	.combout(\Mux17~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~11 .lut_mask = 16'hBBC0;
defparam \Mux17~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y36_N19
dffeas \Reg[8][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][14] .is_wysiwyg = "true";
defparam \Reg[8][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N25
dffeas \Reg[10][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][14] .is_wysiwyg = "true";
defparam \Reg[10][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N18
cycloneive_lcell_comb \Mux17~12 (
// Equation(s):
// \Mux17~12_combout  = (ifid_ifinstr_o_21 & (ifid_ifinstr_o_22)) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[10][14]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[8][14]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[8][14]~q ),
	.datad(\Reg[10][14]~q ),
	.cin(gnd),
	.combout(\Mux17~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~12 .lut_mask = 16'hDC98;
defparam \Mux17~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N7
dffeas \Reg[11][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][14] .is_wysiwyg = "true";
defparam \Reg[11][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y35_N21
dffeas \Reg[9][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][14] .is_wysiwyg = "true";
defparam \Reg[9][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N6
cycloneive_lcell_comb \Mux17~13 (
// Equation(s):
// \Mux17~13_combout  = (ifid_ifinstr_o_21 & ((\Mux17~12_combout  & (\Reg[11][14]~q )) # (!\Mux17~12_combout  & ((\Reg[9][14]~q ))))) # (!ifid_ifinstr_o_21 & (\Mux17~12_combout ))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux17~12_combout ),
	.datac(\Reg[11][14]~q ),
	.datad(\Reg[9][14]~q ),
	.cin(gnd),
	.combout(\Mux17~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~13 .lut_mask = 16'hE6C4;
defparam \Mux17~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N4
cycloneive_lcell_comb \Reg[2][14]~feeder (
// Equation(s):
// \Reg[2][14]~feeder_combout  = \wdat~25_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat11),
	.cin(gnd),
	.combout(\Reg[2][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[2][14]~feeder .lut_mask = 16'hFF00;
defparam \Reg[2][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y36_N5
dffeas \Reg[2][14] (
	.clk(!CLK),
	.d(\Reg[2][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][14] .is_wysiwyg = "true";
defparam \Reg[2][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N25
dffeas \Reg[3][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][14] .is_wysiwyg = "true";
defparam \Reg[3][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N11
dffeas \Reg[1][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][14] .is_wysiwyg = "true";
defparam \Reg[1][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N24
cycloneive_lcell_comb \Mux17~14 (
// Equation(s):
// \Mux17~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[3][14]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[1][14]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[3][14]~q ),
	.datad(\Reg[1][14]~q ),
	.cin(gnd),
	.combout(\Mux17~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~14 .lut_mask = 16'hA280;
defparam \Mux17~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N6
cycloneive_lcell_comb \Mux17~15 (
// Equation(s):
// \Mux17~15_combout  = (\Mux17~14_combout ) # ((!ifid_ifinstr_o_21 & (\Reg[2][14]~q  & ifid_ifinstr_o_22)))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[2][14]~q ),
	.datac(\Mux17~14_combout ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux17~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~15 .lut_mask = 16'hF4F0;
defparam \Mux17~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N0
cycloneive_lcell_comb \Mux17~16 (
// Equation(s):
// \Mux17~16_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Mux17~13_combout )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & ((\Mux17~15_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Mux17~13_combout ),
	.datad(\Mux17~15_combout ),
	.cin(gnd),
	.combout(\Mux17~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~16 .lut_mask = 16'hB9A8;
defparam \Mux17~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N19
dffeas \Reg[19][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][13] .is_wysiwyg = "true";
defparam \Reg[19][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y29_N13
dffeas \Reg[23][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][13] .is_wysiwyg = "true";
defparam \Reg[23][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N12
cycloneive_lcell_comb \Mux18~7 (
// Equation(s):
// \Mux18~7_combout  = (ifid_ifinstr_o_23 & (((\Reg[23][13]~q ) # (ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (\Reg[19][13]~q  & ((!ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[19][13]~q ),
	.datac(\Reg[23][13]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux18~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~7 .lut_mask = 16'hAAE4;
defparam \Mux18~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N0
cycloneive_lcell_comb \Reg[27][13]~feeder (
// Equation(s):
// \Reg[27][13]~feeder_combout  = \wdat~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat12),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[27][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[27][13]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[27][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N1
dffeas \Reg[27][13] (
	.clk(!CLK),
	.d(\Reg[27][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][13] .is_wysiwyg = "true";
defparam \Reg[27][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y29_N3
dffeas \Reg[31][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][13] .is_wysiwyg = "true";
defparam \Reg[31][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N2
cycloneive_lcell_comb \Mux18~8 (
// Equation(s):
// \Mux18~8_combout  = (\Mux18~7_combout  & (((\Reg[31][13]~q ) # (!ifid_ifinstr_o_24)))) # (!\Mux18~7_combout  & (\Reg[27][13]~q  & ((ifid_ifinstr_o_24))))

	.dataa(\Mux18~7_combout ),
	.datab(\Reg[27][13]~q ),
	.datac(\Reg[31][13]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux18~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~8 .lut_mask = 16'hE4AA;
defparam \Mux18~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N8
cycloneive_lcell_comb \Reg[21][13]~feeder (
// Equation(s):
// \Reg[21][13]~feeder_combout  = \wdat~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat12),
	.cin(gnd),
	.combout(\Reg[21][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[21][13]~feeder .lut_mask = 16'hFF00;
defparam \Reg[21][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y38_N9
dffeas \Reg[21][13] (
	.clk(!CLK),
	.d(\Reg[21][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][13] .is_wysiwyg = "true";
defparam \Reg[21][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N27
dffeas \Reg[17][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][13] .is_wysiwyg = "true";
defparam \Reg[17][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N26
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// \Mux18~0_combout  = (ifid_ifinstr_o_23 & ((\Reg[21][13]~q ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((\Reg[17][13]~q  & !ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[21][13]~q ),
	.datac(\Reg[17][13]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'hAAD8;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N22
cycloneive_lcell_comb \Reg[29][13]~feeder (
// Equation(s):
// \Reg[29][13]~feeder_combout  = \wdat~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat12),
	.cin(gnd),
	.combout(\Reg[29][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[29][13]~feeder .lut_mask = 16'hFF00;
defparam \Reg[29][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y38_N23
dffeas \Reg[29][13] (
	.clk(!CLK),
	.d(\Reg[29][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][13] .is_wysiwyg = "true";
defparam \Reg[29][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N16
cycloneive_lcell_comb \Reg[25][13]~feeder (
// Equation(s):
// \Reg[25][13]~feeder_combout  = \wdat~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat12),
	.cin(gnd),
	.combout(\Reg[25][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][13]~feeder .lut_mask = 16'hFF00;
defparam \Reg[25][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N17
dffeas \Reg[25][13] (
	.clk(!CLK),
	.d(\Reg[25][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][13] .is_wysiwyg = "true";
defparam \Reg[25][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N24
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// \Mux18~1_combout  = (ifid_ifinstr_o_24 & ((\Mux18~0_combout  & (\Reg[29][13]~q )) # (!\Mux18~0_combout  & ((\Reg[25][13]~q ))))) # (!ifid_ifinstr_o_24 & (\Mux18~0_combout ))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux18~0_combout ),
	.datac(\Reg[29][13]~q ),
	.datad(\Reg[25][13]~q ),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'hE6C4;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N18
cycloneive_lcell_comb \Reg[16][13]~feeder (
// Equation(s):
// \Reg[16][13]~feeder_combout  = \wdat~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat12),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[16][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[16][13]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[16][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N19
dffeas \Reg[16][13] (
	.clk(!CLK),
	.d(\Reg[16][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][13] .is_wysiwyg = "true";
defparam \Reg[16][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N9
dffeas \Reg[24][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][13] .is_wysiwyg = "true";
defparam \Reg[24][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N8
cycloneive_lcell_comb \Mux18~4 (
// Equation(s):
// \Mux18~4_combout  = (ifid_ifinstr_o_24 & (((\Reg[24][13]~q ) # (ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & (\Reg[16][13]~q  & ((!ifid_ifinstr_o_23))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[16][13]~q ),
	.datac(\Reg[24][13]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux18~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~4 .lut_mask = 16'hAAE4;
defparam \Mux18~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N20
cycloneive_lcell_comb \Reg[20][13]~feeder (
// Equation(s):
// \Reg[20][13]~feeder_combout  = \wdat~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat12),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[20][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[20][13]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[20][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N21
dffeas \Reg[20][13] (
	.clk(!CLK),
	.d(\Reg[20][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][13] .is_wysiwyg = "true";
defparam \Reg[20][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N16
cycloneive_lcell_comb \Mux18~5 (
// Equation(s):
// \Mux18~5_combout  = (ifid_ifinstr_o_23 & ((\Mux18~4_combout  & (\Reg[28][13]~q )) # (!\Mux18~4_combout  & ((\Reg[20][13]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux18~4_combout ))))

	.dataa(\Reg[28][13]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Mux18~4_combout ),
	.datad(\Reg[20][13]~q ),
	.cin(gnd),
	.combout(\Mux18~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~5 .lut_mask = 16'hBCB0;
defparam \Mux18~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N16
cycloneive_lcell_comb \Reg[30][13]~feeder (
// Equation(s):
// \Reg[30][13]~feeder_combout  = \wdat~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat12),
	.cin(gnd),
	.combout(\Reg[30][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[30][13]~feeder .lut_mask = 16'hFF00;
defparam \Reg[30][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y36_N17
dffeas \Reg[30][13] (
	.clk(!CLK),
	.d(\Reg[30][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][13] .is_wysiwyg = "true";
defparam \Reg[30][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y30_N9
dffeas \Reg[26][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][13] .is_wysiwyg = "true";
defparam \Reg[26][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y30_N11
dffeas \Reg[18][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][13] .is_wysiwyg = "true";
defparam \Reg[18][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N8
cycloneive_lcell_comb \Mux18~2 (
// Equation(s):
// \Mux18~2_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[26][13]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & ((\Reg[18][13]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[26][13]~q ),
	.datad(\Reg[18][13]~q ),
	.cin(gnd),
	.combout(\Mux18~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~2 .lut_mask = 16'hB9A8;
defparam \Mux18~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N14
cycloneive_lcell_comb \Mux18~3 (
// Equation(s):
// \Mux18~3_combout  = (ifid_ifinstr_o_23 & ((\Mux18~2_combout  & ((\Reg[30][13]~q ))) # (!\Mux18~2_combout  & (\Reg[22][13]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux18~2_combout ))))

	.dataa(\Reg[22][13]~q ),
	.datab(\Reg[30][13]~q ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux18~2_combout ),
	.cin(gnd),
	.combout(\Mux18~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~3 .lut_mask = 16'hCFA0;
defparam \Mux18~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N28
cycloneive_lcell_comb \Mux18~6 (
// Equation(s):
// \Mux18~6_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Mux18~3_combout ))) # (!ifid_ifinstr_o_22 & (\Mux18~5_combout ))))

	.dataa(\Mux18~5_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux18~3_combout ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux18~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~6 .lut_mask = 16'hFC22;
defparam \Mux18~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y36_N25
dffeas \Reg[3][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][13] .is_wysiwyg = "true";
defparam \Reg[3][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N3
dffeas \Reg[1][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][13] .is_wysiwyg = "true";
defparam \Reg[1][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N24
cycloneive_lcell_comb \Mux18~14 (
// Equation(s):
// \Mux18~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[3][13]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[1][13]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[3][13]~q ),
	.datad(\Reg[1][13]~q ),
	.cin(gnd),
	.combout(\Mux18~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~14 .lut_mask = 16'hC480;
defparam \Mux18~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N29
dffeas \Reg[2][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][13] .is_wysiwyg = "true";
defparam \Reg[2][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N8
cycloneive_lcell_comb \Mux18~15 (
// Equation(s):
// \Mux18~15_combout  = (\Mux18~14_combout ) # ((ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & \Reg[2][13]~q )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux18~14_combout ),
	.datad(\Reg[2][13]~q ),
	.cin(gnd),
	.combout(\Mux18~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~15 .lut_mask = 16'hF2F0;
defparam \Mux18~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N27
dffeas \Reg[7][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][13] .is_wysiwyg = "true";
defparam \Reg[7][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y39_N21
dffeas \Reg[6][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][13] .is_wysiwyg = "true";
defparam \Reg[6][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N26
cycloneive_lcell_comb \Mux18~13 (
// Equation(s):
// \Mux18~13_combout  = (\Mux18~12_combout  & (((\Reg[7][13]~q )) # (!ifid_ifinstr_o_22))) # (!\Mux18~12_combout  & (ifid_ifinstr_o_22 & ((\Reg[6][13]~q ))))

	.dataa(\Mux18~12_combout ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[7][13]~q ),
	.datad(\Reg[6][13]~q ),
	.cin(gnd),
	.combout(\Mux18~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~13 .lut_mask = 16'hE6A2;
defparam \Mux18~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N10
cycloneive_lcell_comb \Mux18~16 (
// Equation(s):
// \Mux18~16_combout  = (ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24) # ((\Mux18~13_combout )))) # (!ifid_ifinstr_o_23 & (!ifid_ifinstr_o_24 & (\Mux18~15_combout )))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Mux18~15_combout ),
	.datad(\Mux18~13_combout ),
	.cin(gnd),
	.combout(\Mux18~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~16 .lut_mask = 16'hBA98;
defparam \Mux18~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N15
dffeas \Reg[14][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][13] .is_wysiwyg = "true";
defparam \Reg[14][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N12
cycloneive_lcell_comb \Reg[15][13]~feeder (
// Equation(s):
// \Reg[15][13]~feeder_combout  = \wdat~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat12),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[15][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[15][13]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[15][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y28_N13
dffeas \Reg[15][13] (
	.clk(!CLK),
	.d(\Reg[15][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][13] .is_wysiwyg = "true";
defparam \Reg[15][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N9
dffeas \Reg[13][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][13] .is_wysiwyg = "true";
defparam \Reg[13][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N11
dffeas \Reg[12][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][13] .is_wysiwyg = "true";
defparam \Reg[12][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N10
cycloneive_lcell_comb \Mux18~17 (
// Equation(s):
// \Mux18~17_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[13][13]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[12][13]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[13][13]~q ),
	.datac(\Reg[12][13]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux18~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~17 .lut_mask = 16'hEE50;
defparam \Mux18~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N8
cycloneive_lcell_comb \Mux18~18 (
// Equation(s):
// \Mux18~18_combout  = (ifid_ifinstr_o_22 & ((\Mux18~17_combout  & ((\Reg[15][13]~q ))) # (!\Mux18~17_combout  & (\Reg[14][13]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux18~17_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[14][13]~q ),
	.datac(\Reg[15][13]~q ),
	.datad(\Mux18~17_combout ),
	.cin(gnd),
	.combout(\Mux18~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~18 .lut_mask = 16'hF588;
defparam \Mux18~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y36_N13
dffeas \Reg[10][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][13] .is_wysiwyg = "true";
defparam \Reg[10][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N7
dffeas \Reg[8][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][13] .is_wysiwyg = "true";
defparam \Reg[8][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N12
cycloneive_lcell_comb \Mux18~10 (
// Equation(s):
// \Mux18~10_combout  = (ifid_ifinstr_o_21 & (ifid_ifinstr_o_22)) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[10][13]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[8][13]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[10][13]~q ),
	.datad(\Reg[8][13]~q ),
	.cin(gnd),
	.combout(\Mux18~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~10 .lut_mask = 16'hD9C8;
defparam \Mux18~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N1
dffeas \Reg[9][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][13] .is_wysiwyg = "true";
defparam \Reg[9][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y36_N31
dffeas \Reg[11][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][13] .is_wysiwyg = "true";
defparam \Reg[11][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N0
cycloneive_lcell_comb \Mux18~11 (
// Equation(s):
// \Mux18~11_combout  = (\Mux18~10_combout  & (((\Reg[11][13]~q )) # (!ifid_ifinstr_o_21))) # (!\Mux18~10_combout  & (ifid_ifinstr_o_21 & (\Reg[9][13]~q )))

	.dataa(\Mux18~10_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[9][13]~q ),
	.datad(\Reg[11][13]~q ),
	.cin(gnd),
	.combout(\Mux18~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~11 .lut_mask = 16'hEA62;
defparam \Mux18~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N30
cycloneive_lcell_comb \Reg[25][12]~feeder (
// Equation(s):
// \Reg[25][12]~feeder_combout  = \wdat~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat13),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[25][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][12]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[25][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N31
dffeas \Reg[25][12] (
	.clk(!CLK),
	.d(\Reg[25][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][12] .is_wysiwyg = "true";
defparam \Reg[25][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N17
dffeas \Reg[17][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][12] .is_wysiwyg = "true";
defparam \Reg[17][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N16
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[25][12]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[17][12]~q )))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[25][12]~q ),
	.datac(\Reg[17][12]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'hEE50;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y37_N15
dffeas \Reg[29][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][12] .is_wysiwyg = "true";
defparam \Reg[29][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y37_N23
dffeas \Reg[21][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][12] .is_wysiwyg = "true";
defparam \Reg[21][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N14
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// \Mux19~1_combout  = (ifid_ifinstr_o_23 & ((\Mux19~0_combout  & (\Reg[29][12]~q )) # (!\Mux19~0_combout  & ((\Reg[21][12]~q ))))) # (!ifid_ifinstr_o_23 & (\Mux19~0_combout ))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux19~0_combout ),
	.datac(\Reg[29][12]~q ),
	.datad(\Reg[21][12]~q ),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'hE6C4;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y29_N27
dffeas \Reg[31][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][12] .is_wysiwyg = "true";
defparam \Reg[31][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N17
dffeas \Reg[23][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][12] .is_wysiwyg = "true";
defparam \Reg[23][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N31
dffeas \Reg[19][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][12] .is_wysiwyg = "true";
defparam \Reg[19][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N28
cycloneive_lcell_comb \Reg[27][12]~feeder (
// Equation(s):
// \Reg[27][12]~feeder_combout  = \wdat~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat13),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[27][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[27][12]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[27][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y29_N29
dffeas \Reg[27][12] (
	.clk(!CLK),
	.d(\Reg[27][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][12] .is_wysiwyg = "true";
defparam \Reg[27][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N30
cycloneive_lcell_comb \Mux19~7 (
// Equation(s):
// \Mux19~7_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[27][12]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & (\Reg[19][12]~q )))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[19][12]~q ),
	.datad(\Reg[27][12]~q ),
	.cin(gnd),
	.combout(\Mux19~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~7 .lut_mask = 16'hBA98;
defparam \Mux19~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N22
cycloneive_lcell_comb \Mux19~8 (
// Equation(s):
// \Mux19~8_combout  = (ifid_ifinstr_o_23 & ((\Mux19~7_combout  & (\Reg[31][12]~q )) # (!\Mux19~7_combout  & ((\Reg[23][12]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux19~7_combout ))))

	.dataa(\Reg[31][12]~q ),
	.datab(\Reg[23][12]~q ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux19~7_combout ),
	.cin(gnd),
	.combout(\Mux19~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~8 .lut_mask = 16'hAFC0;
defparam \Mux19~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y36_N9
dffeas \Reg[22][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][12] .is_wysiwyg = "true";
defparam \Reg[22][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N8
cycloneive_lcell_comb \Mux19~2 (
// Equation(s):
// \Mux19~2_combout  = (ifid_ifinstr_o_23 & (((\Reg[22][12]~q ) # (ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (\Reg[18][12]~q  & ((!ifid_ifinstr_o_24))))

	.dataa(\Reg[18][12]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[22][12]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~2 .lut_mask = 16'hCCE2;
defparam \Mux19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y36_N23
dffeas \Reg[30][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][12] .is_wysiwyg = "true";
defparam \Reg[30][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N24
cycloneive_lcell_comb \Reg[26][12]~feeder (
// Equation(s):
// \Reg[26][12]~feeder_combout  = \wdat~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat13),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[26][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[26][12]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[26][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N25
dffeas \Reg[26][12] (
	.clk(!CLK),
	.d(\Reg[26][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][12] .is_wysiwyg = "true";
defparam \Reg[26][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N22
cycloneive_lcell_comb \Mux19~3 (
// Equation(s):
// \Mux19~3_combout  = (ifid_ifinstr_o_24 & ((\Mux19~2_combout  & (\Reg[30][12]~q )) # (!\Mux19~2_combout  & ((\Reg[26][12]~q ))))) # (!ifid_ifinstr_o_24 & (\Mux19~2_combout ))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux19~2_combout ),
	.datac(\Reg[30][12]~q ),
	.datad(\Reg[26][12]~q ),
	.cin(gnd),
	.combout(\Mux19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~3 .lut_mask = 16'hE6C4;
defparam \Mux19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y34_N13
dffeas \Reg[20][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][12] .is_wysiwyg = "true";
defparam \Reg[20][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N23
dffeas \Reg[16][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][12] .is_wysiwyg = "true";
defparam \Reg[16][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N12
cycloneive_lcell_comb \Mux19~4 (
// Equation(s):
// \Mux19~4_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & (\Reg[20][12]~q )) # (!ifid_ifinstr_o_23 & ((\Reg[16][12]~q )))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[20][12]~q ),
	.datad(\Reg[16][12]~q ),
	.cin(gnd),
	.combout(\Mux19~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~4 .lut_mask = 16'hD9C8;
defparam \Mux19~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y34_N27
dffeas \Reg[28][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][12] .is_wysiwyg = "true";
defparam \Reg[28][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N24
cycloneive_lcell_comb \Mux19~5 (
// Equation(s):
// \Mux19~5_combout  = (ifid_ifinstr_o_24 & ((\Mux19~4_combout  & ((\Reg[28][12]~q ))) # (!\Mux19~4_combout  & (\Reg[24][12]~q )))) # (!ifid_ifinstr_o_24 & (((\Mux19~4_combout ))))

	.dataa(\Reg[24][12]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Mux19~4_combout ),
	.datad(\Reg[28][12]~q ),
	.cin(gnd),
	.combout(\Mux19~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~5 .lut_mask = 16'hF838;
defparam \Mux19~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N28
cycloneive_lcell_comb \Mux19~6 (
// Equation(s):
// \Mux19~6_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Mux19~3_combout )) # (!ifid_ifinstr_o_22 & ((\Mux19~5_combout )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux19~3_combout ),
	.datac(\Mux19~5_combout ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux19~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~6 .lut_mask = 16'hEE50;
defparam \Mux19~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N24
cycloneive_lcell_comb \Reg[15][12]~feeder (
// Equation(s):
// \Reg[15][12]~feeder_combout  = \wdat~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat13),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[15][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[15][12]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[15][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N25
dffeas \Reg[15][12] (
	.clk(!CLK),
	.d(\Reg[15][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][12] .is_wysiwyg = "true";
defparam \Reg[15][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N7
dffeas \Reg[14][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][12] .is_wysiwyg = "true";
defparam \Reg[14][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N1
dffeas \Reg[13][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][12] .is_wysiwyg = "true";
defparam \Reg[13][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N7
dffeas \Reg[12][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][12] .is_wysiwyg = "true";
defparam \Reg[12][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N6
cycloneive_lcell_comb \Mux19~17 (
// Equation(s):
// \Mux19~17_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[13][12]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[12][12]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[13][12]~q ),
	.datac(\Reg[12][12]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux19~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~17 .lut_mask = 16'hEE50;
defparam \Mux19~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N6
cycloneive_lcell_comb \Mux19~18 (
// Equation(s):
// \Mux19~18_combout  = (ifid_ifinstr_o_22 & ((\Mux19~17_combout  & (\Reg[15][12]~q )) # (!\Mux19~17_combout  & ((\Reg[14][12]~q ))))) # (!ifid_ifinstr_o_22 & (((\Mux19~17_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[15][12]~q ),
	.datac(\Reg[14][12]~q ),
	.datad(\Mux19~17_combout ),
	.cin(gnd),
	.combout(\Mux19~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~18 .lut_mask = 16'hDDA0;
defparam \Mux19~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y39_N1
dffeas \Reg[5][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][12] .is_wysiwyg = "true";
defparam \Reg[5][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y39_N7
dffeas \Reg[4][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][12] .is_wysiwyg = "true";
defparam \Reg[4][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N0
cycloneive_lcell_comb \Mux19~10 (
// Equation(s):
// \Mux19~10_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[5][12]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[4][12]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[5][12]~q ),
	.datad(\Reg[4][12]~q ),
	.cin(gnd),
	.combout(\Mux19~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~10 .lut_mask = 16'hD9C8;
defparam \Mux19~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y39_N1
dffeas \Reg[6][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][12] .is_wysiwyg = "true";
defparam \Reg[6][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N3
dffeas \Reg[7][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][12] .is_wysiwyg = "true";
defparam \Reg[7][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N0
cycloneive_lcell_comb \Mux19~11 (
// Equation(s):
// \Mux19~11_combout  = (ifid_ifinstr_o_22 & ((\Mux19~10_combout  & ((\Reg[7][12]~q ))) # (!\Mux19~10_combout  & (\Reg[6][12]~q )))) # (!ifid_ifinstr_o_22 & (\Mux19~10_combout ))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Mux19~10_combout ),
	.datac(\Reg[6][12]~q ),
	.datad(\Reg[7][12]~q ),
	.cin(gnd),
	.combout(\Mux19~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~11 .lut_mask = 16'hEC64;
defparam \Mux19~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N29
dffeas \Reg[9][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][12] .is_wysiwyg = "true";
defparam \Reg[9][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N31
dffeas \Reg[11][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][12] .is_wysiwyg = "true";
defparam \Reg[11][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N23
dffeas \Reg[8][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][12] .is_wysiwyg = "true";
defparam \Reg[8][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N29
dffeas \Reg[10][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][12] .is_wysiwyg = "true";
defparam \Reg[10][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N22
cycloneive_lcell_comb \Mux19~12 (
// Equation(s):
// \Mux19~12_combout  = (ifid_ifinstr_o_21 & (ifid_ifinstr_o_22)) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[10][12]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[8][12]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[8][12]~q ),
	.datad(\Reg[10][12]~q ),
	.cin(gnd),
	.combout(\Mux19~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~12 .lut_mask = 16'hDC98;
defparam \Mux19~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N30
cycloneive_lcell_comb \Mux19~13 (
// Equation(s):
// \Mux19~13_combout  = (ifid_ifinstr_o_21 & ((\Mux19~12_combout  & ((\Reg[11][12]~q ))) # (!\Mux19~12_combout  & (\Reg[9][12]~q )))) # (!ifid_ifinstr_o_21 & (((\Mux19~12_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[9][12]~q ),
	.datac(\Reg[11][12]~q ),
	.datad(\Mux19~12_combout ),
	.cin(gnd),
	.combout(\Mux19~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~13 .lut_mask = 16'hF588;
defparam \Mux19~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N19
dffeas \Reg[2][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][12] .is_wysiwyg = "true";
defparam \Reg[2][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N13
dffeas \Reg[3][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][12] .is_wysiwyg = "true";
defparam \Reg[3][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N3
dffeas \Reg[1][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][12] .is_wysiwyg = "true";
defparam \Reg[1][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N12
cycloneive_lcell_comb \Mux19~14 (
// Equation(s):
// \Mux19~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[3][12]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[1][12]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[3][12]~q ),
	.datad(\Reg[1][12]~q ),
	.cin(gnd),
	.combout(\Mux19~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~14 .lut_mask = 16'hA280;
defparam \Mux19~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N10
cycloneive_lcell_comb \Mux19~15 (
// Equation(s):
// \Mux19~15_combout  = (\Mux19~14_combout ) # ((ifid_ifinstr_o_22 & (\Reg[2][12]~q  & !ifid_ifinstr_o_21)))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[2][12]~q ),
	.datac(\Mux19~14_combout ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux19~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~15 .lut_mask = 16'hF0F8;
defparam \Mux19~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N16
cycloneive_lcell_comb \Mux19~16 (
// Equation(s):
// \Mux19~16_combout  = (ifid_ifinstr_o_24 & ((\Mux19~13_combout ) # ((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & (((!ifid_ifinstr_o_23 & \Mux19~15_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux19~13_combout ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux19~15_combout ),
	.cin(gnd),
	.combout(\Mux19~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~16 .lut_mask = 16'hADA8;
defparam \Mux19~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N24
cycloneive_lcell_comb \Reg[20][11]~feeder (
// Equation(s):
// \Reg[20][11]~feeder_combout  = \wdat~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat14),
	.cin(gnd),
	.combout(\Reg[20][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[20][11]~feeder .lut_mask = 16'hFF00;
defparam \Reg[20][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N25
dffeas \Reg[20][11] (
	.clk(!CLK),
	.d(\Reg[20][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][11] .is_wysiwyg = "true";
defparam \Reg[20][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N23
dffeas \Reg[28][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][11] .is_wysiwyg = "true";
defparam \Reg[28][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N30
cycloneive_lcell_comb \Mux20~5 (
// Equation(s):
// \Mux20~5_combout  = (\Mux20~4_combout  & (((\Reg[28][11]~q ) # (!ifid_ifinstr_o_23)))) # (!\Mux20~4_combout  & (\Reg[20][11]~q  & (ifid_ifinstr_o_23)))

	.dataa(\Mux20~4_combout ),
	.datab(\Reg[20][11]~q ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Reg[28][11]~q ),
	.cin(gnd),
	.combout(\Mux20~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~5 .lut_mask = 16'hEA4A;
defparam \Mux20~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N19
dffeas \Reg[18][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][11] .is_wysiwyg = "true";
defparam \Reg[18][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y30_N13
dffeas \Reg[26][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][11] .is_wysiwyg = "true";
defparam \Reg[26][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N12
cycloneive_lcell_comb \Mux20~2 (
// Equation(s):
// \Mux20~2_combout  = (ifid_ifinstr_o_24 & (((\Reg[26][11]~q ) # (ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & (\Reg[18][11]~q  & ((!ifid_ifinstr_o_23))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[18][11]~q ),
	.datac(\Reg[26][11]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux20~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~2 .lut_mask = 16'hAAE4;
defparam \Mux20~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N28
cycloneive_lcell_comb \Reg[30][11]~feeder (
// Equation(s):
// \Reg[30][11]~feeder_combout  = \wdat~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat14),
	.cin(gnd),
	.combout(\Reg[30][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[30][11]~feeder .lut_mask = 16'hFF00;
defparam \Reg[30][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N29
dffeas \Reg[30][11] (
	.clk(!CLK),
	.d(\Reg[30][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][11] .is_wysiwyg = "true";
defparam \Reg[30][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N2
cycloneive_lcell_comb \Mux20~3 (
// Equation(s):
// \Mux20~3_combout  = (\Mux20~2_combout  & (((\Reg[30][11]~q ) # (!ifid_ifinstr_o_23)))) # (!\Mux20~2_combout  & (\Reg[22][11]~q  & (ifid_ifinstr_o_23)))

	.dataa(\Reg[22][11]~q ),
	.datab(\Mux20~2_combout ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Reg[30][11]~q ),
	.cin(gnd),
	.combout(\Mux20~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~3 .lut_mask = 16'hEC2C;
defparam \Mux20~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N6
cycloneive_lcell_comb \Mux20~6 (
// Equation(s):
// \Mux20~6_combout  = (ifid_ifinstr_o_22 & (((\Mux20~3_combout ) # (ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & (\Mux20~5_combout  & ((!ifid_ifinstr_o_21))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Mux20~5_combout ),
	.datac(\Mux20~3_combout ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux20~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~6 .lut_mask = 16'hAAE4;
defparam \Mux20~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y37_N31
dffeas \Reg[29][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][11] .is_wysiwyg = "true";
defparam \Reg[29][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N21
dffeas \Reg[17][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][11] .is_wysiwyg = "true";
defparam \Reg[17][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N0
cycloneive_lcell_comb \Reg[21][11]~feeder (
// Equation(s):
// \Reg[21][11]~feeder_combout  = \wdat~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat14),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[21][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[21][11]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[21][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N1
dffeas \Reg[21][11] (
	.clk(!CLK),
	.d(\Reg[21][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][11] .is_wysiwyg = "true";
defparam \Reg[21][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N10
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// \Mux20~0_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[21][11]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[17][11]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[17][11]~q ),
	.datad(\Reg[21][11]~q ),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'hDC98;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N0
cycloneive_lcell_comb \Reg[25][11]~feeder (
// Equation(s):
// \Reg[25][11]~feeder_combout  = \wdat~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat14),
	.cin(gnd),
	.combout(\Reg[25][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][11]~feeder .lut_mask = 16'hFF00;
defparam \Reg[25][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y32_N1
dffeas \Reg[25][11] (
	.clk(!CLK),
	.d(\Reg[25][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][11] .is_wysiwyg = "true";
defparam \Reg[25][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N22
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// \Mux20~1_combout  = (ifid_ifinstr_o_24 & ((\Mux20~0_combout  & (\Reg[29][11]~q )) # (!\Mux20~0_combout  & ((\Reg[25][11]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux20~0_combout ))))

	.dataa(\Reg[29][11]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Mux20~0_combout ),
	.datad(\Reg[25][11]~q ),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'hBCB0;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N15
dffeas \Reg[31][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][11] .is_wysiwyg = "true";
defparam \Reg[31][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N20
cycloneive_lcell_comb \Reg[23][11]~feeder (
// Equation(s):
// \Reg[23][11]~feeder_combout  = \wdat~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat14),
	.cin(gnd),
	.combout(\Reg[23][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[23][11]~feeder .lut_mask = 16'hFF00;
defparam \Reg[23][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N21
dffeas \Reg[23][11] (
	.clk(!CLK),
	.d(\Reg[23][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][11] .is_wysiwyg = "true";
defparam \Reg[23][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N22
cycloneive_lcell_comb \Reg[19][11]~feeder (
// Equation(s):
// \Reg[19][11]~feeder_combout  = \wdat~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat14),
	.cin(gnd),
	.combout(\Reg[19][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[19][11]~feeder .lut_mask = 16'hFF00;
defparam \Reg[19][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N23
dffeas \Reg[19][11] (
	.clk(!CLK),
	.d(\Reg[19][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][11] .is_wysiwyg = "true";
defparam \Reg[19][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N8
cycloneive_lcell_comb \Mux20~7 (
// Equation(s):
// \Mux20~7_combout  = (ifid_ifinstr_o_23 & ((\Reg[23][11]~q ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((\Reg[19][11]~q  & !ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[23][11]~q ),
	.datac(\Reg[19][11]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux20~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~7 .lut_mask = 16'hAAD8;
defparam \Mux20~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N13
dffeas \Reg[27][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][11] .is_wysiwyg = "true";
defparam \Reg[27][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N30
cycloneive_lcell_comb \Mux20~8 (
// Equation(s):
// \Mux20~8_combout  = (ifid_ifinstr_o_24 & ((\Mux20~7_combout  & (\Reg[31][11]~q )) # (!\Mux20~7_combout  & ((\Reg[27][11]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux20~7_combout ))))

	.dataa(\Reg[31][11]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Mux20~7_combout ),
	.datad(\Reg[27][11]~q ),
	.cin(gnd),
	.combout(\Mux20~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~8 .lut_mask = 16'hBCB0;
defparam \Mux20~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N13
dffeas \Reg[13][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][11] .is_wysiwyg = "true";
defparam \Reg[13][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N12
cycloneive_lcell_comb \Mux20~17 (
// Equation(s):
// \Mux20~17_combout  = (ifid_ifinstr_o_21 & (((\Reg[13][11]~q ) # (ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & (\Reg[12][11]~q  & ((!ifid_ifinstr_o_22))))

	.dataa(\Reg[12][11]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[13][11]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux20~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~17 .lut_mask = 16'hCCE2;
defparam \Mux20~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N30
cycloneive_lcell_comb \Reg[15][11]~feeder (
// Equation(s):
// \Reg[15][11]~feeder_combout  = \wdat~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat14),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[15][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[15][11]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[15][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y36_N31
dffeas \Reg[15][11] (
	.clk(!CLK),
	.d(\Reg[15][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][11] .is_wysiwyg = "true";
defparam \Reg[15][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N5
dffeas \Reg[14][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][11] .is_wysiwyg = "true";
defparam \Reg[14][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N4
cycloneive_lcell_comb \Mux20~18 (
// Equation(s):
// \Mux20~18_combout  = (\Mux20~17_combout  & ((\Reg[15][11]~q ) # ((!ifid_ifinstr_o_22)))) # (!\Mux20~17_combout  & (((\Reg[14][11]~q  & ifid_ifinstr_o_22))))

	.dataa(\Mux20~17_combout ),
	.datab(\Reg[15][11]~q ),
	.datac(\Reg[14][11]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux20~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~18 .lut_mask = 16'hD8AA;
defparam \Mux20~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N4
cycloneive_lcell_comb \Reg[9][11]~feeder (
// Equation(s):
// \Reg[9][11]~feeder_combout  = \wdat~31_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat14),
	.cin(gnd),
	.combout(\Reg[9][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[9][11]~feeder .lut_mask = 16'hFF00;
defparam \Reg[9][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y32_N5
dffeas \Reg[9][11] (
	.clk(!CLK),
	.d(\Reg[9][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][11] .is_wysiwyg = "true";
defparam \Reg[9][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y36_N21
dffeas \Reg[11][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][11] .is_wysiwyg = "true";
defparam \Reg[11][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N9
dffeas \Reg[10][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][11] .is_wysiwyg = "true";
defparam \Reg[10][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N8
cycloneive_lcell_comb \Mux20~10 (
// Equation(s):
// \Mux20~10_combout  = (ifid_ifinstr_o_22 & (((\Reg[10][11]~q ) # (ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & (\Reg[8][11]~q  & ((!ifid_ifinstr_o_21))))

	.dataa(\Reg[8][11]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[10][11]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux20~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~10 .lut_mask = 16'hCCE2;
defparam \Mux20~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N6
cycloneive_lcell_comb \Mux20~11 (
// Equation(s):
// \Mux20~11_combout  = (ifid_ifinstr_o_21 & ((\Mux20~10_combout  & ((\Reg[11][11]~q ))) # (!\Mux20~10_combout  & (\Reg[9][11]~q )))) # (!ifid_ifinstr_o_21 & (((\Mux20~10_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[9][11]~q ),
	.datac(\Reg[11][11]~q ),
	.datad(\Mux20~10_combout ),
	.cin(gnd),
	.combout(\Mux20~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~11 .lut_mask = 16'hF588;
defparam \Mux20~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y39_N15
dffeas \Reg[4][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][11] .is_wysiwyg = "true";
defparam \Reg[4][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y39_N17
dffeas \Reg[5][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][11] .is_wysiwyg = "true";
defparam \Reg[5][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N14
cycloneive_lcell_comb \Mux20~12 (
// Equation(s):
// \Mux20~12_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[5][11]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[4][11]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[4][11]~q ),
	.datad(\Reg[5][11]~q ),
	.cin(gnd),
	.combout(\Mux20~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~12 .lut_mask = 16'hDC98;
defparam \Mux20~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y39_N27
dffeas \Reg[7][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][11] .is_wysiwyg = "true";
defparam \Reg[7][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N29
dffeas \Reg[6][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][11] .is_wysiwyg = "true";
defparam \Reg[6][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N26
cycloneive_lcell_comb \Mux20~13 (
// Equation(s):
// \Mux20~13_combout  = (ifid_ifinstr_o_22 & ((\Mux20~12_combout  & (\Reg[7][11]~q )) # (!\Mux20~12_combout  & ((\Reg[6][11]~q ))))) # (!ifid_ifinstr_o_22 & (\Mux20~12_combout ))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Mux20~12_combout ),
	.datac(\Reg[7][11]~q ),
	.datad(\Reg[6][11]~q ),
	.cin(gnd),
	.combout(\Mux20~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~13 .lut_mask = 16'hE6C4;
defparam \Mux20~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N23
dffeas \Reg[2][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][11] .is_wysiwyg = "true";
defparam \Reg[2][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N15
dffeas \Reg[1][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][11] .is_wysiwyg = "true";
defparam \Reg[1][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N29
dffeas \Reg[3][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][11] .is_wysiwyg = "true";
defparam \Reg[3][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N28
cycloneive_lcell_comb \Mux20~14 (
// Equation(s):
// \Mux20~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][11]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][11]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[1][11]~q ),
	.datac(\Reg[3][11]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux20~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~14 .lut_mask = 16'hA088;
defparam \Mux20~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N4
cycloneive_lcell_comb \Mux20~15 (
// Equation(s):
// \Mux20~15_combout  = (\Mux20~14_combout ) # ((ifid_ifinstr_o_22 & (\Reg[2][11]~q  & !ifid_ifinstr_o_21)))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[2][11]~q ),
	.datac(\Mux20~14_combout ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux20~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~15 .lut_mask = 16'hF0F8;
defparam \Mux20~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N18
cycloneive_lcell_comb \Mux20~16 (
// Equation(s):
// \Mux20~16_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & (\Mux20~13_combout )) # (!ifid_ifinstr_o_23 & ((\Mux20~15_combout )))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux20~13_combout ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux20~15_combout ),
	.cin(gnd),
	.combout(\Mux20~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~16 .lut_mask = 16'hE5E0;
defparam \Mux20~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N30
cycloneive_lcell_comb \Reg[21][10]~feeder (
// Equation(s):
// \Reg[21][10]~feeder_combout  = \wdat~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat15),
	.cin(gnd),
	.combout(\Reg[21][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[21][10]~feeder .lut_mask = 16'hFF00;
defparam \Reg[21][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N31
dffeas \Reg[21][10] (
	.clk(!CLK),
	.d(\Reg[21][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][10] .is_wysiwyg = "true";
defparam \Reg[21][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N2
cycloneive_lcell_comb \Reg[29][10]~feeder (
// Equation(s):
// \Reg[29][10]~feeder_combout  = \wdat~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat15),
	.cin(gnd),
	.combout(\Reg[29][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[29][10]~feeder .lut_mask = 16'hFF00;
defparam \Reg[29][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y38_N3
dffeas \Reg[29][10] (
	.clk(!CLK),
	.d(\Reg[29][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][10] .is_wysiwyg = "true";
defparam \Reg[29][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N25
dffeas \Reg[17][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][10] .is_wysiwyg = "true";
defparam \Reg[17][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N24
cycloneive_lcell_comb \Reg[25][10]~feeder (
// Equation(s):
// \Reg[25][10]~feeder_combout  = \wdat~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat15),
	.cin(gnd),
	.combout(\Reg[25][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][10]~feeder .lut_mask = 16'hFF00;
defparam \Reg[25][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N25
dffeas \Reg[25][10] (
	.clk(!CLK),
	.d(\Reg[25][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][10] .is_wysiwyg = "true";
defparam \Reg[25][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N6
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// \Mux21~0_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23) # (\Reg[25][10]~q )))) # (!ifid_ifinstr_o_24 & (\Reg[17][10]~q  & (!ifid_ifinstr_o_23)))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[17][10]~q ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Reg[25][10]~q ),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hAEA4;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N8
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// \Mux21~1_combout  = (ifid_ifinstr_o_23 & ((\Mux21~0_combout  & ((\Reg[29][10]~q ))) # (!\Mux21~0_combout  & (\Reg[21][10]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux21~0_combout ))))

	.dataa(\Reg[21][10]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[29][10]~q ),
	.datad(\Mux21~0_combout ),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'hF388;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N1
dffeas \Reg[26][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][10] .is_wysiwyg = "true";
defparam \Reg[26][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y30_N31
dffeas \Reg[18][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][10] .is_wysiwyg = "true";
defparam \Reg[18][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y36_N25
dffeas \Reg[22][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][10] .is_wysiwyg = "true";
defparam \Reg[22][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N24
cycloneive_lcell_comb \Mux21~2 (
// Equation(s):
// \Mux21~2_combout  = (ifid_ifinstr_o_23 & (((\Reg[22][10]~q ) # (ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (\Reg[18][10]~q  & ((!ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[18][10]~q ),
	.datac(\Reg[22][10]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux21~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~2 .lut_mask = 16'hAAE4;
defparam \Mux21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N0
cycloneive_lcell_comb \Mux21~3 (
// Equation(s):
// \Mux21~3_combout  = (ifid_ifinstr_o_24 & ((\Mux21~2_combout  & (\Reg[30][10]~q )) # (!\Mux21~2_combout  & ((\Reg[26][10]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux21~2_combout ))))

	.dataa(\Reg[30][10]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[26][10]~q ),
	.datad(\Mux21~2_combout ),
	.cin(gnd),
	.combout(\Mux21~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~3 .lut_mask = 16'hBBC0;
defparam \Mux21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y34_N9
dffeas \Reg[20][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][10] .is_wysiwyg = "true";
defparam \Reg[20][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N6
cycloneive_lcell_comb \Reg[16][10]~feeder (
// Equation(s):
// \Reg[16][10]~feeder_combout  = \wdat~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat15),
	.cin(gnd),
	.combout(\Reg[16][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[16][10]~feeder .lut_mask = 16'hFF00;
defparam \Reg[16][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N7
dffeas \Reg[16][10] (
	.clk(!CLK),
	.d(\Reg[16][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][10] .is_wysiwyg = "true";
defparam \Reg[16][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N8
cycloneive_lcell_comb \Mux21~4 (
// Equation(s):
// \Mux21~4_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & (\Reg[20][10]~q )) # (!ifid_ifinstr_o_23 & ((\Reg[16][10]~q )))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[20][10]~q ),
	.datad(\Reg[16][10]~q ),
	.cin(gnd),
	.combout(\Mux21~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~4 .lut_mask = 16'hD9C8;
defparam \Mux21~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N7
dffeas \Reg[28][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][10] .is_wysiwyg = "true";
defparam \Reg[28][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N20
cycloneive_lcell_comb \Reg[24][10]~feeder (
// Equation(s):
// \Reg[24][10]~feeder_combout  = \wdat~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat15),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[24][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[24][10]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[24][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N21
dffeas \Reg[24][10] (
	.clk(!CLK),
	.d(\Reg[24][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][10] .is_wysiwyg = "true";
defparam \Reg[24][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N6
cycloneive_lcell_comb \Mux21~5 (
// Equation(s):
// \Mux21~5_combout  = (ifid_ifinstr_o_24 & ((\Mux21~4_combout  & (\Reg[28][10]~q )) # (!\Mux21~4_combout  & ((\Reg[24][10]~q ))))) # (!ifid_ifinstr_o_24 & (\Mux21~4_combout ))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux21~4_combout ),
	.datac(\Reg[28][10]~q ),
	.datad(\Reg[24][10]~q ),
	.cin(gnd),
	.combout(\Mux21~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~5 .lut_mask = 16'hE6C4;
defparam \Mux21~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N8
cycloneive_lcell_comb \Mux21~6 (
// Equation(s):
// \Mux21~6_combout  = (ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21) # ((\Mux21~3_combout )))) # (!ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & ((\Mux21~5_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux21~3_combout ),
	.datad(\Mux21~5_combout ),
	.cin(gnd),
	.combout(\Mux21~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~6 .lut_mask = 16'hB9A8;
defparam \Mux21~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N25
dffeas \Reg[27][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][10] .is_wysiwyg = "true";
defparam \Reg[27][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N11
dffeas \Reg[19][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][10] .is_wysiwyg = "true";
defparam \Reg[19][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N24
cycloneive_lcell_comb \Mux21~7 (
// Equation(s):
// \Mux21~7_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[27][10]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[19][10]~q )))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[27][10]~q ),
	.datad(\Reg[19][10]~q ),
	.cin(gnd),
	.combout(\Mux21~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~7 .lut_mask = 16'hD9C8;
defparam \Mux21~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N1
dffeas \Reg[23][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][10] .is_wysiwyg = "true";
defparam \Reg[23][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y29_N9
dffeas \Reg[31][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][10] .is_wysiwyg = "true";
defparam \Reg[31][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N0
cycloneive_lcell_comb \Mux21~8 (
// Equation(s):
// \Mux21~8_combout  = (ifid_ifinstr_o_23 & ((\Mux21~7_combout  & ((\Reg[31][10]~q ))) # (!\Mux21~7_combout  & (\Reg[23][10]~q )))) # (!ifid_ifinstr_o_23 & (\Mux21~7_combout ))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux21~7_combout ),
	.datac(\Reg[23][10]~q ),
	.datad(\Reg[31][10]~q ),
	.cin(gnd),
	.combout(\Mux21~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~8 .lut_mask = 16'hEC64;
defparam \Mux21~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y39_N11
dffeas \Reg[7][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][10] .is_wysiwyg = "true";
defparam \Reg[7][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y39_N5
dffeas \Reg[5][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][10] .is_wysiwyg = "true";
defparam \Reg[5][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y39_N31
dffeas \Reg[4][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][10] .is_wysiwyg = "true";
defparam \Reg[4][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N4
cycloneive_lcell_comb \Mux21~10 (
// Equation(s):
// \Mux21~10_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[5][10]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[4][10]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[5][10]~q ),
	.datad(\Reg[4][10]~q ),
	.cin(gnd),
	.combout(\Mux21~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~10 .lut_mask = 16'hD9C8;
defparam \Mux21~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y39_N13
dffeas \Reg[6][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][10] .is_wysiwyg = "true";
defparam \Reg[6][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N12
cycloneive_lcell_comb \Mux21~11 (
// Equation(s):
// \Mux21~11_combout  = (\Mux21~10_combout  & ((\Reg[7][10]~q ) # ((!ifid_ifinstr_o_22)))) # (!\Mux21~10_combout  & (((\Reg[6][10]~q  & ifid_ifinstr_o_22))))

	.dataa(\Reg[7][10]~q ),
	.datab(\Mux21~10_combout ),
	.datac(\Reg[6][10]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux21~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~11 .lut_mask = 16'hB8CC;
defparam \Mux21~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N1
dffeas \Reg[13][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][10] .is_wysiwyg = "true";
defparam \Reg[13][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N0
cycloneive_lcell_comb \Mux21~17 (
// Equation(s):
// \Mux21~17_combout  = (ifid_ifinstr_o_21 & (((\Reg[13][10]~q ) # (ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & (\Reg[12][10]~q  & ((!ifid_ifinstr_o_22))))

	.dataa(\Reg[12][10]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[13][10]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux21~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~17 .lut_mask = 16'hCCE2;
defparam \Mux21~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N11
dffeas \Reg[14][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][10] .is_wysiwyg = "true";
defparam \Reg[14][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N13
dffeas \Reg[15][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][10] .is_wysiwyg = "true";
defparam \Reg[15][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N10
cycloneive_lcell_comb \Mux21~18 (
// Equation(s):
// \Mux21~18_combout  = (\Mux21~17_combout  & (((\Reg[15][10]~q )) # (!ifid_ifinstr_o_22))) # (!\Mux21~17_combout  & (ifid_ifinstr_o_22 & (\Reg[14][10]~q )))

	.dataa(\Mux21~17_combout ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[14][10]~q ),
	.datad(\Reg[15][10]~q ),
	.cin(gnd),
	.combout(\Mux21~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~18 .lut_mask = 16'hEA62;
defparam \Mux21~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N11
dffeas \Reg[2][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][10] .is_wysiwyg = "true";
defparam \Reg[2][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N31
dffeas \Reg[3][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][10] .is_wysiwyg = "true";
defparam \Reg[3][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y36_N21
dffeas \Reg[1][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][10] .is_wysiwyg = "true";
defparam \Reg[1][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N30
cycloneive_lcell_comb \Mux21~14 (
// Equation(s):
// \Mux21~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[3][10]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[1][10]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[3][10]~q ),
	.datad(\Reg[1][10]~q ),
	.cin(gnd),
	.combout(\Mux21~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~14 .lut_mask = 16'hA280;
defparam \Mux21~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N4
cycloneive_lcell_comb \Mux21~15 (
// Equation(s):
// \Mux21~15_combout  = (\Mux21~14_combout ) # ((ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & \Reg[2][10]~q )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[2][10]~q ),
	.datad(\Mux21~14_combout ),
	.cin(gnd),
	.combout(\Mux21~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~15 .lut_mask = 16'hFF20;
defparam \Mux21~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y36_N1
dffeas \Reg[11][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][10] .is_wysiwyg = "true";
defparam \Reg[11][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N3
dffeas \Reg[8][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][10] .is_wysiwyg = "true";
defparam \Reg[8][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N17
dffeas \Reg[10][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][10] .is_wysiwyg = "true";
defparam \Reg[10][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N2
cycloneive_lcell_comb \Mux21~12 (
// Equation(s):
// \Mux21~12_combout  = (ifid_ifinstr_o_21 & (ifid_ifinstr_o_22)) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[10][10]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[8][10]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[8][10]~q ),
	.datad(\Reg[10][10]~q ),
	.cin(gnd),
	.combout(\Mux21~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~12 .lut_mask = 16'hDC98;
defparam \Mux21~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N0
cycloneive_lcell_comb \Mux21~13 (
// Equation(s):
// \Mux21~13_combout  = (ifid_ifinstr_o_21 & ((\Mux21~12_combout  & ((\Reg[11][10]~q ))) # (!\Mux21~12_combout  & (\Reg[9][10]~q )))) # (!ifid_ifinstr_o_21 & (((\Mux21~12_combout ))))

	.dataa(\Reg[9][10]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[11][10]~q ),
	.datad(\Mux21~12_combout ),
	.cin(gnd),
	.combout(\Mux21~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~13 .lut_mask = 16'hF388;
defparam \Mux21~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N18
cycloneive_lcell_comb \Mux21~16 (
// Equation(s):
// \Mux21~16_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Mux21~13_combout ))) # (!ifid_ifinstr_o_24 & (\Mux21~15_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux21~15_combout ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Mux21~13_combout ),
	.cin(gnd),
	.combout(\Mux21~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~16 .lut_mask = 16'hF4A4;
defparam \Mux21~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N29
dffeas \Reg[25][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][9] .is_wysiwyg = "true";
defparam \Reg[25][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y37_N11
dffeas \Reg[29][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][9] .is_wysiwyg = "true";
defparam \Reg[29][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y37_N9
dffeas \Reg[21][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][9] .is_wysiwyg = "true";
defparam \Reg[21][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N11
dffeas \Reg[17][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][9] .is_wysiwyg = "true";
defparam \Reg[17][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N10
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// \Mux22~0_combout  = (ifid_ifinstr_o_23 & ((\Reg[21][9]~q ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((\Reg[17][9]~q  & !ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[21][9]~q ),
	.datac(\Reg[17][9]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'hAAD8;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N10
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// \Mux22~1_combout  = (ifid_ifinstr_o_24 & ((\Mux22~0_combout  & ((\Reg[29][9]~q ))) # (!\Mux22~0_combout  & (\Reg[25][9]~q )))) # (!ifid_ifinstr_o_24 & (((\Mux22~0_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[25][9]~q ),
	.datac(\Reg[29][9]~q ),
	.datad(\Mux22~0_combout ),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'hF588;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N9
dffeas \Reg[30][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][9] .is_wysiwyg = "true";
defparam \Reg[30][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y33_N17
dffeas \Reg[18][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][9] .is_wysiwyg = "true";
defparam \Reg[18][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N18
cycloneive_lcell_comb \Reg[26][9]~feeder (
// Equation(s):
// \Reg[26][9]~feeder_combout  = \wdat~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat16),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[26][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[26][9]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[26][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N19
dffeas \Reg[26][9] (
	.clk(!CLK),
	.d(\Reg[26][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][9] .is_wysiwyg = "true";
defparam \Reg[26][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N16
cycloneive_lcell_comb \Mux22~2 (
// Equation(s):
// \Mux22~2_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[26][9]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & (\Reg[18][9]~q )))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[18][9]~q ),
	.datad(\Reg[26][9]~q ),
	.cin(gnd),
	.combout(\Mux22~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~2 .lut_mask = 16'hBA98;
defparam \Mux22~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N2
cycloneive_lcell_comb \Mux22~3 (
// Equation(s):
// \Mux22~3_combout  = (ifid_ifinstr_o_23 & ((\Mux22~2_combout  & ((\Reg[30][9]~q ))) # (!\Mux22~2_combout  & (\Reg[22][9]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux22~2_combout ))))

	.dataa(\Reg[22][9]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[30][9]~q ),
	.datad(\Mux22~2_combout ),
	.cin(gnd),
	.combout(\Mux22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~3 .lut_mask = 16'hF388;
defparam \Mux22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N14
cycloneive_lcell_comb \Reg[20][9]~feeder (
// Equation(s):
// \Reg[20][9]~feeder_combout  = \wdat~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat16),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[20][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[20][9]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[20][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N15
dffeas \Reg[20][9] (
	.clk(!CLK),
	.d(\Reg[20][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][9] .is_wysiwyg = "true";
defparam \Reg[20][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N13
dffeas \Reg[24][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][9] .is_wysiwyg = "true";
defparam \Reg[24][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N12
cycloneive_lcell_comb \Mux22~4 (
// Equation(s):
// \Mux22~4_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Reg[24][9]~q ))) # (!ifid_ifinstr_o_24 & (\Reg[16][9]~q ))))

	.dataa(\Reg[16][9]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[24][9]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux22~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~4 .lut_mask = 16'hFC22;
defparam \Mux22~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N0
cycloneive_lcell_comb \Mux22~5 (
// Equation(s):
// \Mux22~5_combout  = (ifid_ifinstr_o_23 & ((\Mux22~4_combout  & (\Reg[28][9]~q )) # (!\Mux22~4_combout  & ((\Reg[20][9]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux22~4_combout ))))

	.dataa(\Reg[28][9]~q ),
	.datab(\Reg[20][9]~q ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux22~4_combout ),
	.cin(gnd),
	.combout(\Mux22~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~5 .lut_mask = 16'hAFC0;
defparam \Mux22~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N14
cycloneive_lcell_comb \Mux22~6 (
// Equation(s):
// \Mux22~6_combout  = (ifid_ifinstr_o_21 & (ifid_ifinstr_o_22)) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Mux22~3_combout )) # (!ifid_ifinstr_o_22 & ((\Mux22~5_combout )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Mux22~3_combout ),
	.datad(\Mux22~5_combout ),
	.cin(gnd),
	.combout(\Mux22~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~6 .lut_mask = 16'hD9C8;
defparam \Mux22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N8
cycloneive_lcell_comb \Reg[31][9]~feeder (
// Equation(s):
// \Reg[31][9]~feeder_combout  = \wdat~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat16),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[31][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[31][9]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[31][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N9
dffeas \Reg[31][9] (
	.clk(!CLK),
	.d(\Reg[31][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][9] .is_wysiwyg = "true";
defparam \Reg[31][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N17
dffeas \Reg[27][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][9] .is_wysiwyg = "true";
defparam \Reg[27][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N23
dffeas \Reg[19][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][9] .is_wysiwyg = "true";
defparam \Reg[19][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N4
cycloneive_lcell_comb \Reg[23][9]~feeder (
// Equation(s):
// \Reg[23][9]~feeder_combout  = \wdat~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat16),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[23][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[23][9]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[23][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N5
dffeas \Reg[23][9] (
	.clk(!CLK),
	.d(\Reg[23][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][9] .is_wysiwyg = "true";
defparam \Reg[23][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N14
cycloneive_lcell_comb \Mux22~7 (
// Equation(s):
// \Mux22~7_combout  = (ifid_ifinstr_o_23 & (((\Reg[23][9]~q ) # (ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (\Reg[19][9]~q  & ((!ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[19][9]~q ),
	.datac(\Reg[23][9]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux22~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~7 .lut_mask = 16'hAAE4;
defparam \Mux22~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N16
cycloneive_lcell_comb \Mux22~8 (
// Equation(s):
// \Mux22~8_combout  = (ifid_ifinstr_o_24 & ((\Mux22~7_combout  & (\Reg[31][9]~q )) # (!\Mux22~7_combout  & ((\Reg[27][9]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux22~7_combout ))))

	.dataa(\Reg[31][9]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[27][9]~q ),
	.datad(\Mux22~7_combout ),
	.cin(gnd),
	.combout(\Mux22~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~8 .lut_mask = 16'hBBC0;
defparam \Mux22~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N3
dffeas \Reg[14][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][9] .is_wysiwyg = "true";
defparam \Reg[14][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N2
cycloneive_lcell_comb \Reg[15][9]~feeder (
// Equation(s):
// \Reg[15][9]~feeder_combout  = \wdat~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat16),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[15][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[15][9]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[15][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y28_N3
dffeas \Reg[15][9] (
	.clk(!CLK),
	.d(\Reg[15][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][9] .is_wysiwyg = "true";
defparam \Reg[15][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N21
dffeas \Reg[13][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][9] .is_wysiwyg = "true";
defparam \Reg[13][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N15
dffeas \Reg[12][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][9] .is_wysiwyg = "true";
defparam \Reg[12][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N14
cycloneive_lcell_comb \Mux22~17 (
// Equation(s):
// \Mux22~17_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[13][9]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[12][9]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[13][9]~q ),
	.datac(\Reg[12][9]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux22~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~17 .lut_mask = 16'hEE50;
defparam \Mux22~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N12
cycloneive_lcell_comb \Mux22~18 (
// Equation(s):
// \Mux22~18_combout  = (ifid_ifinstr_o_22 & ((\Mux22~17_combout  & ((\Reg[15][9]~q ))) # (!\Mux22~17_combout  & (\Reg[14][9]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux22~17_combout ))))

	.dataa(\Reg[14][9]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[15][9]~q ),
	.datad(\Mux22~17_combout ),
	.cin(gnd),
	.combout(\Mux22~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~18 .lut_mask = 16'hF388;
defparam \Mux22~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N7
dffeas \Reg[11][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][9] .is_wysiwyg = "true";
defparam \Reg[11][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N21
dffeas \Reg[10][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][9] .is_wysiwyg = "true";
defparam \Reg[10][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N11
dffeas \Reg[8][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][9] .is_wysiwyg = "true";
defparam \Reg[8][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N20
cycloneive_lcell_comb \Mux22~10 (
// Equation(s):
// \Mux22~10_combout  = (ifid_ifinstr_o_21 & (ifid_ifinstr_o_22)) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[10][9]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[8][9]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[10][9]~q ),
	.datad(\Reg[8][9]~q ),
	.cin(gnd),
	.combout(\Mux22~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~10 .lut_mask = 16'hD9C8;
defparam \Mux22~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N5
dffeas \Reg[9][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][9] .is_wysiwyg = "true";
defparam \Reg[9][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N4
cycloneive_lcell_comb \Mux22~11 (
// Equation(s):
// \Mux22~11_combout  = (\Mux22~10_combout  & ((\Reg[11][9]~q ) # ((!ifid_ifinstr_o_21)))) # (!\Mux22~10_combout  & (((\Reg[9][9]~q  & ifid_ifinstr_o_21))))

	.dataa(\Reg[11][9]~q ),
	.datab(\Mux22~10_combout ),
	.datac(\Reg[9][9]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux22~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~11 .lut_mask = 16'hB8CC;
defparam \Mux22~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y39_N5
dffeas \Reg[6][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][9] .is_wysiwyg = "true";
defparam \Reg[6][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N19
dffeas \Reg[7][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][9] .is_wysiwyg = "true";
defparam \Reg[7][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y39_N3
dffeas \Reg[4][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][9] .is_wysiwyg = "true";
defparam \Reg[4][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y39_N29
dffeas \Reg[5][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][9] .is_wysiwyg = "true";
defparam \Reg[5][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N2
cycloneive_lcell_comb \Mux22~12 (
// Equation(s):
// \Mux22~12_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[5][9]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[4][9]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[4][9]~q ),
	.datad(\Reg[5][9]~q ),
	.cin(gnd),
	.combout(\Mux22~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~12 .lut_mask = 16'hDC98;
defparam \Mux22~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N18
cycloneive_lcell_comb \Mux22~13 (
// Equation(s):
// \Mux22~13_combout  = (ifid_ifinstr_o_22 & ((\Mux22~12_combout  & ((\Reg[7][9]~q ))) # (!\Mux22~12_combout  & (\Reg[6][9]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux22~12_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[6][9]~q ),
	.datac(\Reg[7][9]~q ),
	.datad(\Mux22~12_combout ),
	.cin(gnd),
	.combout(\Mux22~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~13 .lut_mask = 16'hF588;
defparam \Mux22~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N4
cycloneive_lcell_comb \Reg[2][9]~feeder (
// Equation(s):
// \Reg[2][9]~feeder_combout  = \wdat~35_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat16),
	.cin(gnd),
	.combout(\Reg[2][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[2][9]~feeder .lut_mask = 16'hFF00;
defparam \Reg[2][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N5
dffeas \Reg[2][9] (
	.clk(!CLK),
	.d(\Reg[2][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][9] .is_wysiwyg = "true";
defparam \Reg[2][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N22
cycloneive_lcell_comb \Mux22~15 (
// Equation(s):
// \Mux22~15_combout  = (\Mux22~14_combout ) # ((!ifid_ifinstr_o_21 & (\Reg[2][9]~q  & ifid_ifinstr_o_22)))

	.dataa(\Mux22~14_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[2][9]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux22~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~15 .lut_mask = 16'hBAAA;
defparam \Mux22~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N10
cycloneive_lcell_comb \Mux22~16 (
// Equation(s):
// \Mux22~16_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & (\Mux22~13_combout )) # (!ifid_ifinstr_o_23 & ((\Mux22~15_combout )))))

	.dataa(\Mux22~13_combout ),
	.datab(ifid_ifinstr_o_24),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux22~15_combout ),
	.cin(gnd),
	.combout(\Mux22~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~16 .lut_mask = 16'hE3E0;
defparam \Mux22~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N16
cycloneive_lcell_comb \Mux59~0 (
// Equation(s):
// \Mux59~0_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19) # (\Reg[21][4]~q )))) # (!ifid_ifinstr_o_18 & (\Reg[17][4]~q  & (!ifid_ifinstr_o_19)))

	.dataa(\Reg[17][4]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(ifid_ifinstr_o_19),
	.datad(\Reg[21][4]~q ),
	.cin(gnd),
	.combout(\Mux59~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~0 .lut_mask = 16'hCEC2;
defparam \Mux59~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N2
cycloneive_lcell_comb \Mux59~1 (
// Equation(s):
// \Mux59~1_combout  = (ifid_ifinstr_o_19 & ((\Mux59~0_combout  & (\Reg[29][4]~q )) # (!\Mux59~0_combout  & ((\Reg[25][4]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux59~0_combout ))))

	.dataa(\Reg[29][4]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[25][4]~q ),
	.datad(\Mux59~0_combout ),
	.cin(gnd),
	.combout(\Mux59~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~1 .lut_mask = 16'hBBC0;
defparam \Mux59~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N18
cycloneive_lcell_comb \Mux59~7 (
// Equation(s):
// \Mux59~7_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Reg[23][4]~q ))) # (!ifid_ifinstr_o_18 & (\Reg[19][4]~q ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[19][4]~q ),
	.datad(\Reg[23][4]~q ),
	.cin(gnd),
	.combout(\Mux59~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~7 .lut_mask = 16'hDC98;
defparam \Mux59~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N10
cycloneive_lcell_comb \Mux59~8 (
// Equation(s):
// \Mux59~8_combout  = (\Mux59~7_combout  & (((\Reg[31][4]~q ) # (!ifid_ifinstr_o_19)))) # (!\Mux59~7_combout  & (\Reg[27][4]~q  & ((ifid_ifinstr_o_19))))

	.dataa(\Mux59~7_combout ),
	.datab(\Reg[27][4]~q ),
	.datac(\Reg[31][4]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux59~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~8 .lut_mask = 16'hE4AA;
defparam \Mux59~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N31
dffeas \Reg[26][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat3),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][4] .is_wysiwyg = "true";
defparam \Reg[26][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N30
cycloneive_lcell_comb \Reg[18][4]~feeder (
// Equation(s):
// \Reg[18][4]~feeder_combout  = \wdat~7_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat3),
	.cin(gnd),
	.combout(\Reg[18][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[18][4]~feeder .lut_mask = 16'hFF00;
defparam \Reg[18][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N31
dffeas \Reg[18][4] (
	.clk(!CLK),
	.d(\Reg[18][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][4] .is_wysiwyg = "true";
defparam \Reg[18][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N30
cycloneive_lcell_comb \Mux59~2 (
// Equation(s):
// \Mux59~2_combout  = (ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18) # ((\Reg[26][4]~q )))) # (!ifid_ifinstr_o_19 & (!ifid_ifinstr_o_18 & ((\Reg[18][4]~q ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[26][4]~q ),
	.datad(\Reg[18][4]~q ),
	.cin(gnd),
	.combout(\Mux59~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~2 .lut_mask = 16'hB9A8;
defparam \Mux59~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N22
cycloneive_lcell_comb \Mux59~3 (
// Equation(s):
// \Mux59~3_combout  = (ifid_ifinstr_o_18 & ((\Mux59~2_combout  & ((\Reg[30][4]~q ))) # (!\Mux59~2_combout  & (\Reg[22][4]~q )))) # (!ifid_ifinstr_o_18 & (((\Mux59~2_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[22][4]~q ),
	.datac(\Reg[30][4]~q ),
	.datad(\Mux59~2_combout ),
	.cin(gnd),
	.combout(\Mux59~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~3 .lut_mask = 16'hF588;
defparam \Mux59~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N6
cycloneive_lcell_comb \Mux59~4 (
// Equation(s):
// \Mux59~4_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[24][4]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[16][4]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[16][4]~q ),
	.datad(\Reg[24][4]~q ),
	.cin(gnd),
	.combout(\Mux59~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~4 .lut_mask = 16'hDC98;
defparam \Mux59~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N6
cycloneive_lcell_comb \Mux59~5 (
// Equation(s):
// \Mux59~5_combout  = (ifid_ifinstr_o_18 & ((\Mux59~4_combout  & ((\Reg[28][4]~q ))) # (!\Mux59~4_combout  & (\Reg[20][4]~q )))) # (!ifid_ifinstr_o_18 & (((\Mux59~4_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[20][4]~q ),
	.datac(\Reg[28][4]~q ),
	.datad(\Mux59~4_combout ),
	.cin(gnd),
	.combout(\Mux59~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~5 .lut_mask = 16'hF588;
defparam \Mux59~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N12
cycloneive_lcell_comb \Mux59~6 (
// Equation(s):
// \Mux59~6_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Mux59~3_combout )) # (!ifid_ifinstr_o_17 & ((\Mux59~5_combout )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux59~3_combout ),
	.datad(\Mux59~5_combout ),
	.cin(gnd),
	.combout(\Mux59~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~6 .lut_mask = 16'hD9C8;
defparam \Mux59~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N16
cycloneive_lcell_comb \Mux59~17 (
// Equation(s):
// \Mux59~17_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17) # ((\Reg[13][4]~q )))) # (!ifid_ifinstr_o_16 & (!ifid_ifinstr_o_17 & (\Reg[12][4]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[12][4]~q ),
	.datad(\Reg[13][4]~q ),
	.cin(gnd),
	.combout(\Mux59~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~17 .lut_mask = 16'hBA98;
defparam \Mux59~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N0
cycloneive_lcell_comb \Mux59~18 (
// Equation(s):
// \Mux59~18_combout  = (\Mux59~17_combout  & ((\Reg[15][4]~q ) # ((!ifid_ifinstr_o_17)))) # (!\Mux59~17_combout  & (((\Reg[14][4]~q  & ifid_ifinstr_o_17))))

	.dataa(\Reg[15][4]~q ),
	.datab(\Mux59~17_combout ),
	.datac(\Reg[14][4]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux59~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~18 .lut_mask = 16'hB8CC;
defparam \Mux59~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N2
cycloneive_lcell_comb \Mux59~15 (
// Equation(s):
// \Mux59~15_combout  = (\Mux59~14_combout ) # ((!ifid_ifinstr_o_16 & (\Reg[2][4]~q  & ifid_ifinstr_o_17)))

	.dataa(\Mux59~14_combout ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[2][4]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux59~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~15 .lut_mask = 16'hBAAA;
defparam \Mux59~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N20
cycloneive_lcell_comb \Mux59~13 (
// Equation(s):
// \Mux59~13_combout  = (\Mux59~12_combout  & (((\Reg[7][4]~q )) # (!ifid_ifinstr_o_17))) # (!\Mux59~12_combout  & (ifid_ifinstr_o_17 & ((\Reg[6][4]~q ))))

	.dataa(\Mux59~12_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[7][4]~q ),
	.datad(\Reg[6][4]~q ),
	.cin(gnd),
	.combout(\Mux59~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~13 .lut_mask = 16'hE6A2;
defparam \Mux59~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N4
cycloneive_lcell_comb \Mux59~16 (
// Equation(s):
// \Mux59~16_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19) # (\Mux59~13_combout )))) # (!ifid_ifinstr_o_18 & (\Mux59~15_combout  & (!ifid_ifinstr_o_19)))

	.dataa(\Mux59~15_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux59~13_combout ),
	.cin(gnd),
	.combout(\Mux59~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~16 .lut_mask = 16'hCEC2;
defparam \Mux59~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N8
cycloneive_lcell_comb \Mux59~10 (
// Equation(s):
// \Mux59~10_combout  = (ifid_ifinstr_o_17 & (((\Reg[10][4]~q ) # (ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & (\Reg[8][4]~q  & ((!ifid_ifinstr_o_16))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[8][4]~q ),
	.datac(\Reg[10][4]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux59~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~10 .lut_mask = 16'hAAE4;
defparam \Mux59~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N12
cycloneive_lcell_comb \Mux59~11 (
// Equation(s):
// \Mux59~11_combout  = (ifid_ifinstr_o_16 & ((\Mux59~10_combout  & ((\Reg[11][4]~q ))) # (!\Mux59~10_combout  & (\Reg[9][4]~q )))) # (!ifid_ifinstr_o_16 & (\Mux59~10_combout ))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux59~10_combout ),
	.datac(\Reg[9][4]~q ),
	.datad(\Reg[11][4]~q ),
	.cin(gnd),
	.combout(\Mux59~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~11 .lut_mask = 16'hEC64;
defparam \Mux59~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N18
cycloneive_lcell_comb \Reg[31][31]~feeder (
// Equation(s):
// \Reg[31][31]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat17),
	.cin(gnd),
	.combout(\Reg[31][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[31][31]~feeder .lut_mask = 16'hFF00;
defparam \Reg[31][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N19
dffeas \Reg[31][31] (
	.clk(!CLK),
	.d(\Reg[31][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][31] .is_wysiwyg = "true";
defparam \Reg[31][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N19
dffeas \Reg[27][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][31] .is_wysiwyg = "true";
defparam \Reg[27][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N5
dffeas \Reg[23][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][31] .is_wysiwyg = "true";
defparam \Reg[23][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N4
cycloneive_lcell_comb \Mux0~7 (
// Equation(s):
// \Mux0~7_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[23][31]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[19][31]~q ))))

	.dataa(\Reg[19][31]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[23][31]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~7 .lut_mask = 16'hFC22;
defparam \Mux0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N18
cycloneive_lcell_comb \Mux0~8 (
// Equation(s):
// \Mux0~8_combout  = (ifid_ifinstr_o_24 & ((\Mux0~7_combout  & (\Reg[31][31]~q )) # (!\Mux0~7_combout  & ((\Reg[27][31]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux0~7_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[31][31]~q ),
	.datac(\Reg[27][31]~q ),
	.datad(\Mux0~7_combout ),
	.cin(gnd),
	.combout(\Mux0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~8 .lut_mask = 16'hDDA0;
defparam \Mux0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N6
cycloneive_lcell_comb \Reg[25][31]~feeder (
// Equation(s):
// \Reg[25][31]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat17),
	.cin(gnd),
	.combout(\Reg[25][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][31]~feeder .lut_mask = 16'hFF00;
defparam \Reg[25][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N7
dffeas \Reg[25][31] (
	.clk(!CLK),
	.d(\Reg[25][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][31] .is_wysiwyg = "true";
defparam \Reg[25][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N13
dffeas \Reg[29][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][31] .is_wysiwyg = "true";
defparam \Reg[29][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N0
cycloneive_lcell_comb \Reg[17][31]~feeder (
// Equation(s):
// \Reg[17][31]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat17),
	.cin(gnd),
	.combout(\Reg[17][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[17][31]~feeder .lut_mask = 16'hFF00;
defparam \Reg[17][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N1
dffeas \Reg[17][31] (
	.clk(!CLK),
	.d(\Reg[17][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][31] .is_wysiwyg = "true";
defparam \Reg[17][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N7
dffeas \Reg[21][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][31] .is_wysiwyg = "true";
defparam \Reg[21][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N6
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// \Mux0~0_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[21][31]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[17][31]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[17][31]~q ),
	.datac(\Reg[21][31]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'hFA44;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N12
cycloneive_lcell_comb \Mux0~1 (
// Equation(s):
// \Mux0~1_combout  = (ifid_ifinstr_o_24 & ((\Mux0~0_combout  & ((\Reg[29][31]~q ))) # (!\Mux0~0_combout  & (\Reg[25][31]~q )))) # (!ifid_ifinstr_o_24 & (((\Mux0~0_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[25][31]~q ),
	.datac(\Reg[29][31]~q ),
	.datad(\Mux0~0_combout ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~1 .lut_mask = 16'hF588;
defparam \Mux0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N30
cycloneive_lcell_comb \Reg[22][31]~feeder (
// Equation(s):
// \Reg[22][31]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat17),
	.cin(gnd),
	.combout(\Reg[22][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[22][31]~feeder .lut_mask = 16'hFF00;
defparam \Reg[22][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y31_N31
dffeas \Reg[22][31] (
	.clk(!CLK),
	.d(\Reg[22][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][31] .is_wysiwyg = "true";
defparam \Reg[22][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N9
dffeas \Reg[26][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][31] .is_wysiwyg = "true";
defparam \Reg[26][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N3
dffeas \Reg[18][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][31] .is_wysiwyg = "true";
defparam \Reg[18][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N8
cycloneive_lcell_comb \Mux0~2 (
// Equation(s):
// \Mux0~2_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[26][31]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[18][31]~q )))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[26][31]~q ),
	.datad(\Reg[18][31]~q ),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~2 .lut_mask = 16'hD9C8;
defparam \Mux0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N8
cycloneive_lcell_comb \Mux0~3 (
// Equation(s):
// \Mux0~3_combout  = (ifid_ifinstr_o_23 & ((\Mux0~2_combout  & (\Reg[30][31]~q )) # (!\Mux0~2_combout  & ((\Reg[22][31]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux0~2_combout ))))

	.dataa(\Reg[30][31]~q ),
	.datab(\Reg[22][31]~q ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux0~2_combout ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~3 .lut_mask = 16'hAFC0;
defparam \Mux0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N12
cycloneive_lcell_comb \Reg[20][31]~feeder (
// Equation(s):
// \Reg[20][31]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat17),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[20][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[20][31]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[20][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y34_N13
dffeas \Reg[20][31] (
	.clk(!CLK),
	.d(\Reg[20][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][31] .is_wysiwyg = "true";
defparam \Reg[20][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N19
dffeas \Reg[28][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][31] .is_wysiwyg = "true";
defparam \Reg[28][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N28
cycloneive_lcell_comb \Mux0~5 (
// Equation(s):
// \Mux0~5_combout  = (\Mux0~4_combout  & (((\Reg[28][31]~q )) # (!ifid_ifinstr_o_23))) # (!\Mux0~4_combout  & (ifid_ifinstr_o_23 & (\Reg[20][31]~q )))

	.dataa(\Mux0~4_combout ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[20][31]~q ),
	.datad(\Reg[28][31]~q ),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~5 .lut_mask = 16'hEA62;
defparam \Mux0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N24
cycloneive_lcell_comb \Mux0~6 (
// Equation(s):
// \Mux0~6_combout  = (ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21) # ((\Mux0~3_combout )))) # (!ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & ((\Mux0~5_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux0~3_combout ),
	.datad(\Mux0~5_combout ),
	.cin(gnd),
	.combout(\Mux0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~6 .lut_mask = 16'hB9A8;
defparam \Mux0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N31
dffeas \Reg[15][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][31] .is_wysiwyg = "true";
defparam \Reg[15][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N5
dffeas \Reg[12][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][31] .is_wysiwyg = "true";
defparam \Reg[12][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N7
dffeas \Reg[13][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][31] .is_wysiwyg = "true";
defparam \Reg[13][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N6
cycloneive_lcell_comb \Mux0~17 (
// Equation(s):
// \Mux0~17_combout  = (ifid_ifinstr_o_21 & (((\Reg[13][31]~q ) # (ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & (\Reg[12][31]~q  & ((!ifid_ifinstr_o_22))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[12][31]~q ),
	.datac(\Reg[13][31]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~17 .lut_mask = 16'hAAE4;
defparam \Mux0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N9
dffeas \Reg[14][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][31] .is_wysiwyg = "true";
defparam \Reg[14][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N8
cycloneive_lcell_comb \Mux0~18 (
// Equation(s):
// \Mux0~18_combout  = (\Mux0~17_combout  & ((\Reg[15][31]~q ) # ((!ifid_ifinstr_o_22)))) # (!\Mux0~17_combout  & (((\Reg[14][31]~q  & ifid_ifinstr_o_22))))

	.dataa(\Reg[15][31]~q ),
	.datab(\Mux0~17_combout ),
	.datac(\Reg[14][31]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~18 .lut_mask = 16'hB8CC;
defparam \Mux0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N11
dffeas \Reg[11][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][31] .is_wysiwyg = "true";
defparam \Reg[11][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y33_N29
dffeas \Reg[9][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][31] .is_wysiwyg = "true";
defparam \Reg[9][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N29
dffeas \Reg[10][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][31] .is_wysiwyg = "true";
defparam \Reg[10][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N28
cycloneive_lcell_comb \Mux0~10 (
// Equation(s):
// \Mux0~10_combout  = (ifid_ifinstr_o_22 & (((\Reg[10][31]~q ) # (ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & (\Reg[8][31]~q  & ((!ifid_ifinstr_o_21))))

	.dataa(\Reg[8][31]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[10][31]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~10 .lut_mask = 16'hCCE2;
defparam \Mux0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N28
cycloneive_lcell_comb \Mux0~11 (
// Equation(s):
// \Mux0~11_combout  = (ifid_ifinstr_o_21 & ((\Mux0~10_combout  & (\Reg[11][31]~q )) # (!\Mux0~10_combout  & ((\Reg[9][31]~q ))))) # (!ifid_ifinstr_o_21 & (((\Mux0~10_combout ))))

	.dataa(\Reg[11][31]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[9][31]~q ),
	.datad(\Mux0~10_combout ),
	.cin(gnd),
	.combout(\Mux0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~11 .lut_mask = 16'hBBC0;
defparam \Mux0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N0
cycloneive_lcell_comb \Reg[2][31]~feeder (
// Equation(s):
// \Reg[2][31]~feeder_combout  = \wdat~37_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat17),
	.cin(gnd),
	.combout(\Reg[2][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[2][31]~feeder .lut_mask = 16'hFF00;
defparam \Reg[2][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N1
dffeas \Reg[2][31] (
	.clk(!CLK),
	.d(\Reg[2][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][31] .is_wysiwyg = "true";
defparam \Reg[2][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N9
dffeas \Reg[3][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][31] .is_wysiwyg = "true";
defparam \Reg[3][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N7
dffeas \Reg[1][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][31] .is_wysiwyg = "true";
defparam \Reg[1][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N8
cycloneive_lcell_comb \Mux0~14 (
// Equation(s):
// \Mux0~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[3][31]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[1][31]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[3][31]~q ),
	.datad(\Reg[1][31]~q ),
	.cin(gnd),
	.combout(\Mux0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~14 .lut_mask = 16'hA280;
defparam \Mux0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N18
cycloneive_lcell_comb \Mux0~15 (
// Equation(s):
// \Mux0~15_combout  = (\Mux0~14_combout ) # ((!ifid_ifinstr_o_21 & (\Reg[2][31]~q  & ifid_ifinstr_o_22)))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[2][31]~q ),
	.datac(ifid_ifinstr_o_22),
	.datad(\Mux0~14_combout ),
	.cin(gnd),
	.combout(\Mux0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~15 .lut_mask = 16'hFF40;
defparam \Mux0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y39_N25
dffeas \Reg[6][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][31] .is_wysiwyg = "true";
defparam \Reg[6][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N23
dffeas \Reg[7][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][31] .is_wysiwyg = "true";
defparam \Reg[7][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N7
dffeas \Reg[4][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][31] .is_wysiwyg = "true";
defparam \Reg[4][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N1
dffeas \Reg[5][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][31] .is_wysiwyg = "true";
defparam \Reg[5][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N6
cycloneive_lcell_comb \Mux0~12 (
// Equation(s):
// \Mux0~12_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22) # ((\Reg[5][31]~q )))) # (!ifid_ifinstr_o_21 & (!ifid_ifinstr_o_22 & (\Reg[4][31]~q )))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[4][31]~q ),
	.datad(\Reg[5][31]~q ),
	.cin(gnd),
	.combout(\Mux0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~12 .lut_mask = 16'hBA98;
defparam \Mux0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N22
cycloneive_lcell_comb \Mux0~13 (
// Equation(s):
// \Mux0~13_combout  = (ifid_ifinstr_o_22 & ((\Mux0~12_combout  & ((\Reg[7][31]~q ))) # (!\Mux0~12_combout  & (\Reg[6][31]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux0~12_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[6][31]~q ),
	.datac(\Reg[7][31]~q ),
	.datad(\Mux0~12_combout ),
	.cin(gnd),
	.combout(\Mux0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~13 .lut_mask = 16'hF588;
defparam \Mux0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N28
cycloneive_lcell_comb \Mux0~16 (
// Equation(s):
// \Mux0~16_combout  = (ifid_ifinstr_o_23 & (((\Mux0~13_combout ) # (ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (\Mux0~15_combout  & ((!ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Mux0~15_combout ),
	.datac(\Mux0~13_combout ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~16 .lut_mask = 16'hAAE4;
defparam \Mux0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N22
cycloneive_lcell_comb \Reg[29][29]~feeder (
// Equation(s):
// \Reg[29][29]~feeder_combout  = \wdat~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat18),
	.cin(gnd),
	.combout(\Reg[29][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[29][29]~feeder .lut_mask = 16'hFF00;
defparam \Reg[29][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y38_N23
dffeas \Reg[29][29] (
	.clk(!CLK),
	.d(\Reg[29][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][29] .is_wysiwyg = "true";
defparam \Reg[29][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N28
cycloneive_lcell_comb \Reg[25][29]~feeder (
// Equation(s):
// \Reg[25][29]~feeder_combout  = \wdat~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat18),
	.cin(gnd),
	.combout(\Reg[25][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][29]~feeder .lut_mask = 16'hFF00;
defparam \Reg[25][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y38_N29
dffeas \Reg[25][29] (
	.clk(!CLK),
	.d(\Reg[25][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][29] .is_wysiwyg = "true";
defparam \Reg[25][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N2
cycloneive_lcell_comb \Reg[21][29]~feeder (
// Equation(s):
// \Reg[21][29]~feeder_combout  = \wdat~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat18),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[21][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[21][29]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[21][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N3
dffeas \Reg[21][29] (
	.clk(!CLK),
	.d(\Reg[21][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][29] .is_wysiwyg = "true";
defparam \Reg[21][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N1
dffeas \Reg[17][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][29] .is_wysiwyg = "true";
defparam \Reg[17][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N4
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// \Mux2~0_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & (\Reg[21][29]~q )) # (!ifid_ifinstr_o_23 & ((\Reg[17][29]~q )))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[21][29]~q ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Reg[17][29]~q ),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'hE5E0;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N4
cycloneive_lcell_comb \Mux2~1 (
// Equation(s):
// \Mux2~1_combout  = (\Mux2~0_combout  & ((\Reg[29][29]~q ) # ((!ifid_ifinstr_o_24)))) # (!\Mux2~0_combout  & (((\Reg[25][29]~q  & ifid_ifinstr_o_24))))

	.dataa(\Reg[29][29]~q ),
	.datab(\Reg[25][29]~q ),
	.datac(\Mux2~0_combout ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~1 .lut_mask = 16'hACF0;
defparam \Mux2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N10
cycloneive_lcell_comb \Reg[23][29]~feeder (
// Equation(s):
// \Reg[23][29]~feeder_combout  = \wdat~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat18),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[23][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[23][29]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[23][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N11
dffeas \Reg[23][29] (
	.clk(!CLK),
	.d(\Reg[23][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][29] .is_wysiwyg = "true";
defparam \Reg[23][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N29
dffeas \Reg[19][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][29] .is_wysiwyg = "true";
defparam \Reg[19][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N28
cycloneive_lcell_comb \Mux2~7 (
// Equation(s):
// \Mux2~7_combout  = (ifid_ifinstr_o_23 & ((\Reg[23][29]~q ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((\Reg[19][29]~q  & !ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[23][29]~q ),
	.datac(\Reg[19][29]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~7 .lut_mask = 16'hAAD8;
defparam \Mux2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N11
dffeas \Reg[31][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][29] .is_wysiwyg = "true";
defparam \Reg[31][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N5
dffeas \Reg[27][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][29] .is_wysiwyg = "true";
defparam \Reg[27][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N18
cycloneive_lcell_comb \Mux2~8 (
// Equation(s):
// \Mux2~8_combout  = (\Mux2~7_combout  & ((\Reg[31][29]~q ) # ((!ifid_ifinstr_o_24)))) # (!\Mux2~7_combout  & (((ifid_ifinstr_o_24 & \Reg[27][29]~q ))))

	.dataa(\Mux2~7_combout ),
	.datab(\Reg[31][29]~q ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Reg[27][29]~q ),
	.cin(gnd),
	.combout(\Mux2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~8 .lut_mask = 16'hDA8A;
defparam \Mux2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N25
dffeas \Reg[22][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][29] .is_wysiwyg = "true";
defparam \Reg[22][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N19
dffeas \Reg[30][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][29] .is_wysiwyg = "true";
defparam \Reg[30][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y33_N27
dffeas \Reg[18][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][29] .is_wysiwyg = "true";
defparam \Reg[18][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N13
dffeas \Reg[26][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][29] .is_wysiwyg = "true";
defparam \Reg[26][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N26
cycloneive_lcell_comb \Mux2~2 (
// Equation(s):
// \Mux2~2_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[26][29]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & (\Reg[18][29]~q )))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[18][29]~q ),
	.datad(\Reg[26][29]~q ),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~2 .lut_mask = 16'hBA98;
defparam \Mux2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N22
cycloneive_lcell_comb \Mux2~3 (
// Equation(s):
// \Mux2~3_combout  = (ifid_ifinstr_o_23 & ((\Mux2~2_combout  & ((\Reg[30][29]~q ))) # (!\Mux2~2_combout  & (\Reg[22][29]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux2~2_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[22][29]~q ),
	.datac(\Reg[30][29]~q ),
	.datad(\Mux2~2_combout ),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~3 .lut_mask = 16'hF588;
defparam \Mux2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N19
dffeas \Reg[28][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][29] .is_wysiwyg = "true";
defparam \Reg[28][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N25
dffeas \Reg[24][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][29] .is_wysiwyg = "true";
defparam \Reg[24][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N24
cycloneive_lcell_comb \Mux2~4 (
// Equation(s):
// \Mux2~4_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Reg[24][29]~q ))) # (!ifid_ifinstr_o_24 & (\Reg[16][29]~q ))))

	.dataa(\Reg[16][29]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[24][29]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~4 .lut_mask = 16'hFC22;
defparam \Mux2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N18
cycloneive_lcell_comb \Mux2~5 (
// Equation(s):
// \Mux2~5_combout  = (ifid_ifinstr_o_23 & ((\Mux2~4_combout  & ((\Reg[28][29]~q ))) # (!\Mux2~4_combout  & (\Reg[20][29]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux2~4_combout ))))

	.dataa(\Reg[20][29]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[28][29]~q ),
	.datad(\Mux2~4_combout ),
	.cin(gnd),
	.combout(\Mux2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~5 .lut_mask = 16'hF388;
defparam \Mux2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N16
cycloneive_lcell_comb \Mux2~6 (
// Equation(s):
// \Mux2~6_combout  = (ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21) # ((\Mux2~3_combout )))) # (!ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & ((\Mux2~5_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux2~3_combout ),
	.datad(\Mux2~5_combout ),
	.cin(gnd),
	.combout(\Mux2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~6 .lut_mask = 16'hB9A8;
defparam \Mux2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N15
dffeas \Reg[2][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][29] .is_wysiwyg = "true";
defparam \Reg[2][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N9
dffeas \Reg[3][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][29] .is_wysiwyg = "true";
defparam \Reg[3][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N8
cycloneive_lcell_comb \Mux2~14 (
// Equation(s):
// \Mux2~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][29]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][29]~q ))))

	.dataa(\Reg[1][29]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[3][29]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux2~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~14 .lut_mask = 16'hC088;
defparam \Mux2~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N28
cycloneive_lcell_comb \Mux2~15 (
// Equation(s):
// \Mux2~15_combout  = (\Mux2~14_combout ) # ((!ifid_ifinstr_o_21 & (\Reg[2][29]~q  & ifid_ifinstr_o_22)))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[2][29]~q ),
	.datac(\Mux2~14_combout ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux2~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~15 .lut_mask = 16'hF4F0;
defparam \Mux2~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N31
dffeas \Reg[4][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][29] .is_wysiwyg = "true";
defparam \Reg[4][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N1
dffeas \Reg[5][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][29] .is_wysiwyg = "true";
defparam \Reg[5][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N30
cycloneive_lcell_comb \Mux2~12 (
// Equation(s):
// \Mux2~12_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[5][29]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[4][29]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[4][29]~q ),
	.datad(\Reg[5][29]~q ),
	.cin(gnd),
	.combout(\Mux2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~12 .lut_mask = 16'hDC98;
defparam \Mux2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N23
dffeas \Reg[6][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][29] .is_wysiwyg = "true";
defparam \Reg[6][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N28
cycloneive_lcell_comb \Reg[7][29]~feeder (
// Equation(s):
// \Reg[7][29]~feeder_combout  = \wdat~39_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat18),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[7][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[7][29]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[7][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N29
dffeas \Reg[7][29] (
	.clk(!CLK),
	.d(\Reg[7][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][29] .is_wysiwyg = "true";
defparam \Reg[7][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N22
cycloneive_lcell_comb \Mux2~13 (
// Equation(s):
// \Mux2~13_combout  = (ifid_ifinstr_o_22 & ((\Mux2~12_combout  & ((\Reg[7][29]~q ))) # (!\Mux2~12_combout  & (\Reg[6][29]~q )))) # (!ifid_ifinstr_o_22 & (\Mux2~12_combout ))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Mux2~12_combout ),
	.datac(\Reg[6][29]~q ),
	.datad(\Reg[7][29]~q ),
	.cin(gnd),
	.combout(\Mux2~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~13 .lut_mask = 16'hEC64;
defparam \Mux2~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N12
cycloneive_lcell_comb \Mux2~16 (
// Equation(s):
// \Mux2~16_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Mux2~13_combout ))) # (!ifid_ifinstr_o_23 & (\Mux2~15_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux2~15_combout ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux2~13_combout ),
	.cin(gnd),
	.combout(\Mux2~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~16 .lut_mask = 16'hF4A4;
defparam \Mux2~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N23
dffeas \Reg[15][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][29] .is_wysiwyg = "true";
defparam \Reg[15][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N29
dffeas \Reg[14][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][29] .is_wysiwyg = "true";
defparam \Reg[14][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N3
dffeas \Reg[12][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][29] .is_wysiwyg = "true";
defparam \Reg[12][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N9
dffeas \Reg[13][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][29] .is_wysiwyg = "true";
defparam \Reg[13][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N8
cycloneive_lcell_comb \Mux2~17 (
// Equation(s):
// \Mux2~17_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[13][29]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[12][29]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[12][29]~q ),
	.datac(\Reg[13][29]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux2~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~17 .lut_mask = 16'hFA44;
defparam \Mux2~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N28
cycloneive_lcell_comb \Mux2~18 (
// Equation(s):
// \Mux2~18_combout  = (ifid_ifinstr_o_22 & ((\Mux2~17_combout  & (\Reg[15][29]~q )) # (!\Mux2~17_combout  & ((\Reg[14][29]~q ))))) # (!ifid_ifinstr_o_22 & (((\Mux2~17_combout ))))

	.dataa(\Reg[15][29]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[14][29]~q ),
	.datad(\Mux2~17_combout ),
	.cin(gnd),
	.combout(\Mux2~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~18 .lut_mask = 16'hBBC0;
defparam \Mux2~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N23
dffeas \Reg[11][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][29] .is_wysiwyg = "true";
defparam \Reg[11][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y33_N9
dffeas \Reg[9][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][29] .is_wysiwyg = "true";
defparam \Reg[9][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N9
dffeas \Reg[10][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][29] .is_wysiwyg = "true";
defparam \Reg[10][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N3
dffeas \Reg[8][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][29] .is_wysiwyg = "true";
defparam \Reg[8][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N8
cycloneive_lcell_comb \Mux2~10 (
// Equation(s):
// \Mux2~10_combout  = (ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21) # ((\Reg[10][29]~q )))) # (!ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & ((\Reg[8][29]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[10][29]~q ),
	.datad(\Reg[8][29]~q ),
	.cin(gnd),
	.combout(\Mux2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~10 .lut_mask = 16'hB9A8;
defparam \Mux2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N8
cycloneive_lcell_comb \Mux2~11 (
// Equation(s):
// \Mux2~11_combout  = (ifid_ifinstr_o_21 & ((\Mux2~10_combout  & (\Reg[11][29]~q )) # (!\Mux2~10_combout  & ((\Reg[9][29]~q ))))) # (!ifid_ifinstr_o_21 & (((\Mux2~10_combout ))))

	.dataa(\Reg[11][29]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[9][29]~q ),
	.datad(\Mux2~10_combout ),
	.cin(gnd),
	.combout(\Mux2~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~11 .lut_mask = 16'hBBC0;
defparam \Mux2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N5
dffeas \Reg[21][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][30] .is_wysiwyg = "true";
defparam \Reg[21][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N21
dffeas \Reg[29][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][30] .is_wysiwyg = "true";
defparam \Reg[29][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N15
dffeas \Reg[25][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][30] .is_wysiwyg = "true";
defparam \Reg[25][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N7
dffeas \Reg[17][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][30] .is_wysiwyg = "true";
defparam \Reg[17][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N6
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// \Mux1~0_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[25][30]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[17][30]~q )))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[25][30]~q ),
	.datac(\Reg[17][30]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'hEE50;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N20
cycloneive_lcell_comb \Mux1~1 (
// Equation(s):
// \Mux1~1_combout  = (ifid_ifinstr_o_23 & ((\Mux1~0_combout  & ((\Reg[29][30]~q ))) # (!\Mux1~0_combout  & (\Reg[21][30]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux1~0_combout ))))

	.dataa(\Reg[21][30]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[29][30]~q ),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~1 .lut_mask = 16'hF388;
defparam \Mux1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N17
dffeas \Reg[24][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][30] .is_wysiwyg = "true";
defparam \Reg[24][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y34_N3
dffeas \Reg[28][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][30] .is_wysiwyg = "true";
defparam \Reg[28][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N0
cycloneive_lcell_comb \Reg[16][30]~feeder (
// Equation(s):
// \Reg[16][30]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat19),
	.cin(gnd),
	.combout(\Reg[16][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[16][30]~feeder .lut_mask = 16'hFF00;
defparam \Reg[16][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N1
dffeas \Reg[16][30] (
	.clk(!CLK),
	.d(\Reg[16][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][30] .is_wysiwyg = "true";
defparam \Reg[16][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y34_N21
dffeas \Reg[20][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][30] .is_wysiwyg = "true";
defparam \Reg[20][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N20
cycloneive_lcell_comb \Mux1~4 (
// Equation(s):
// \Mux1~4_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[20][30]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[16][30]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[16][30]~q ),
	.datac(\Reg[20][30]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~4 .lut_mask = 16'hFA44;
defparam \Mux1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N2
cycloneive_lcell_comb \Mux1~5 (
// Equation(s):
// \Mux1~5_combout  = (ifid_ifinstr_o_24 & ((\Mux1~4_combout  & ((\Reg[28][30]~q ))) # (!\Mux1~4_combout  & (\Reg[24][30]~q )))) # (!ifid_ifinstr_o_24 & (((\Mux1~4_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[24][30]~q ),
	.datac(\Reg[28][30]~q ),
	.datad(\Mux1~4_combout ),
	.cin(gnd),
	.combout(\Mux1~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~5 .lut_mask = 16'hF588;
defparam \Mux1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y36_N1
dffeas \Reg[22][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][30] .is_wysiwyg = "true";
defparam \Reg[22][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y30_N17
dffeas \Reg[18][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][30] .is_wysiwyg = "true";
defparam \Reg[18][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N0
cycloneive_lcell_comb \Mux1~2 (
// Equation(s):
// \Mux1~2_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & (\Reg[22][30]~q )) # (!ifid_ifinstr_o_23 & ((\Reg[18][30]~q )))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[22][30]~q ),
	.datad(\Reg[18][30]~q ),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~2 .lut_mask = 16'hD9C8;
defparam \Mux1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y36_N31
dffeas \Reg[30][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][30] .is_wysiwyg = "true";
defparam \Reg[30][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N8
cycloneive_lcell_comb \Reg[26][30]~feeder (
// Equation(s):
// \Reg[26][30]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat19),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[26][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[26][30]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[26][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y36_N9
dffeas \Reg[26][30] (
	.clk(!CLK),
	.d(\Reg[26][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][30] .is_wysiwyg = "true";
defparam \Reg[26][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N16
cycloneive_lcell_comb \Mux1~3 (
// Equation(s):
// \Mux1~3_combout  = (ifid_ifinstr_o_24 & ((\Mux1~2_combout  & (\Reg[30][30]~q )) # (!\Mux1~2_combout  & ((\Reg[26][30]~q ))))) # (!ifid_ifinstr_o_24 & (\Mux1~2_combout ))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux1~2_combout ),
	.datac(\Reg[30][30]~q ),
	.datad(\Reg[26][30]~q ),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~3 .lut_mask = 16'hE6C4;
defparam \Mux1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N22
cycloneive_lcell_comb \Mux1~6 (
// Equation(s):
// \Mux1~6_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Mux1~3_combout ))) # (!ifid_ifinstr_o_22 & (\Mux1~5_combout ))))

	.dataa(\Mux1~5_combout ),
	.datab(\Mux1~3_combout ),
	.datac(ifid_ifinstr_o_21),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux1~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~6 .lut_mask = 16'hFC0A;
defparam \Mux1~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N31
dffeas \Reg[31][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][30] .is_wysiwyg = "true";
defparam \Reg[31][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N9
dffeas \Reg[23][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][30] .is_wysiwyg = "true";
defparam \Reg[23][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N15
dffeas \Reg[19][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][30] .is_wysiwyg = "true";
defparam \Reg[19][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N14
cycloneive_lcell_comb \Mux1~7 (
// Equation(s):
// \Mux1~7_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[27][30]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[19][30]~q )))))

	.dataa(\Reg[27][30]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[19][30]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux1~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~7 .lut_mask = 16'hEE30;
defparam \Mux1~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N28
cycloneive_lcell_comb \Mux1~8 (
// Equation(s):
// \Mux1~8_combout  = (ifid_ifinstr_o_23 & ((\Mux1~7_combout  & (\Reg[31][30]~q )) # (!\Mux1~7_combout  & ((\Reg[23][30]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux1~7_combout ))))

	.dataa(\Reg[31][30]~q ),
	.datab(\Reg[23][30]~q ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux1~7_combout ),
	.cin(gnd),
	.combout(\Mux1~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~8 .lut_mask = 16'hAFC0;
defparam \Mux1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N12
cycloneive_lcell_comb \Reg[6][30]~feeder (
// Equation(s):
// \Reg[6][30]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat19),
	.cin(gnd),
	.combout(\Reg[6][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[6][30]~feeder .lut_mask = 16'hFF00;
defparam \Reg[6][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N13
dffeas \Reg[6][30] (
	.clk(!CLK),
	.d(\Reg[6][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][30] .is_wysiwyg = "true";
defparam \Reg[6][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y39_N21
dffeas \Reg[5][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][30] .is_wysiwyg = "true";
defparam \Reg[5][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y39_N27
dffeas \Reg[4][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][30] .is_wysiwyg = "true";
defparam \Reg[4][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N20
cycloneive_lcell_comb \Mux1~10 (
// Equation(s):
// \Mux1~10_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[5][30]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[4][30]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[5][30]~q ),
	.datad(\Reg[4][30]~q ),
	.cin(gnd),
	.combout(\Mux1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~10 .lut_mask = 16'hD9C8;
defparam \Mux1~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N17
dffeas \Reg[7][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][30] .is_wysiwyg = "true";
defparam \Reg[7][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N10
cycloneive_lcell_comb \Mux1~11 (
// Equation(s):
// \Mux1~11_combout  = (ifid_ifinstr_o_22 & ((\Mux1~10_combout  & ((\Reg[7][30]~q ))) # (!\Mux1~10_combout  & (\Reg[6][30]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux1~10_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[6][30]~q ),
	.datac(\Mux1~10_combout ),
	.datad(\Reg[7][30]~q ),
	.cin(gnd),
	.combout(\Mux1~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~11 .lut_mask = 16'hF858;
defparam \Mux1~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N27
dffeas \Reg[15][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][30] .is_wysiwyg = "true";
defparam \Reg[15][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N20
cycloneive_lcell_comb \Reg[13][30]~feeder (
// Equation(s):
// \Reg[13][30]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat19),
	.cin(gnd),
	.combout(\Reg[13][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[13][30]~feeder .lut_mask = 16'hFF00;
defparam \Reg[13][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N21
dffeas \Reg[13][30] (
	.clk(!CLK),
	.d(\Reg[13][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][30] .is_wysiwyg = "true";
defparam \Reg[13][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N29
dffeas \Reg[12][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][30] .is_wysiwyg = "true";
defparam \Reg[12][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N28
cycloneive_lcell_comb \Mux1~17 (
// Equation(s):
// \Mux1~17_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[13][30]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[12][30]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[13][30]~q ),
	.datac(\Reg[12][30]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux1~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~17 .lut_mask = 16'hEE50;
defparam \Mux1~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N17
dffeas \Reg[14][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][30] .is_wysiwyg = "true";
defparam \Reg[14][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N16
cycloneive_lcell_comb \Mux1~18 (
// Equation(s):
// \Mux1~18_combout  = (\Mux1~17_combout  & ((\Reg[15][30]~q ) # ((!ifid_ifinstr_o_22)))) # (!\Mux1~17_combout  & (((\Reg[14][30]~q  & ifid_ifinstr_o_22))))

	.dataa(\Reg[15][30]~q ),
	.datab(\Mux1~17_combout ),
	.datac(\Reg[14][30]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux1~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~18 .lut_mask = 16'hB8CC;
defparam \Mux1~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N7
dffeas \Reg[2][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][30] .is_wysiwyg = "true";
defparam \Reg[2][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N6
cycloneive_lcell_comb \Mux1~15 (
// Equation(s):
// \Mux1~15_combout  = (\Mux1~14_combout ) # ((!ifid_ifinstr_o_21 & (\Reg[2][30]~q  & ifid_ifinstr_o_22)))

	.dataa(\Mux1~14_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[2][30]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux1~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~15 .lut_mask = 16'hBAAA;
defparam \Mux1~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N3
dffeas \Reg[11][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][30] .is_wysiwyg = "true";
defparam \Reg[11][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y33_N21
dffeas \Reg[9][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][30] .is_wysiwyg = "true";
defparam \Reg[9][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N2
cycloneive_lcell_comb \Mux1~13 (
// Equation(s):
// \Mux1~13_combout  = (\Mux1~12_combout  & (((\Reg[11][30]~q )) # (!ifid_ifinstr_o_21))) # (!\Mux1~12_combout  & (ifid_ifinstr_o_21 & ((\Reg[9][30]~q ))))

	.dataa(\Mux1~12_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[11][30]~q ),
	.datad(\Reg[9][30]~q ),
	.cin(gnd),
	.combout(\Mux1~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~13 .lut_mask = 16'hE6A2;
defparam \Mux1~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N20
cycloneive_lcell_comb \Mux1~16 (
// Equation(s):
// \Mux1~16_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Mux1~13_combout )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & (\Mux1~15_combout )))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Mux1~15_combout ),
	.datad(\Mux1~13_combout ),
	.cin(gnd),
	.combout(\Mux1~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~16 .lut_mask = 16'hBA98;
defparam \Mux1~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y29_N17
dffeas \Reg[31][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][28] .is_wysiwyg = "true";
defparam \Reg[31][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N1
dffeas \Reg[23][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][28] .is_wysiwyg = "true";
defparam \Reg[23][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N27
dffeas \Reg[19][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][28] .is_wysiwyg = "true";
defparam \Reg[19][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N18
cycloneive_lcell_comb \Reg[27][28]~feeder (
// Equation(s):
// \Reg[27][28]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat20),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[27][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[27][28]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[27][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y29_N19
dffeas \Reg[27][28] (
	.clk(!CLK),
	.d(\Reg[27][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][28] .is_wysiwyg = "true";
defparam \Reg[27][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N26
cycloneive_lcell_comb \Mux3~7 (
// Equation(s):
// \Mux3~7_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[27][28]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & (\Reg[19][28]~q )))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[19][28]~q ),
	.datad(\Reg[27][28]~q ),
	.cin(gnd),
	.combout(\Mux3~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~7 .lut_mask = 16'hBA98;
defparam \Mux3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N2
cycloneive_lcell_comb \Mux3~8 (
// Equation(s):
// \Mux3~8_combout  = (ifid_ifinstr_o_23 & ((\Mux3~7_combout  & (\Reg[31][28]~q )) # (!\Mux3~7_combout  & ((\Reg[23][28]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux3~7_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[31][28]~q ),
	.datac(\Reg[23][28]~q ),
	.datad(\Mux3~7_combout ),
	.cin(gnd),
	.combout(\Mux3~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~8 .lut_mask = 16'hDDA0;
defparam \Mux3~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N12
cycloneive_lcell_comb \Reg[29][28]~feeder (
// Equation(s):
// \Reg[29][28]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat20),
	.cin(gnd),
	.combout(\Reg[29][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[29][28]~feeder .lut_mask = 16'hFF00;
defparam \Reg[29][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N13
dffeas \Reg[29][28] (
	.clk(!CLK),
	.d(\Reg[29][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][28] .is_wysiwyg = "true";
defparam \Reg[29][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N16
cycloneive_lcell_comb \Reg[21][28]~feeder (
// Equation(s):
// \Reg[21][28]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat20),
	.cin(gnd),
	.combout(\Reg[21][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[21][28]~feeder .lut_mask = 16'hFF00;
defparam \Reg[21][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N17
dffeas \Reg[21][28] (
	.clk(!CLK),
	.d(\Reg[21][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][28] .is_wysiwyg = "true";
defparam \Reg[21][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N0
cycloneive_lcell_comb \Reg[17][28]~feeder (
// Equation(s):
// \Reg[17][28]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat20),
	.cin(gnd),
	.combout(\Reg[17][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[17][28]~feeder .lut_mask = 16'hFF00;
defparam \Reg[17][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N1
dffeas \Reg[17][28] (
	.clk(!CLK),
	.d(\Reg[17][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][28] .is_wysiwyg = "true";
defparam \Reg[17][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N2
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[25][28]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[17][28]~q )))))

	.dataa(\Reg[25][28]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[17][28]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hEE30;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N6
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// \Mux3~1_combout  = (ifid_ifinstr_o_23 & ((\Mux3~0_combout  & (\Reg[29][28]~q )) # (!\Mux3~0_combout  & ((\Reg[21][28]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux3~0_combout ))))

	.dataa(\Reg[29][28]~q ),
	.datab(\Reg[21][28]~q ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux3~0_combout ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'hAFC0;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y34_N15
dffeas \Reg[28][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][28] .is_wysiwyg = "true";
defparam \Reg[28][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N30
cycloneive_lcell_comb \Reg[24][28]~feeder (
// Equation(s):
// \Reg[24][28]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat20),
	.cin(gnd),
	.combout(\Reg[24][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[24][28]~feeder .lut_mask = 16'hFF00;
defparam \Reg[24][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N31
dffeas \Reg[24][28] (
	.clk(!CLK),
	.d(\Reg[24][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][28] .is_wysiwyg = "true";
defparam \Reg[24][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y34_N29
dffeas \Reg[20][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][28] .is_wysiwyg = "true";
defparam \Reg[20][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y33_N9
dffeas \Reg[16][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][28] .is_wysiwyg = "true";
defparam \Reg[16][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N28
cycloneive_lcell_comb \Mux3~4 (
// Equation(s):
// \Mux3~4_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & (\Reg[20][28]~q )) # (!ifid_ifinstr_o_23 & ((\Reg[16][28]~q )))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[20][28]~q ),
	.datad(\Reg[16][28]~q ),
	.cin(gnd),
	.combout(\Mux3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~4 .lut_mask = 16'hD9C8;
defparam \Mux3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N20
cycloneive_lcell_comb \Mux3~5 (
// Equation(s):
// \Mux3~5_combout  = (ifid_ifinstr_o_24 & ((\Mux3~4_combout  & (\Reg[28][28]~q )) # (!\Mux3~4_combout  & ((\Reg[24][28]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux3~4_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[28][28]~q ),
	.datac(\Reg[24][28]~q ),
	.datad(\Mux3~4_combout ),
	.cin(gnd),
	.combout(\Mux3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~5 .lut_mask = 16'hDDA0;
defparam \Mux3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N17
dffeas \Reg[26][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][28] .is_wysiwyg = "true";
defparam \Reg[26][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y36_N5
dffeas \Reg[30][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][28] .is_wysiwyg = "true";
defparam \Reg[30][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y33_N27
dffeas \Reg[22][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][28] .is_wysiwyg = "true";
defparam \Reg[22][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N6
cycloneive_lcell_comb \Reg[18][28]~feeder (
// Equation(s):
// \Reg[18][28]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat20),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[18][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[18][28]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[18][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N7
dffeas \Reg[18][28] (
	.clk(!CLK),
	.d(\Reg[18][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][28] .is_wysiwyg = "true";
defparam \Reg[18][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N26
cycloneive_lcell_comb \Mux3~2 (
// Equation(s):
// \Mux3~2_combout  = (ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24) # ((\Reg[22][28]~q )))) # (!ifid_ifinstr_o_23 & (!ifid_ifinstr_o_24 & ((\Reg[18][28]~q ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[22][28]~q ),
	.datad(\Reg[18][28]~q ),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~2 .lut_mask = 16'hB9A8;
defparam \Mux3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N20
cycloneive_lcell_comb \Mux3~3 (
// Equation(s):
// \Mux3~3_combout  = (ifid_ifinstr_o_24 & ((\Mux3~2_combout  & ((\Reg[30][28]~q ))) # (!\Mux3~2_combout  & (\Reg[26][28]~q )))) # (!ifid_ifinstr_o_24 & (((\Mux3~2_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[26][28]~q ),
	.datac(\Reg[30][28]~q ),
	.datad(\Mux3~2_combout ),
	.cin(gnd),
	.combout(\Mux3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~3 .lut_mask = 16'hF588;
defparam \Mux3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N2
cycloneive_lcell_comb \Mux3~6 (
// Equation(s):
// \Mux3~6_combout  = (ifid_ifinstr_o_21 & (ifid_ifinstr_o_22)) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Mux3~3_combout ))) # (!ifid_ifinstr_o_22 & (\Mux3~5_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Mux3~5_combout ),
	.datad(\Mux3~3_combout ),
	.cin(gnd),
	.combout(\Mux3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~6 .lut_mask = 16'hDC98;
defparam \Mux3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N30
cycloneive_lcell_comb \Reg[6][28]~feeder (
// Equation(s):
// \Reg[6][28]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat20),
	.cin(gnd),
	.combout(\Reg[6][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[6][28]~feeder .lut_mask = 16'hFF00;
defparam \Reg[6][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N31
dffeas \Reg[6][28] (
	.clk(!CLK),
	.d(\Reg[6][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][28] .is_wysiwyg = "true";
defparam \Reg[6][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N15
dffeas \Reg[4][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][28] .is_wysiwyg = "true";
defparam \Reg[4][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N13
dffeas \Reg[5][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][28] .is_wysiwyg = "true";
defparam \Reg[5][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N12
cycloneive_lcell_comb \Mux3~10 (
// Equation(s):
// \Mux3~10_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[5][28]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[4][28]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[4][28]~q ),
	.datac(\Reg[5][28]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux3~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~10 .lut_mask = 16'hFA44;
defparam \Mux3~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N13
dffeas \Reg[7][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][28] .is_wysiwyg = "true";
defparam \Reg[7][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N28
cycloneive_lcell_comb \Mux3~11 (
// Equation(s):
// \Mux3~11_combout  = (\Mux3~10_combout  & (((\Reg[7][28]~q ) # (!ifid_ifinstr_o_22)))) # (!\Mux3~10_combout  & (\Reg[6][28]~q  & (ifid_ifinstr_o_22)))

	.dataa(\Reg[6][28]~q ),
	.datab(\Mux3~10_combout ),
	.datac(ifid_ifinstr_o_22),
	.datad(\Reg[7][28]~q ),
	.cin(gnd),
	.combout(\Mux3~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~11 .lut_mask = 16'hEC2C;
defparam \Mux3~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N7
dffeas \Reg[15][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][28] .is_wysiwyg = "true";
defparam \Reg[15][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N25
dffeas \Reg[12][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][28] .is_wysiwyg = "true";
defparam \Reg[12][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N19
dffeas \Reg[13][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][28] .is_wysiwyg = "true";
defparam \Reg[13][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N18
cycloneive_lcell_comb \Mux3~17 (
// Equation(s):
// \Mux3~17_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[13][28]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[12][28]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[12][28]~q ),
	.datac(\Reg[13][28]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux3~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~17 .lut_mask = 16'hFA44;
defparam \Mux3~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N1
dffeas \Reg[14][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][28] .is_wysiwyg = "true";
defparam \Reg[14][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N0
cycloneive_lcell_comb \Mux3~18 (
// Equation(s):
// \Mux3~18_combout  = (\Mux3~17_combout  & ((\Reg[15][28]~q ) # ((!ifid_ifinstr_o_22)))) # (!\Mux3~17_combout  & (((\Reg[14][28]~q  & ifid_ifinstr_o_22))))

	.dataa(\Reg[15][28]~q ),
	.datab(\Mux3~17_combout ),
	.datac(\Reg[14][28]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux3~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~18 .lut_mask = 16'hB8CC;
defparam \Mux3~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N25
dffeas \Reg[9][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][28] .is_wysiwyg = "true";
defparam \Reg[9][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y33_N15
dffeas \Reg[11][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][28] .is_wysiwyg = "true";
defparam \Reg[11][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N14
cycloneive_lcell_comb \Mux3~13 (
// Equation(s):
// \Mux3~13_combout  = (\Mux3~12_combout  & (((\Reg[11][28]~q ) # (!ifid_ifinstr_o_21)))) # (!\Mux3~12_combout  & (\Reg[9][28]~q  & ((ifid_ifinstr_o_21))))

	.dataa(\Mux3~12_combout ),
	.datab(\Reg[9][28]~q ),
	.datac(\Reg[11][28]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux3~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~13 .lut_mask = 16'hE4AA;
defparam \Mux3~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N17
dffeas \Reg[1][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][28] .is_wysiwyg = "true";
defparam \Reg[1][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N11
dffeas \Reg[3][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][28] .is_wysiwyg = "true";
defparam \Reg[3][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N16
cycloneive_lcell_comb \Mux3~14 (
// Equation(s):
// \Mux3~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][28]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][28]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[1][28]~q ),
	.datad(\Reg[3][28]~q ),
	.cin(gnd),
	.combout(\Mux3~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~14 .lut_mask = 16'hC840;
defparam \Mux3~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N31
dffeas \Reg[2][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][28] .is_wysiwyg = "true";
defparam \Reg[2][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N14
cycloneive_lcell_comb \Mux3~15 (
// Equation(s):
// \Mux3~15_combout  = (\Mux3~14_combout ) # ((ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & \Reg[2][28]~q )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux3~14_combout ),
	.datad(\Reg[2][28]~q ),
	.cin(gnd),
	.combout(\Mux3~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~15 .lut_mask = 16'hF2F0;
defparam \Mux3~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N10
cycloneive_lcell_comb \Mux3~16 (
// Equation(s):
// \Mux3~16_combout  = (ifid_ifinstr_o_24 & ((\Mux3~13_combout ) # ((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & (((\Mux3~15_combout  & !ifid_ifinstr_o_23))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux3~13_combout ),
	.datac(\Mux3~15_combout ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux3~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~16 .lut_mask = 16'hAAD8;
defparam \Mux3~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N5
dffeas \Reg[23][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][26] .is_wysiwyg = "true";
defparam \Reg[23][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N26
cycloneive_lcell_comb \Reg[31][26]~feeder (
// Equation(s):
// \Reg[31][26]~feeder_combout  = \wdat~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat21),
	.cin(gnd),
	.combout(\Reg[31][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[31][26]~feeder .lut_mask = 16'hFF00;
defparam \Reg[31][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N27
dffeas \Reg[31][26] (
	.clk(!CLK),
	.d(\Reg[31][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][26] .is_wysiwyg = "true";
defparam \Reg[31][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N23
dffeas \Reg[19][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][26] .is_wysiwyg = "true";
defparam \Reg[19][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N22
cycloneive_lcell_comb \Mux5~7 (
// Equation(s):
// \Mux5~7_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[27][26]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[19][26]~q )))))

	.dataa(\Reg[27][26]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[19][26]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux5~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~7 .lut_mask = 16'hEE30;
defparam \Mux5~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N8
cycloneive_lcell_comb \Mux5~8 (
// Equation(s):
// \Mux5~8_combout  = (ifid_ifinstr_o_23 & ((\Mux5~7_combout  & ((\Reg[31][26]~q ))) # (!\Mux5~7_combout  & (\Reg[23][26]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux5~7_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[23][26]~q ),
	.datac(\Reg[31][26]~q ),
	.datad(\Mux5~7_combout ),
	.cin(gnd),
	.combout(\Mux5~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~8 .lut_mask = 16'hF588;
defparam \Mux5~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N10
cycloneive_lcell_comb \Reg[16][26]~feeder (
// Equation(s):
// \Reg[16][26]~feeder_combout  = \wdat~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat21),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[16][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[16][26]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[16][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y34_N11
dffeas \Reg[16][26] (
	.clk(!CLK),
	.d(\Reg[16][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][26] .is_wysiwyg = "true";
defparam \Reg[16][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y34_N25
dffeas \Reg[20][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][26] .is_wysiwyg = "true";
defparam \Reg[20][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N24
cycloneive_lcell_comb \Mux5~4 (
// Equation(s):
// \Mux5~4_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[20][26]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[16][26]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[16][26]~q ),
	.datac(\Reg[20][26]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~4 .lut_mask = 16'hFA44;
defparam \Mux5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y34_N7
dffeas \Reg[28][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][26] .is_wysiwyg = "true";
defparam \Reg[28][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y34_N1
dffeas \Reg[24][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][26] .is_wysiwyg = "true";
defparam \Reg[24][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N6
cycloneive_lcell_comb \Mux5~5 (
// Equation(s):
// \Mux5~5_combout  = (ifid_ifinstr_o_24 & ((\Mux5~4_combout  & (\Reg[28][26]~q )) # (!\Mux5~4_combout  & ((\Reg[24][26]~q ))))) # (!ifid_ifinstr_o_24 & (\Mux5~4_combout ))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux5~4_combout ),
	.datac(\Reg[28][26]~q ),
	.datad(\Reg[24][26]~q ),
	.cin(gnd),
	.combout(\Mux5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~5 .lut_mask = 16'hE6C4;
defparam \Mux5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N29
dffeas \Reg[18][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][26] .is_wysiwyg = "true";
defparam \Reg[18][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N26
cycloneive_lcell_comb \Reg[22][26]~feeder (
// Equation(s):
// \Reg[22][26]~feeder_combout  = \wdat~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat21),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[22][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[22][26]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[22][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N27
dffeas \Reg[22][26] (
	.clk(!CLK),
	.d(\Reg[22][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][26] .is_wysiwyg = "true";
defparam \Reg[22][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N28
cycloneive_lcell_comb \Mux5~2 (
// Equation(s):
// \Mux5~2_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[22][26]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[18][26]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[18][26]~q ),
	.datad(\Reg[22][26]~q ),
	.cin(gnd),
	.combout(\Mux5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~2 .lut_mask = 16'hDC98;
defparam \Mux5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N15
dffeas \Reg[26][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][26] .is_wysiwyg = "true";
defparam \Reg[26][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N16
cycloneive_lcell_comb \Mux5~3 (
// Equation(s):
// \Mux5~3_combout  = (ifid_ifinstr_o_24 & ((\Mux5~2_combout  & (\Reg[30][26]~q )) # (!\Mux5~2_combout  & ((\Reg[26][26]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux5~2_combout ))))

	.dataa(\Reg[30][26]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Mux5~2_combout ),
	.datad(\Reg[26][26]~q ),
	.cin(gnd),
	.combout(\Mux5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~3 .lut_mask = 16'hBCB0;
defparam \Mux5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N14
cycloneive_lcell_comb \Mux5~6 (
// Equation(s):
// \Mux5~6_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Mux5~3_combout ))) # (!ifid_ifinstr_o_22 & (\Mux5~5_combout ))))

	.dataa(\Mux5~5_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(ifid_ifinstr_o_22),
	.datad(\Mux5~3_combout ),
	.cin(gnd),
	.combout(\Mux5~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~6 .lut_mask = 16'hF2C2;
defparam \Mux5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N21
dffeas \Reg[25][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][26] .is_wysiwyg = "true";
defparam \Reg[25][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N11
dffeas \Reg[17][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][26] .is_wysiwyg = "true";
defparam \Reg[17][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N20
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// \Mux5~0_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[25][26]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & ((\Reg[17][26]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[25][26]~q ),
	.datad(\Reg[17][26]~q ),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'hB9A8;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N29
dffeas \Reg[29][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][26] .is_wysiwyg = "true";
defparam \Reg[29][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N29
dffeas \Reg[21][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][26] .is_wysiwyg = "true";
defparam \Reg[21][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N28
cycloneive_lcell_comb \Mux5~1 (
// Equation(s):
// \Mux5~1_combout  = (\Mux5~0_combout  & ((\Reg[29][26]~q ) # ((!ifid_ifinstr_o_23)))) # (!\Mux5~0_combout  & (((\Reg[21][26]~q  & ifid_ifinstr_o_23))))

	.dataa(\Mux5~0_combout ),
	.datab(\Reg[29][26]~q ),
	.datac(\Reg[21][26]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~1 .lut_mask = 16'hD8AA;
defparam \Mux5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y37_N14
cycloneive_lcell_comb \Reg[12][26]~feeder (
// Equation(s):
// \Reg[12][26]~feeder_combout  = \wdat~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat21),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[12][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[12][26]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[12][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y37_N15
dffeas \Reg[12][26] (
	.clk(!CLK),
	.d(\Reg[12][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][26] .is_wysiwyg = "true";
defparam \Reg[12][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y37_N1
dffeas \Reg[13][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][26] .is_wysiwyg = "true";
defparam \Reg[13][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y37_N0
cycloneive_lcell_comb \Mux5~17 (
// Equation(s):
// \Mux5~17_combout  = (ifid_ifinstr_o_21 & (((\Reg[13][26]~q ) # (ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & (\Reg[12][26]~q  & ((!ifid_ifinstr_o_22))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[12][26]~q ),
	.datac(\Reg[13][26]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux5~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~17 .lut_mask = 16'hAAE4;
defparam \Mux5~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N19
dffeas \Reg[15][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][26] .is_wysiwyg = "true";
defparam \Reg[15][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N25
dffeas \Reg[14][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][26] .is_wysiwyg = "true";
defparam \Reg[14][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N18
cycloneive_lcell_comb \Mux5~18 (
// Equation(s):
// \Mux5~18_combout  = (\Mux5~17_combout  & (((\Reg[15][26]~q )) # (!ifid_ifinstr_o_22))) # (!\Mux5~17_combout  & (ifid_ifinstr_o_22 & ((\Reg[14][26]~q ))))

	.dataa(\Mux5~17_combout ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[15][26]~q ),
	.datad(\Reg[14][26]~q ),
	.cin(gnd),
	.combout(\Mux5~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~18 .lut_mask = 16'hE6A2;
defparam \Mux5~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y39_N15
dffeas \Reg[7][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][26] .is_wysiwyg = "true";
defparam \Reg[7][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N17
dffeas \Reg[6][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][26] .is_wysiwyg = "true";
defparam \Reg[6][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N5
dffeas \Reg[5][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][26] .is_wysiwyg = "true";
defparam \Reg[5][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N4
cycloneive_lcell_comb \Mux5~10 (
// Equation(s):
// \Mux5~10_combout  = (ifid_ifinstr_o_21 & (((\Reg[5][26]~q ) # (ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & (\Reg[4][26]~q  & ((!ifid_ifinstr_o_22))))

	.dataa(\Reg[4][26]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[5][26]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux5~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~10 .lut_mask = 16'hCCE2;
defparam \Mux5~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N16
cycloneive_lcell_comb \Mux5~11 (
// Equation(s):
// \Mux5~11_combout  = (ifid_ifinstr_o_22 & ((\Mux5~10_combout  & (\Reg[7][26]~q )) # (!\Mux5~10_combout  & ((\Reg[6][26]~q ))))) # (!ifid_ifinstr_o_22 & (((\Mux5~10_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[7][26]~q ),
	.datac(\Reg[6][26]~q ),
	.datad(\Mux5~10_combout ),
	.cin(gnd),
	.combout(\Mux5~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~11 .lut_mask = 16'hDDA0;
defparam \Mux5~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y35_N1
dffeas \Reg[3][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][26] .is_wysiwyg = "true";
defparam \Reg[3][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y35_N19
dffeas \Reg[1][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][26] .is_wysiwyg = "true";
defparam \Reg[1][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N0
cycloneive_lcell_comb \Mux5~14 (
// Equation(s):
// \Mux5~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[3][26]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[1][26]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[3][26]~q ),
	.datad(\Reg[1][26]~q ),
	.cin(gnd),
	.combout(\Mux5~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~14 .lut_mask = 16'hA280;
defparam \Mux5~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y36_N29
dffeas \Reg[2][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][26] .is_wysiwyg = "true";
defparam \Reg[2][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N28
cycloneive_lcell_comb \Mux5~15 (
// Equation(s):
// \Mux5~15_combout  = (\Mux5~14_combout ) # ((!ifid_ifinstr_o_21 & (\Reg[2][26]~q  & ifid_ifinstr_o_22)))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux5~14_combout ),
	.datac(\Reg[2][26]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux5~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~15 .lut_mask = 16'hDCCC;
defparam \Mux5~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N8
cycloneive_lcell_comb \Reg[11][26]~feeder (
// Equation(s):
// \Reg[11][26]~feeder_combout  = \wdat~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat21),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[11][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[11][26]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[11][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y36_N9
dffeas \Reg[11][26] (
	.clk(!CLK),
	.d(\Reg[11][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][26] .is_wysiwyg = "true";
defparam \Reg[11][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N23
dffeas \Reg[8][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][26] .is_wysiwyg = "true";
defparam \Reg[8][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N13
dffeas \Reg[10][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat21),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][26] .is_wysiwyg = "true";
defparam \Reg[10][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N22
cycloneive_lcell_comb \Mux5~12 (
// Equation(s):
// \Mux5~12_combout  = (ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21) # ((\Reg[10][26]~q )))) # (!ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & (\Reg[8][26]~q )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[8][26]~q ),
	.datad(\Reg[10][26]~q ),
	.cin(gnd),
	.combout(\Mux5~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~12 .lut_mask = 16'hBA98;
defparam \Mux5~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N2
cycloneive_lcell_comb \Reg[9][26]~feeder (
// Equation(s):
// \Reg[9][26]~feeder_combout  = \wdat~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat21),
	.cin(gnd),
	.combout(\Reg[9][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[9][26]~feeder .lut_mask = 16'hFF00;
defparam \Reg[9][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y32_N3
dffeas \Reg[9][26] (
	.clk(!CLK),
	.d(\Reg[9][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][26] .is_wysiwyg = "true";
defparam \Reg[9][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N2
cycloneive_lcell_comb \Mux5~13 (
// Equation(s):
// \Mux5~13_combout  = (ifid_ifinstr_o_21 & ((\Mux5~12_combout  & (\Reg[11][26]~q )) # (!\Mux5~12_combout  & ((\Reg[9][26]~q ))))) # (!ifid_ifinstr_o_21 & (((\Mux5~12_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[11][26]~q ),
	.datac(\Mux5~12_combout ),
	.datad(\Reg[9][26]~q ),
	.cin(gnd),
	.combout(\Mux5~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~13 .lut_mask = 16'hDAD0;
defparam \Mux5~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N22
cycloneive_lcell_comb \Mux5~16 (
// Equation(s):
// \Mux5~16_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23) # (\Mux5~13_combout )))) # (!ifid_ifinstr_o_24 & (\Mux5~15_combout  & (!ifid_ifinstr_o_23)))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux5~15_combout ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux5~13_combout ),
	.cin(gnd),
	.combout(\Mux5~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~16 .lut_mask = 16'hAEA4;
defparam \Mux5~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N5
dffeas \Reg[25][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][27] .is_wysiwyg = "true";
defparam \Reg[25][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N21
dffeas \Reg[29][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][27] .is_wysiwyg = "true";
defparam \Reg[29][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N7
dffeas \Reg[17][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][27] .is_wysiwyg = "true";
defparam \Reg[17][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N15
dffeas \Reg[21][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][27] .is_wysiwyg = "true";
defparam \Reg[21][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N6
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// \Mux4~0_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[21][27]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[17][27]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[17][27]~q ),
	.datad(\Reg[21][27]~q ),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'hDC98;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N20
cycloneive_lcell_comb \Mux4~1 (
// Equation(s):
// \Mux4~1_combout  = (ifid_ifinstr_o_24 & ((\Mux4~0_combout  & ((\Reg[29][27]~q ))) # (!\Mux4~0_combout  & (\Reg[25][27]~q )))) # (!ifid_ifinstr_o_24 & (((\Mux4~0_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[25][27]~q ),
	.datac(\Reg[29][27]~q ),
	.datad(\Mux4~0_combout ),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~1 .lut_mask = 16'hF588;
defparam \Mux4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N9
dffeas \Reg[27][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][27] .is_wysiwyg = "true";
defparam \Reg[27][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N6
cycloneive_lcell_comb \Reg[23][27]~feeder (
// Equation(s):
// \Reg[23][27]~feeder_combout  = \wdat~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat22),
	.cin(gnd),
	.combout(\Reg[23][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[23][27]~feeder .lut_mask = 16'hFF00;
defparam \Reg[23][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N7
dffeas \Reg[23][27] (
	.clk(!CLK),
	.d(\Reg[23][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][27] .is_wysiwyg = "true";
defparam \Reg[23][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N25
dffeas \Reg[19][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][27] .is_wysiwyg = "true";
defparam \Reg[19][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N24
cycloneive_lcell_comb \Mux4~7 (
// Equation(s):
// \Mux4~7_combout  = (ifid_ifinstr_o_23 & ((\Reg[23][27]~q ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((\Reg[19][27]~q  & !ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[23][27]~q ),
	.datac(\Reg[19][27]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux4~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~7 .lut_mask = 16'hAAD8;
defparam \Mux4~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N23
dffeas \Reg[31][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][27] .is_wysiwyg = "true";
defparam \Reg[31][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N26
cycloneive_lcell_comb \Mux4~8 (
// Equation(s):
// \Mux4~8_combout  = (\Mux4~7_combout  & (((\Reg[31][27]~q ) # (!ifid_ifinstr_o_24)))) # (!\Mux4~7_combout  & (\Reg[27][27]~q  & (ifid_ifinstr_o_24)))

	.dataa(\Reg[27][27]~q ),
	.datab(\Mux4~7_combout ),
	.datac(ifid_ifinstr_o_24),
	.datad(\Reg[31][27]~q ),
	.cin(gnd),
	.combout(\Mux4~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~8 .lut_mask = 16'hEC2C;
defparam \Mux4~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N2
cycloneive_lcell_comb \Reg[20][27]~feeder (
// Equation(s):
// \Reg[20][27]~feeder_combout  = \wdat~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat22),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[20][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[20][27]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[20][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N3
dffeas \Reg[20][27] (
	.clk(!CLK),
	.d(\Reg[20][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][27] .is_wysiwyg = "true";
defparam \Reg[20][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N1
dffeas \Reg[24][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][27] .is_wysiwyg = "true";
defparam \Reg[24][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N0
cycloneive_lcell_comb \Mux4~4 (
// Equation(s):
// \Mux4~4_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Reg[24][27]~q ))) # (!ifid_ifinstr_o_24 & (\Reg[16][27]~q ))))

	.dataa(\Reg[16][27]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[24][27]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~4 .lut_mask = 16'hFC22;
defparam \Mux4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N10
cycloneive_lcell_comb \Mux4~5 (
// Equation(s):
// \Mux4~5_combout  = (\Mux4~4_combout  & ((\Reg[28][27]~q ) # ((!ifid_ifinstr_o_23)))) # (!\Mux4~4_combout  & (((\Reg[20][27]~q  & ifid_ifinstr_o_23))))

	.dataa(\Reg[28][27]~q ),
	.datab(\Reg[20][27]~q ),
	.datac(\Mux4~4_combout ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~5 .lut_mask = 16'hACF0;
defparam \Mux4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N3
dffeas \Reg[22][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][27] .is_wysiwyg = "true";
defparam \Reg[22][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N5
dffeas \Reg[18][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][27] .is_wysiwyg = "true";
defparam \Reg[18][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N2
cycloneive_lcell_comb \Reg[26][27]~feeder (
// Equation(s):
// \Reg[26][27]~feeder_combout  = \wdat~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat22),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[26][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[26][27]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[26][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N3
dffeas \Reg[26][27] (
	.clk(!CLK),
	.d(\Reg[26][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][27] .is_wysiwyg = "true";
defparam \Reg[26][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N4
cycloneive_lcell_comb \Mux4~2 (
// Equation(s):
// \Mux4~2_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[26][27]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & (\Reg[18][27]~q )))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[18][27]~q ),
	.datad(\Reg[26][27]~q ),
	.cin(gnd),
	.combout(\Mux4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~2 .lut_mask = 16'hBA98;
defparam \Mux4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N20
cycloneive_lcell_comb \Mux4~3 (
// Equation(s):
// \Mux4~3_combout  = (\Mux4~2_combout  & ((\Reg[30][27]~q ) # ((!ifid_ifinstr_o_23)))) # (!\Mux4~2_combout  & (((\Reg[22][27]~q  & ifid_ifinstr_o_23))))

	.dataa(\Reg[30][27]~q ),
	.datab(\Reg[22][27]~q ),
	.datac(\Mux4~2_combout ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~3 .lut_mask = 16'hACF0;
defparam \Mux4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N16
cycloneive_lcell_comb \Mux4~6 (
// Equation(s):
// \Mux4~6_combout  = (ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21) # ((\Mux4~3_combout )))) # (!ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & (\Mux4~5_combout )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux4~5_combout ),
	.datad(\Mux4~3_combout ),
	.cin(gnd),
	.combout(\Mux4~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~6 .lut_mask = 16'hBA98;
defparam \Mux4~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y31_N19
dffeas \Reg[11][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][27] .is_wysiwyg = "true";
defparam \Reg[11][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y32_N29
dffeas \Reg[9][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][27] .is_wysiwyg = "true";
defparam \Reg[9][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N1
dffeas \Reg[10][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][27] .is_wysiwyg = "true";
defparam \Reg[10][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N7
dffeas \Reg[8][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][27] .is_wysiwyg = "true";
defparam \Reg[8][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N0
cycloneive_lcell_comb \Mux4~10 (
// Equation(s):
// \Mux4~10_combout  = (ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21) # ((\Reg[10][27]~q )))) # (!ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & ((\Reg[8][27]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[10][27]~q ),
	.datad(\Reg[8][27]~q ),
	.cin(gnd),
	.combout(\Mux4~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~10 .lut_mask = 16'hB9A8;
defparam \Mux4~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N28
cycloneive_lcell_comb \Mux4~11 (
// Equation(s):
// \Mux4~11_combout  = (ifid_ifinstr_o_21 & ((\Mux4~10_combout  & (\Reg[11][27]~q )) # (!\Mux4~10_combout  & ((\Reg[9][27]~q ))))) # (!ifid_ifinstr_o_21 & (((\Mux4~10_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[11][27]~q ),
	.datac(\Reg[9][27]~q ),
	.datad(\Mux4~10_combout ),
	.cin(gnd),
	.combout(\Mux4~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~11 .lut_mask = 16'hDDA0;
defparam \Mux4~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N12
cycloneive_lcell_comb \Reg[14][27]~feeder (
// Equation(s):
// \Reg[14][27]~feeder_combout  = \wdat~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat22),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[14][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[14][27]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[14][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N13
dffeas \Reg[14][27] (
	.clk(!CLK),
	.d(\Reg[14][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][27] .is_wysiwyg = "true";
defparam \Reg[14][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N27
dffeas \Reg[12][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][27] .is_wysiwyg = "true";
defparam \Reg[12][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N8
cycloneive_lcell_comb \Mux4~17 (
// Equation(s):
// \Mux4~17_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[13][27]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[12][27]~q )))))

	.dataa(\Reg[13][27]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[12][27]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux4~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~17 .lut_mask = 16'hEE30;
defparam \Mux4~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N30
cycloneive_lcell_comb \Reg[15][27]~feeder (
// Equation(s):
// \Reg[15][27]~feeder_combout  = \wdat~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat22),
	.cin(gnd),
	.combout(\Reg[15][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[15][27]~feeder .lut_mask = 16'hFF00;
defparam \Reg[15][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N31
dffeas \Reg[15][27] (
	.clk(!CLK),
	.d(\Reg[15][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][27] .is_wysiwyg = "true";
defparam \Reg[15][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N14
cycloneive_lcell_comb \Mux4~18 (
// Equation(s):
// \Mux4~18_combout  = (ifid_ifinstr_o_22 & ((\Mux4~17_combout  & ((\Reg[15][27]~q ))) # (!\Mux4~17_combout  & (\Reg[14][27]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux4~17_combout ))))

	.dataa(\Reg[14][27]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Mux4~17_combout ),
	.datad(\Reg[15][27]~q ),
	.cin(gnd),
	.combout(\Mux4~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~18 .lut_mask = 16'hF838;
defparam \Mux4~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y39_N9
dffeas \Reg[6][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][27] .is_wysiwyg = "true";
defparam \Reg[6][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y39_N7
dffeas \Reg[7][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][27] .is_wysiwyg = "true";
defparam \Reg[7][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N25
dffeas \Reg[5][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][27] .is_wysiwyg = "true";
defparam \Reg[5][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N7
dffeas \Reg[4][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][27] .is_wysiwyg = "true";
defparam \Reg[4][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N6
cycloneive_lcell_comb \Mux4~12 (
// Equation(s):
// \Mux4~12_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[5][27]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[4][27]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[5][27]~q ),
	.datac(\Reg[4][27]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux4~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~12 .lut_mask = 16'hEE50;
defparam \Mux4~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N6
cycloneive_lcell_comb \Mux4~13 (
// Equation(s):
// \Mux4~13_combout  = (ifid_ifinstr_o_22 & ((\Mux4~12_combout  & ((\Reg[7][27]~q ))) # (!\Mux4~12_combout  & (\Reg[6][27]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux4~12_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[6][27]~q ),
	.datac(\Reg[7][27]~q ),
	.datad(\Mux4~12_combout ),
	.cin(gnd),
	.combout(\Mux4~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~13 .lut_mask = 16'hF588;
defparam \Mux4~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N21
dffeas \Reg[3][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][27] .is_wysiwyg = "true";
defparam \Reg[3][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N3
dffeas \Reg[1][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][27] .is_wysiwyg = "true";
defparam \Reg[1][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N20
cycloneive_lcell_comb \Mux4~14 (
// Equation(s):
// \Mux4~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[3][27]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[1][27]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[3][27]~q ),
	.datad(\Reg[1][27]~q ),
	.cin(gnd),
	.combout(\Mux4~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~14 .lut_mask = 16'hC480;
defparam \Mux4~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y31_N9
dffeas \Reg[2][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][27] .is_wysiwyg = "true";
defparam \Reg[2][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N8
cycloneive_lcell_comb \Mux4~15 (
// Equation(s):
// \Mux4~15_combout  = (\Mux4~14_combout ) # ((ifid_ifinstr_o_22 & (\Reg[2][27]~q  & !ifid_ifinstr_o_21)))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Mux4~14_combout ),
	.datac(\Reg[2][27]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux4~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~15 .lut_mask = 16'hCCEC;
defparam \Mux4~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N2
cycloneive_lcell_comb \Mux4~16 (
// Equation(s):
// \Mux4~16_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & (\Mux4~13_combout )) # (!ifid_ifinstr_o_23 & ((\Mux4~15_combout )))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Mux4~13_combout ),
	.datad(\Mux4~15_combout ),
	.cin(gnd),
	.combout(\Mux4~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~16 .lut_mask = 16'hD9C8;
defparam \Mux4~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N6
cycloneive_lcell_comb \Reg[31][25]~feeder (
// Equation(s):
// \Reg[31][25]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat23),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[31][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[31][25]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[31][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N7
dffeas \Reg[31][25] (
	.clk(!CLK),
	.d(\Reg[31][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][25] .is_wysiwyg = "true";
defparam \Reg[31][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N9
dffeas \Reg[27][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][25] .is_wysiwyg = "true";
defparam \Reg[27][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y29_N29
dffeas \Reg[23][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][25] .is_wysiwyg = "true";
defparam \Reg[23][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N7
dffeas \Reg[19][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][25] .is_wysiwyg = "true";
defparam \Reg[19][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N28
cycloneive_lcell_comb \Mux6~7 (
// Equation(s):
// \Mux6~7_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & (\Reg[23][25]~q )) # (!ifid_ifinstr_o_23 & ((\Reg[19][25]~q )))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[23][25]~q ),
	.datad(\Reg[19][25]~q ),
	.cin(gnd),
	.combout(\Mux6~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~7 .lut_mask = 16'hD9C8;
defparam \Mux6~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N8
cycloneive_lcell_comb \Mux6~8 (
// Equation(s):
// \Mux6~8_combout  = (ifid_ifinstr_o_24 & ((\Mux6~7_combout  & (\Reg[31][25]~q )) # (!\Mux6~7_combout  & ((\Reg[27][25]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux6~7_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[31][25]~q ),
	.datac(\Reg[27][25]~q ),
	.datad(\Mux6~7_combout ),
	.cin(gnd),
	.combout(\Mux6~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~8 .lut_mask = 16'hDDA0;
defparam \Mux6~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N5
dffeas \Reg[22][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][25] .is_wysiwyg = "true";
defparam \Reg[22][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y30_N19
dffeas \Reg[30][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][25] .is_wysiwyg = "true";
defparam \Reg[30][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N25
dffeas \Reg[18][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][25] .is_wysiwyg = "true";
defparam \Reg[18][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N10
cycloneive_lcell_comb \Reg[26][25]~feeder (
// Equation(s):
// \Reg[26][25]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat23),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[26][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[26][25]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[26][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N11
dffeas \Reg[26][25] (
	.clk(!CLK),
	.d(\Reg[26][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][25] .is_wysiwyg = "true";
defparam \Reg[26][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N24
cycloneive_lcell_comb \Mux6~2 (
// Equation(s):
// \Mux6~2_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[26][25]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & (\Reg[18][25]~q )))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[18][25]~q ),
	.datad(\Reg[26][25]~q ),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~2 .lut_mask = 16'hBA98;
defparam \Mux6~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N8
cycloneive_lcell_comb \Mux6~3 (
// Equation(s):
// \Mux6~3_combout  = (ifid_ifinstr_o_23 & ((\Mux6~2_combout  & ((\Reg[30][25]~q ))) # (!\Mux6~2_combout  & (\Reg[22][25]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux6~2_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[22][25]~q ),
	.datac(\Reg[30][25]~q ),
	.datad(\Mux6~2_combout ),
	.cin(gnd),
	.combout(\Mux6~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~3 .lut_mask = 16'hF588;
defparam \Mux6~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N5
dffeas \Reg[28][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][25] .is_wysiwyg = "true";
defparam \Reg[28][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y33_N5
dffeas \Reg[20][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][25] .is_wysiwyg = "true";
defparam \Reg[20][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N11
dffeas \Reg[24][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][25] .is_wysiwyg = "true";
defparam \Reg[24][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N10
cycloneive_lcell_comb \Mux6~4 (
// Equation(s):
// \Mux6~4_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Reg[24][25]~q ))) # (!ifid_ifinstr_o_24 & (\Reg[16][25]~q ))))

	.dataa(\Reg[16][25]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[24][25]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux6~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~4 .lut_mask = 16'hFC22;
defparam \Mux6~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N4
cycloneive_lcell_comb \Mux6~5 (
// Equation(s):
// \Mux6~5_combout  = (ifid_ifinstr_o_23 & ((\Mux6~4_combout  & (\Reg[28][25]~q )) # (!\Mux6~4_combout  & ((\Reg[20][25]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux6~4_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[28][25]~q ),
	.datac(\Reg[20][25]~q ),
	.datad(\Mux6~4_combout ),
	.cin(gnd),
	.combout(\Mux6~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~5 .lut_mask = 16'hDDA0;
defparam \Mux6~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N26
cycloneive_lcell_comb \Mux6~6 (
// Equation(s):
// \Mux6~6_combout  = (ifid_ifinstr_o_21 & (ifid_ifinstr_o_22)) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Mux6~3_combout )) # (!ifid_ifinstr_o_22 & ((\Mux6~5_combout )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Mux6~3_combout ),
	.datad(\Mux6~5_combout ),
	.cin(gnd),
	.combout(\Mux6~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~6 .lut_mask = 16'hD9C8;
defparam \Mux6~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N9
dffeas \Reg[25][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][25] .is_wysiwyg = "true";
defparam \Reg[25][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y37_N23
dffeas \Reg[29][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][25] .is_wysiwyg = "true";
defparam \Reg[29][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N27
dffeas \Reg[17][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][25] .is_wysiwyg = "true";
defparam \Reg[17][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y37_N13
dffeas \Reg[21][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][25] .is_wysiwyg = "true";
defparam \Reg[21][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N26
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// \Mux6~0_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[21][25]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[17][25]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[17][25]~q ),
	.datad(\Reg[21][25]~q ),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'hDC98;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N22
cycloneive_lcell_comb \Mux6~1 (
// Equation(s):
// \Mux6~1_combout  = (ifid_ifinstr_o_24 & ((\Mux6~0_combout  & ((\Reg[29][25]~q ))) # (!\Mux6~0_combout  & (\Reg[25][25]~q )))) # (!ifid_ifinstr_o_24 & (((\Mux6~0_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[25][25]~q ),
	.datac(\Reg[29][25]~q ),
	.datad(\Mux6~0_combout ),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~1 .lut_mask = 16'hF588;
defparam \Mux6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N26
cycloneive_lcell_comb \Reg[9][25]~feeder (
// Equation(s):
// \Reg[9][25]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat23),
	.cin(gnd),
	.combout(\Reg[9][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[9][25]~feeder .lut_mask = 16'hFF00;
defparam \Reg[9][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y32_N27
dffeas \Reg[9][25] (
	.clk(!CLK),
	.d(\Reg[9][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][25] .is_wysiwyg = "true";
defparam \Reg[9][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y31_N7
dffeas \Reg[11][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][25] .is_wysiwyg = "true";
defparam \Reg[11][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N13
dffeas \Reg[10][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][25] .is_wysiwyg = "true";
defparam \Reg[10][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N12
cycloneive_lcell_comb \Mux6~10 (
// Equation(s):
// \Mux6~10_combout  = (ifid_ifinstr_o_22 & (((\Reg[10][25]~q ) # (ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & (\Reg[8][25]~q  & ((!ifid_ifinstr_o_21))))

	.dataa(\Reg[8][25]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[10][25]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux6~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~10 .lut_mask = 16'hCCE2;
defparam \Mux6~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N12
cycloneive_lcell_comb \Mux6~11 (
// Equation(s):
// \Mux6~11_combout  = (\Mux6~10_combout  & (((\Reg[11][25]~q ) # (!ifid_ifinstr_o_21)))) # (!\Mux6~10_combout  & (\Reg[9][25]~q  & ((ifid_ifinstr_o_21))))

	.dataa(\Reg[9][25]~q ),
	.datab(\Reg[11][25]~q ),
	.datac(\Mux6~10_combout ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux6~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~11 .lut_mask = 16'hCAF0;
defparam \Mux6~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y37_N17
dffeas \Reg[13][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][25] .is_wysiwyg = "true";
defparam \Reg[13][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y37_N6
cycloneive_lcell_comb \Reg[12][25]~feeder (
// Equation(s):
// \Reg[12][25]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat23),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[12][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[12][25]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[12][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y37_N7
dffeas \Reg[12][25] (
	.clk(!CLK),
	.d(\Reg[12][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][25] .is_wysiwyg = "true";
defparam \Reg[12][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y37_N16
cycloneive_lcell_comb \Mux6~17 (
// Equation(s):
// \Mux6~17_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[13][25]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[12][25]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[13][25]~q ),
	.datad(\Reg[12][25]~q ),
	.cin(gnd),
	.combout(\Mux6~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~17 .lut_mask = 16'hD9C8;
defparam \Mux6~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y37_N25
dffeas \Reg[14][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][25] .is_wysiwyg = "true";
defparam \Reg[14][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N30
cycloneive_lcell_comb \Reg[15][25]~feeder (
// Equation(s):
// \Reg[15][25]~feeder_combout  = \wdat~49_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat23),
	.cin(gnd),
	.combout(\Reg[15][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[15][25]~feeder .lut_mask = 16'hFF00;
defparam \Reg[15][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N31
dffeas \Reg[15][25] (
	.clk(!CLK),
	.d(\Reg[15][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][25] .is_wysiwyg = "true";
defparam \Reg[15][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N14
cycloneive_lcell_comb \Mux6~18 (
// Equation(s):
// \Mux6~18_combout  = (\Mux6~17_combout  & (((\Reg[15][25]~q )) # (!ifid_ifinstr_o_22))) # (!\Mux6~17_combout  & (ifid_ifinstr_o_22 & (\Reg[14][25]~q )))

	.dataa(\Mux6~17_combout ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[14][25]~q ),
	.datad(\Reg[15][25]~q ),
	.cin(gnd),
	.combout(\Mux6~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~18 .lut_mask = 16'hEA62;
defparam \Mux6~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y35_N3
dffeas \Reg[3][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][25] .is_wysiwyg = "true";
defparam \Reg[3][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y35_N29
dffeas \Reg[1][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][25] .is_wysiwyg = "true";
defparam \Reg[1][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N2
cycloneive_lcell_comb \Mux6~14 (
// Equation(s):
// \Mux6~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[3][25]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[1][25]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[3][25]~q ),
	.datad(\Reg[1][25]~q ),
	.cin(gnd),
	.combout(\Mux6~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~14 .lut_mask = 16'hA280;
defparam \Mux6~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y31_N21
dffeas \Reg[2][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][25] .is_wysiwyg = "true";
defparam \Reg[2][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N10
cycloneive_lcell_comb \Mux6~15 (
// Equation(s):
// \Mux6~15_combout  = (\Mux6~14_combout ) # ((!ifid_ifinstr_o_21 & (ifid_ifinstr_o_22 & \Reg[2][25]~q )))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Mux6~14_combout ),
	.datad(\Reg[2][25]~q ),
	.cin(gnd),
	.combout(\Mux6~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~15 .lut_mask = 16'hF4F0;
defparam \Mux6~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N13
dffeas \Reg[7][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][25] .is_wysiwyg = "true";
defparam \Reg[7][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y39_N7
dffeas \Reg[4][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][25] .is_wysiwyg = "true";
defparam \Reg[4][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y39_N5
dffeas \Reg[5][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][25] .is_wysiwyg = "true";
defparam \Reg[5][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N6
cycloneive_lcell_comb \Mux6~12 (
// Equation(s):
// \Mux6~12_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[5][25]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[4][25]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[4][25]~q ),
	.datad(\Reg[5][25]~q ),
	.cin(gnd),
	.combout(\Mux6~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~12 .lut_mask = 16'hDC98;
defparam \Mux6~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N12
cycloneive_lcell_comb \Mux6~13 (
// Equation(s):
// \Mux6~13_combout  = (ifid_ifinstr_o_22 & ((\Mux6~12_combout  & ((\Reg[7][25]~q ))) # (!\Mux6~12_combout  & (\Reg[6][25]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux6~12_combout ))))

	.dataa(\Reg[6][25]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[7][25]~q ),
	.datad(\Mux6~12_combout ),
	.cin(gnd),
	.combout(\Mux6~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~13 .lut_mask = 16'hF388;
defparam \Mux6~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N20
cycloneive_lcell_comb \Mux6~16 (
// Equation(s):
// \Mux6~16_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Mux6~13_combout ))) # (!ifid_ifinstr_o_23 & (\Mux6~15_combout ))))

	.dataa(\Mux6~15_combout ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Mux6~13_combout ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux6~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~16 .lut_mask = 16'hFC22;
defparam \Mux6~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N26
cycloneive_lcell_comb \Reg[18][24]~feeder (
// Equation(s):
// \Reg[18][24]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat24),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[18][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[18][24]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[18][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N27
dffeas \Reg[18][24] (
	.clk(!CLK),
	.d(\Reg[18][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][24] .is_wysiwyg = "true";
defparam \Reg[18][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N0
cycloneive_lcell_comb \Reg[22][24]~feeder (
// Equation(s):
// \Reg[22][24]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat24),
	.cin(gnd),
	.combout(\Reg[22][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[22][24]~feeder .lut_mask = 16'hFF00;
defparam \Reg[22][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N1
dffeas \Reg[22][24] (
	.clk(!CLK),
	.d(\Reg[22][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][24] .is_wysiwyg = "true";
defparam \Reg[22][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N18
cycloneive_lcell_comb \Mux7~2 (
// Equation(s):
// \Mux7~2_combout  = (ifid_ifinstr_o_23 & (((\Reg[22][24]~q ) # (ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (\Reg[18][24]~q  & ((!ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[18][24]~q ),
	.datac(\Reg[22][24]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~2 .lut_mask = 16'hAAE4;
defparam \Mux7~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N5
dffeas \Reg[26][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][24] .is_wysiwyg = "true";
defparam \Reg[26][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N6
cycloneive_lcell_comb \Reg[30][24]~feeder (
// Equation(s):
// \Reg[30][24]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat24),
	.cin(gnd),
	.combout(\Reg[30][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[30][24]~feeder .lut_mask = 16'hFF00;
defparam \Reg[30][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N7
dffeas \Reg[30][24] (
	.clk(!CLK),
	.d(\Reg[30][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][24] .is_wysiwyg = "true";
defparam \Reg[30][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N4
cycloneive_lcell_comb \Mux7~3 (
// Equation(s):
// \Mux7~3_combout  = (ifid_ifinstr_o_24 & ((\Mux7~2_combout  & ((\Reg[30][24]~q ))) # (!\Mux7~2_combout  & (\Reg[26][24]~q )))) # (!ifid_ifinstr_o_24 & (\Mux7~2_combout ))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux7~2_combout ),
	.datac(\Reg[26][24]~q ),
	.datad(\Reg[30][24]~q ),
	.cin(gnd),
	.combout(\Mux7~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~3 .lut_mask = 16'hEC64;
defparam \Mux7~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y32_N31
dffeas \Reg[16][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][24] .is_wysiwyg = "true";
defparam \Reg[16][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N20
cycloneive_lcell_comb \Mux7~4 (
// Equation(s):
// \Mux7~4_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & (\Reg[20][24]~q )) # (!ifid_ifinstr_o_23 & ((\Reg[16][24]~q )))))

	.dataa(\Reg[20][24]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[16][24]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux7~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~4 .lut_mask = 16'hEE30;
defparam \Mux7~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y32_N1
dffeas \Reg[24][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][24] .is_wysiwyg = "true";
defparam \Reg[24][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N0
cycloneive_lcell_comb \Mux7~5 (
// Equation(s):
// \Mux7~5_combout  = (\Mux7~4_combout  & ((\Reg[28][24]~q ) # ((!ifid_ifinstr_o_24)))) # (!\Mux7~4_combout  & (((\Reg[24][24]~q  & ifid_ifinstr_o_24))))

	.dataa(\Reg[28][24]~q ),
	.datab(\Mux7~4_combout ),
	.datac(\Reg[24][24]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux7~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~5 .lut_mask = 16'hB8CC;
defparam \Mux7~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N26
cycloneive_lcell_comb \Mux7~6 (
// Equation(s):
// \Mux7~6_combout  = (ifid_ifinstr_o_21 & (ifid_ifinstr_o_22)) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Mux7~3_combout )) # (!ifid_ifinstr_o_22 & ((\Mux7~5_combout )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Mux7~3_combout ),
	.datad(\Mux7~5_combout ),
	.cin(gnd),
	.combout(\Mux7~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~6 .lut_mask = 16'hD9C8;
defparam \Mux7~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N15
dffeas \Reg[21][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][24] .is_wysiwyg = "true";
defparam \Reg[21][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N1
dffeas \Reg[29][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][24] .is_wysiwyg = "true";
defparam \Reg[29][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N7
dffeas \Reg[25][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][24] .is_wysiwyg = "true";
defparam \Reg[25][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N29
dffeas \Reg[17][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][24] .is_wysiwyg = "true";
defparam \Reg[17][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N28
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (ifid_ifinstr_o_24 & ((\Reg[25][24]~q ) # ((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & (((\Reg[17][24]~q  & !ifid_ifinstr_o_23))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[25][24]~q ),
	.datac(\Reg[17][24]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hAAD8;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N0
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// \Mux7~1_combout  = (ifid_ifinstr_o_23 & ((\Mux7~0_combout  & ((\Reg[29][24]~q ))) # (!\Mux7~0_combout  & (\Reg[21][24]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux7~0_combout ))))

	.dataa(\Reg[21][24]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[29][24]~q ),
	.datad(\Mux7~0_combout ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hF388;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N11
dffeas \Reg[31][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][24] .is_wysiwyg = "true";
defparam \Reg[31][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N29
dffeas \Reg[27][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][24] .is_wysiwyg = "true";
defparam \Reg[27][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N3
dffeas \Reg[19][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][24] .is_wysiwyg = "true";
defparam \Reg[19][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N28
cycloneive_lcell_comb \Mux7~7 (
// Equation(s):
// \Mux7~7_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[27][24]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[19][24]~q )))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[27][24]~q ),
	.datad(\Reg[19][24]~q ),
	.cin(gnd),
	.combout(\Mux7~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~7 .lut_mask = 16'hD9C8;
defparam \Mux7~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N25
dffeas \Reg[23][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][24] .is_wysiwyg = "true";
defparam \Reg[23][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N24
cycloneive_lcell_comb \Mux7~8 (
// Equation(s):
// \Mux7~8_combout  = (\Mux7~7_combout  & ((\Reg[31][24]~q ) # ((!ifid_ifinstr_o_23)))) # (!\Mux7~7_combout  & (((\Reg[23][24]~q  & ifid_ifinstr_o_23))))

	.dataa(\Reg[31][24]~q ),
	.datab(\Mux7~7_combout ),
	.datac(\Reg[23][24]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux7~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~8 .lut_mask = 16'hB8CC;
defparam \Mux7~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y39_N21
dffeas \Reg[5][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][24] .is_wysiwyg = "true";
defparam \Reg[5][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N20
cycloneive_lcell_comb \Mux7~10 (
// Equation(s):
// \Mux7~10_combout  = (ifid_ifinstr_o_21 & (((\Reg[5][24]~q ) # (ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & (\Reg[4][24]~q  & ((!ifid_ifinstr_o_22))))

	.dataa(\Reg[4][24]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[5][24]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux7~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~10 .lut_mask = 16'hCCE2;
defparam \Mux7~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N27
dffeas \Reg[6][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][24] .is_wysiwyg = "true";
defparam \Reg[6][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N16
cycloneive_lcell_comb \Reg[7][24]~feeder (
// Equation(s):
// \Reg[7][24]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat24),
	.cin(gnd),
	.combout(\Reg[7][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[7][24]~feeder .lut_mask = 16'hFF00;
defparam \Reg[7][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N17
dffeas \Reg[7][24] (
	.clk(!CLK),
	.d(\Reg[7][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][24] .is_wysiwyg = "true";
defparam \Reg[7][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N26
cycloneive_lcell_comb \Mux7~11 (
// Equation(s):
// \Mux7~11_combout  = (\Mux7~10_combout  & (((\Reg[7][24]~q )) # (!ifid_ifinstr_o_22))) # (!\Mux7~10_combout  & (ifid_ifinstr_o_22 & (\Reg[6][24]~q )))

	.dataa(\Mux7~10_combout ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[6][24]~q ),
	.datad(\Reg[7][24]~q ),
	.cin(gnd),
	.combout(\Mux7~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~11 .lut_mask = 16'hEA62;
defparam \Mux7~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y37_N31
dffeas \Reg[14][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][24] .is_wysiwyg = "true";
defparam \Reg[14][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y37_N5
dffeas \Reg[15][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][24] .is_wysiwyg = "true";
defparam \Reg[15][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y37_N19
dffeas \Reg[12][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][24] .is_wysiwyg = "true";
defparam \Reg[12][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y37_N21
dffeas \Reg[13][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][24] .is_wysiwyg = "true";
defparam \Reg[13][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y37_N18
cycloneive_lcell_comb \Mux7~17 (
// Equation(s):
// \Mux7~17_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[13][24]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[12][24]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[12][24]~q ),
	.datad(\Reg[13][24]~q ),
	.cin(gnd),
	.combout(\Mux7~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~17 .lut_mask = 16'hDC98;
defparam \Mux7~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N4
cycloneive_lcell_comb \Mux7~18 (
// Equation(s):
// \Mux7~18_combout  = (ifid_ifinstr_o_22 & ((\Mux7~17_combout  & ((\Reg[15][24]~q ))) # (!\Mux7~17_combout  & (\Reg[14][24]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux7~17_combout ))))

	.dataa(\Reg[14][24]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[15][24]~q ),
	.datad(\Mux7~17_combout ),
	.cin(gnd),
	.combout(\Mux7~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~18 .lut_mask = 16'hF388;
defparam \Mux7~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N27
dffeas \Reg[1][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][24] .is_wysiwyg = "true";
defparam \Reg[1][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N22
cycloneive_lcell_comb \Mux7~14 (
// Equation(s):
// \Mux7~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[3][24]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[1][24]~q )))))

	.dataa(\Reg[3][24]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(ifid_ifinstr_o_22),
	.datad(\Reg[1][24]~q ),
	.cin(gnd),
	.combout(\Mux7~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~14 .lut_mask = 16'h8C80;
defparam \Mux7~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N22
cycloneive_lcell_comb \Reg[2][24]~feeder (
// Equation(s):
// \Reg[2][24]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat24),
	.cin(gnd),
	.combout(\Reg[2][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[2][24]~feeder .lut_mask = 16'hFF00;
defparam \Reg[2][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N23
dffeas \Reg[2][24] (
	.clk(!CLK),
	.d(\Reg[2][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][24] .is_wysiwyg = "true";
defparam \Reg[2][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N20
cycloneive_lcell_comb \Mux7~15 (
// Equation(s):
// \Mux7~15_combout  = (\Mux7~14_combout ) # ((ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & \Reg[2][24]~q )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux7~14_combout ),
	.datad(\Reg[2][24]~q ),
	.cin(gnd),
	.combout(\Mux7~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~15 .lut_mask = 16'hF2F0;
defparam \Mux7~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y32_N29
dffeas \Reg[10][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][24] .is_wysiwyg = "true";
defparam \Reg[10][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N11
dffeas \Reg[8][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][24] .is_wysiwyg = "true";
defparam \Reg[8][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N10
cycloneive_lcell_comb \Mux7~12 (
// Equation(s):
// \Mux7~12_combout  = (ifid_ifinstr_o_22 & ((\Reg[10][24]~q ) # ((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & (((\Reg[8][24]~q  & !ifid_ifinstr_o_21))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[10][24]~q ),
	.datac(\Reg[8][24]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux7~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~12 .lut_mask = 16'hAAD8;
defparam \Mux7~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N19
dffeas \Reg[11][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][24] .is_wysiwyg = "true";
defparam \Reg[11][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N18
cycloneive_lcell_comb \Mux7~13 (
// Equation(s):
// \Mux7~13_combout  = (\Mux7~12_combout  & (((\Reg[11][24]~q ) # (!ifid_ifinstr_o_21)))) # (!\Mux7~12_combout  & (\Reg[9][24]~q  & ((ifid_ifinstr_o_21))))

	.dataa(\Reg[9][24]~q ),
	.datab(\Mux7~12_combout ),
	.datac(\Reg[11][24]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux7~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~13 .lut_mask = 16'hE2CC;
defparam \Mux7~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N10
cycloneive_lcell_comb \Mux7~16 (
// Equation(s):
// \Mux7~16_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Mux7~13_combout ))) # (!ifid_ifinstr_o_24 & (\Mux7~15_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Mux7~15_combout ),
	.datad(\Mux7~13_combout ),
	.cin(gnd),
	.combout(\Mux7~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~16 .lut_mask = 16'hDC98;
defparam \Mux7~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N11
dffeas \Reg[31][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][22] .is_wysiwyg = "true";
defparam \Reg[31][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N21
dffeas \Reg[23][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][22] .is_wysiwyg = "true";
defparam \Reg[23][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N29
dffeas \Reg[27][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][22] .is_wysiwyg = "true";
defparam \Reg[27][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N15
dffeas \Reg[19][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][22] .is_wysiwyg = "true";
defparam \Reg[19][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N28
cycloneive_lcell_comb \Mux9~7 (
// Equation(s):
// \Mux9~7_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[27][22]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[19][22]~q )))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[27][22]~q ),
	.datad(\Reg[19][22]~q ),
	.cin(gnd),
	.combout(\Mux9~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~7 .lut_mask = 16'hD9C8;
defparam \Mux9~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N20
cycloneive_lcell_comb \Mux9~8 (
// Equation(s):
// \Mux9~8_combout  = (ifid_ifinstr_o_23 & ((\Mux9~7_combout  & (\Reg[31][22]~q )) # (!\Mux9~7_combout  & ((\Reg[23][22]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux9~7_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[31][22]~q ),
	.datac(\Reg[23][22]~q ),
	.datad(\Mux9~7_combout ),
	.cin(gnd),
	.combout(\Mux9~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~8 .lut_mask = 16'hDDA0;
defparam \Mux9~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y32_N15
dffeas \Reg[16][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][22] .is_wysiwyg = "true";
defparam \Reg[16][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N14
cycloneive_lcell_comb \Mux9~4 (
// Equation(s):
// \Mux9~4_combout  = (ifid_ifinstr_o_23 & ((\Reg[20][22]~q ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((\Reg[16][22]~q  & !ifid_ifinstr_o_24))))

	.dataa(\Reg[20][22]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[16][22]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux9~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~4 .lut_mask = 16'hCCB8;
defparam \Mux9~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N9
dffeas \Reg[28][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][22] .is_wysiwyg = "true";
defparam \Reg[28][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y32_N17
dffeas \Reg[24][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][22] .is_wysiwyg = "true";
defparam \Reg[24][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N12
cycloneive_lcell_comb \Mux9~5 (
// Equation(s):
// \Mux9~5_combout  = (ifid_ifinstr_o_24 & ((\Mux9~4_combout  & (\Reg[28][22]~q )) # (!\Mux9~4_combout  & ((\Reg[24][22]~q ))))) # (!ifid_ifinstr_o_24 & (\Mux9~4_combout ))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux9~4_combout ),
	.datac(\Reg[28][22]~q ),
	.datad(\Reg[24][22]~q ),
	.cin(gnd),
	.combout(\Mux9~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~5 .lut_mask = 16'hE6C4;
defparam \Mux9~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N20
cycloneive_lcell_comb \Reg[30][22]~feeder (
// Equation(s):
// \Reg[30][22]~feeder_combout  = \wdat~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat25),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[30][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[30][22]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[30][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y36_N21
dffeas \Reg[30][22] (
	.clk(!CLK),
	.d(\Reg[30][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][22] .is_wysiwyg = "true";
defparam \Reg[30][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N29
dffeas \Reg[18][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][22] .is_wysiwyg = "true";
defparam \Reg[18][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y36_N3
dffeas \Reg[22][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][22] .is_wysiwyg = "true";
defparam \Reg[22][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N28
cycloneive_lcell_comb \Mux9~2 (
// Equation(s):
// \Mux9~2_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[22][22]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[18][22]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[18][22]~q ),
	.datad(\Reg[22][22]~q ),
	.cin(gnd),
	.combout(\Mux9~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~2 .lut_mask = 16'hDC98;
defparam \Mux9~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N23
dffeas \Reg[26][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][22] .is_wysiwyg = "true";
defparam \Reg[26][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N10
cycloneive_lcell_comb \Mux9~3 (
// Equation(s):
// \Mux9~3_combout  = (ifid_ifinstr_o_24 & ((\Mux9~2_combout  & (\Reg[30][22]~q )) # (!\Mux9~2_combout  & ((\Reg[26][22]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux9~2_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[30][22]~q ),
	.datac(\Mux9~2_combout ),
	.datad(\Reg[26][22]~q ),
	.cin(gnd),
	.combout(\Mux9~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~3 .lut_mask = 16'hDAD0;
defparam \Mux9~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N22
cycloneive_lcell_comb \Mux9~6 (
// Equation(s):
// \Mux9~6_combout  = (ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21) # ((\Mux9~3_combout )))) # (!ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & (\Mux9~5_combout )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux9~5_combout ),
	.datad(\Mux9~3_combout ),
	.cin(gnd),
	.combout(\Mux9~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~6 .lut_mask = 16'hBA98;
defparam \Mux9~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N17
dffeas \Reg[21][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][22] .is_wysiwyg = "true";
defparam \Reg[21][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y38_N13
dffeas \Reg[29][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][22] .is_wysiwyg = "true";
defparam \Reg[29][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N4
cycloneive_lcell_comb \Reg[17][22]~feeder (
// Equation(s):
// \Reg[17][22]~feeder_combout  = \wdat~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat25),
	.cin(gnd),
	.combout(\Reg[17][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[17][22]~feeder .lut_mask = 16'hFF00;
defparam \Reg[17][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N5
dffeas \Reg[17][22] (
	.clk(!CLK),
	.d(\Reg[17][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][22] .is_wysiwyg = "true";
defparam \Reg[17][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N10
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// \Mux9~0_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[25][22]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[17][22]~q )))))

	.dataa(\Reg[25][22]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[17][22]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hEE30;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N12
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// \Mux9~1_combout  = (ifid_ifinstr_o_23 & ((\Mux9~0_combout  & ((\Reg[29][22]~q ))) # (!\Mux9~0_combout  & (\Reg[21][22]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux9~0_combout ))))

	.dataa(\Reg[21][22]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[29][22]~q ),
	.datad(\Mux9~0_combout ),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'hF388;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y37_N23
dffeas \Reg[12][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][22] .is_wysiwyg = "true";
defparam \Reg[12][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y37_N29
dffeas \Reg[13][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][22] .is_wysiwyg = "true";
defparam \Reg[13][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y37_N22
cycloneive_lcell_comb \Mux9~17 (
// Equation(s):
// \Mux9~17_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[13][22]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[12][22]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[12][22]~q ),
	.datad(\Reg[13][22]~q ),
	.cin(gnd),
	.combout(\Mux9~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~17 .lut_mask = 16'hDC98;
defparam \Mux9~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y37_N21
dffeas \Reg[15][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][22] .is_wysiwyg = "true";
defparam \Reg[15][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y37_N11
dffeas \Reg[14][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][22] .is_wysiwyg = "true";
defparam \Reg[14][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N20
cycloneive_lcell_comb \Mux9~18 (
// Equation(s):
// \Mux9~18_combout  = (ifid_ifinstr_o_22 & ((\Mux9~17_combout  & (\Reg[15][22]~q )) # (!\Mux9~17_combout  & ((\Reg[14][22]~q ))))) # (!ifid_ifinstr_o_22 & (\Mux9~17_combout ))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Mux9~17_combout ),
	.datac(\Reg[15][22]~q ),
	.datad(\Reg[14][22]~q ),
	.cin(gnd),
	.combout(\Mux9~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~18 .lut_mask = 16'hE6C4;
defparam \Mux9~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N30
cycloneive_lcell_comb \Reg[1][22]~feeder (
// Equation(s):
// \Reg[1][22]~feeder_combout  = \wdat~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat25),
	.cin(gnd),
	.combout(\Reg[1][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[1][22]~feeder .lut_mask = 16'hFF00;
defparam \Reg[1][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y35_N31
dffeas \Reg[1][22] (
	.clk(!CLK),
	.d(\Reg[1][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][22] .is_wysiwyg = "true";
defparam \Reg[1][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N13
dffeas \Reg[3][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][22] .is_wysiwyg = "true";
defparam \Reg[3][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N28
cycloneive_lcell_comb \Mux9~14 (
// Equation(s):
// \Mux9~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][22]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][22]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[1][22]~q ),
	.datad(\Reg[3][22]~q ),
	.cin(gnd),
	.combout(\Mux9~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~14 .lut_mask = 16'hC840;
defparam \Mux9~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y31_N17
dffeas \Reg[2][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][22] .is_wysiwyg = "true";
defparam \Reg[2][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N16
cycloneive_lcell_comb \Mux9~15 (
// Equation(s):
// \Mux9~15_combout  = (\Mux9~14_combout ) # ((ifid_ifinstr_o_22 & (\Reg[2][22]~q  & !ifid_ifinstr_o_21)))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Mux9~14_combout ),
	.datac(\Reg[2][22]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux9~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~15 .lut_mask = 16'hCCEC;
defparam \Mux9~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y31_N23
dffeas \Reg[11][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][22] .is_wysiwyg = "true";
defparam \Reg[11][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N5
dffeas \Reg[10][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][22] .is_wysiwyg = "true";
defparam \Reg[10][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N31
dffeas \Reg[8][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][22] .is_wysiwyg = "true";
defparam \Reg[8][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N30
cycloneive_lcell_comb \Mux9~12 (
// Equation(s):
// \Mux9~12_combout  = (ifid_ifinstr_o_22 & ((\Reg[10][22]~q ) # ((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & (((\Reg[8][22]~q  & !ifid_ifinstr_o_21))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[10][22]~q ),
	.datac(\Reg[8][22]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux9~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~12 .lut_mask = 16'hAAD8;
defparam \Mux9~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N22
cycloneive_lcell_comb \Mux9~13 (
// Equation(s):
// \Mux9~13_combout  = (ifid_ifinstr_o_21 & ((\Mux9~12_combout  & ((\Reg[11][22]~q ))) # (!\Mux9~12_combout  & (\Reg[9][22]~q )))) # (!ifid_ifinstr_o_21 & (((\Mux9~12_combout ))))

	.dataa(\Reg[9][22]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[11][22]~q ),
	.datad(\Mux9~12_combout ),
	.cin(gnd),
	.combout(\Mux9~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~13 .lut_mask = 16'hF388;
defparam \Mux9~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N18
cycloneive_lcell_comb \Mux9~16 (
// Equation(s):
// \Mux9~16_combout  = (ifid_ifinstr_o_24 & (((\Mux9~13_combout ) # (ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & (\Mux9~15_combout  & ((!ifid_ifinstr_o_23))))

	.dataa(\Mux9~15_combout ),
	.datab(\Mux9~13_combout ),
	.datac(ifid_ifinstr_o_24),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux9~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~16 .lut_mask = 16'hF0CA;
defparam \Mux9~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y39_N31
dffeas \Reg[7][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][22] .is_wysiwyg = "true";
defparam \Reg[7][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y39_N15
dffeas \Reg[4][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][22] .is_wysiwyg = "true";
defparam \Reg[4][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y39_N25
dffeas \Reg[5][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][22] .is_wysiwyg = "true";
defparam \Reg[5][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N24
cycloneive_lcell_comb \Mux9~10 (
// Equation(s):
// \Mux9~10_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[5][22]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[4][22]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[4][22]~q ),
	.datac(\Reg[5][22]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux9~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~10 .lut_mask = 16'hFA44;
defparam \Mux9~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y39_N21
dffeas \Reg[6][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][22] .is_wysiwyg = "true";
defparam \Reg[6][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N20
cycloneive_lcell_comb \Mux9~11 (
// Equation(s):
// \Mux9~11_combout  = (\Mux9~10_combout  & ((\Reg[7][22]~q ) # ((!ifid_ifinstr_o_22)))) # (!\Mux9~10_combout  & (((\Reg[6][22]~q  & ifid_ifinstr_o_22))))

	.dataa(\Reg[7][22]~q ),
	.datab(\Mux9~10_combout ),
	.datac(\Reg[6][22]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux9~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~11 .lut_mask = 16'hB8CC;
defparam \Mux9~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N27
dffeas \Reg[19][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][23] .is_wysiwyg = "true";
defparam \Reg[19][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y29_N21
dffeas \Reg[23][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][23] .is_wysiwyg = "true";
defparam \Reg[23][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N20
cycloneive_lcell_comb \Mux8~7 (
// Equation(s):
// \Mux8~7_combout  = (ifid_ifinstr_o_23 & (((\Reg[23][23]~q ) # (ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (\Reg[19][23]~q  & ((!ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[19][23]~q ),
	.datac(\Reg[23][23]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux8~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~7 .lut_mask = 16'hAAE4;
defparam \Mux8~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N13
dffeas \Reg[27][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][23] .is_wysiwyg = "true";
defparam \Reg[27][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y29_N23
dffeas \Reg[31][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][23] .is_wysiwyg = "true";
defparam \Reg[31][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N12
cycloneive_lcell_comb \Mux8~8 (
// Equation(s):
// \Mux8~8_combout  = (ifid_ifinstr_o_24 & ((\Mux8~7_combout  & ((\Reg[31][23]~q ))) # (!\Mux8~7_combout  & (\Reg[27][23]~q )))) # (!ifid_ifinstr_o_24 & (\Mux8~7_combout ))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux8~7_combout ),
	.datac(\Reg[27][23]~q ),
	.datad(\Reg[31][23]~q ),
	.cin(gnd),
	.combout(\Mux8~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~8 .lut_mask = 16'hEC64;
defparam \Mux8~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N26
cycloneive_lcell_comb \Reg[29][23]~feeder (
// Equation(s):
// \Reg[29][23]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat26),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[29][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[29][23]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[29][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N27
dffeas \Reg[29][23] (
	.clk(!CLK),
	.d(\Reg[29][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][23] .is_wysiwyg = "true";
defparam \Reg[29][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N22
cycloneive_lcell_comb \Reg[17][23]~feeder (
// Equation(s):
// \Reg[17][23]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat26),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[17][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[17][23]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[17][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N23
dffeas \Reg[17][23] (
	.clk(!CLK),
	.d(\Reg[17][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][23] .is_wysiwyg = "true";
defparam \Reg[17][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N20
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// \Mux8~0_combout  = (ifid_ifinstr_o_23 & ((\Reg[21][23]~q ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((\Reg[17][23]~q  & !ifid_ifinstr_o_24))))

	.dataa(\Reg[21][23]~q ),
	.datab(\Reg[17][23]~q ),
	.datac(ifid_ifinstr_o_23),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hF0AC;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N16
cycloneive_lcell_comb \Reg[25][23]~feeder (
// Equation(s):
// \Reg[25][23]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat26),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[25][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][23]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[25][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N17
dffeas \Reg[25][23] (
	.clk(!CLK),
	.d(\Reg[25][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][23] .is_wysiwyg = "true";
defparam \Reg[25][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N28
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// \Mux8~1_combout  = (\Mux8~0_combout  & ((\Reg[29][23]~q ) # ((!ifid_ifinstr_o_24)))) # (!\Mux8~0_combout  & (((\Reg[25][23]~q  & ifid_ifinstr_o_24))))

	.dataa(\Reg[29][23]~q ),
	.datab(\Mux8~0_combout ),
	.datac(\Reg[25][23]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'hB8CC;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N29
dffeas \Reg[22][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][23] .is_wysiwyg = "true";
defparam \Reg[22][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N29
dffeas \Reg[26][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][23] .is_wysiwyg = "true";
defparam \Reg[26][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N7
dffeas \Reg[18][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][23] .is_wysiwyg = "true";
defparam \Reg[18][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N28
cycloneive_lcell_comb \Mux8~2 (
// Equation(s):
// \Mux8~2_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[26][23]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[18][23]~q )))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[26][23]~q ),
	.datad(\Reg[18][23]~q ),
	.cin(gnd),
	.combout(\Mux8~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~2 .lut_mask = 16'hD9C8;
defparam \Mux8~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N28
cycloneive_lcell_comb \Mux8~3 (
// Equation(s):
// \Mux8~3_combout  = (ifid_ifinstr_o_23 & ((\Mux8~2_combout  & (\Reg[30][23]~q )) # (!\Mux8~2_combout  & ((\Reg[22][23]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux8~2_combout ))))

	.dataa(\Reg[30][23]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[22][23]~q ),
	.datad(\Mux8~2_combout ),
	.cin(gnd),
	.combout(\Mux8~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~3 .lut_mask = 16'hBBC0;
defparam \Mux8~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N7
dffeas \Reg[28][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][23] .is_wysiwyg = "true";
defparam \Reg[28][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y33_N11
dffeas \Reg[16][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][23] .is_wysiwyg = "true";
defparam \Reg[16][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N24
cycloneive_lcell_comb \Reg[24][23]~feeder (
// Equation(s):
// \Reg[24][23]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat26),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[24][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[24][23]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[24][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N25
dffeas \Reg[24][23] (
	.clk(!CLK),
	.d(\Reg[24][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][23] .is_wysiwyg = "true";
defparam \Reg[24][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N10
cycloneive_lcell_comb \Mux8~4 (
// Equation(s):
// \Mux8~4_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Reg[24][23]~q ))) # (!ifid_ifinstr_o_24 & (\Reg[16][23]~q ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[16][23]~q ),
	.datad(\Reg[24][23]~q ),
	.cin(gnd),
	.combout(\Mux8~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~4 .lut_mask = 16'hDC98;
defparam \Mux8~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y33_N21
dffeas \Reg[20][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][23] .is_wysiwyg = "true";
defparam \Reg[20][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N16
cycloneive_lcell_comb \Mux8~5 (
// Equation(s):
// \Mux8~5_combout  = (ifid_ifinstr_o_23 & ((\Mux8~4_combout  & (\Reg[28][23]~q )) # (!\Mux8~4_combout  & ((\Reg[20][23]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux8~4_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[28][23]~q ),
	.datac(\Mux8~4_combout ),
	.datad(\Reg[20][23]~q ),
	.cin(gnd),
	.combout(\Mux8~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~5 .lut_mask = 16'hDAD0;
defparam \Mux8~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N12
cycloneive_lcell_comb \Mux8~6 (
// Equation(s):
// \Mux8~6_combout  = (ifid_ifinstr_o_22 & ((\Mux8~3_combout ) # ((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & (((\Mux8~5_combout  & !ifid_ifinstr_o_21))))

	.dataa(\Mux8~3_combout ),
	.datab(\Mux8~5_combout ),
	.datac(ifid_ifinstr_o_22),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux8~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~6 .lut_mask = 16'hF0AC;
defparam \Mux8~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N24
cycloneive_lcell_comb \Reg[15][23]~feeder (
// Equation(s):
// \Reg[15][23]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat26),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[15][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[15][23]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[15][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N25
dffeas \Reg[15][23] (
	.clk(!CLK),
	.d(\Reg[15][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][23] .is_wysiwyg = "true";
defparam \Reg[15][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y37_N7
dffeas \Reg[14][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][23] .is_wysiwyg = "true";
defparam \Reg[14][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y37_N5
dffeas \Reg[13][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][23] .is_wysiwyg = "true";
defparam \Reg[13][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y37_N27
dffeas \Reg[12][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][23] .is_wysiwyg = "true";
defparam \Reg[12][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y37_N26
cycloneive_lcell_comb \Mux8~17 (
// Equation(s):
// \Mux8~17_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[13][23]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[12][23]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[13][23]~q ),
	.datac(\Reg[12][23]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux8~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~17 .lut_mask = 16'hEE50;
defparam \Mux8~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N6
cycloneive_lcell_comb \Mux8~18 (
// Equation(s):
// \Mux8~18_combout  = (ifid_ifinstr_o_22 & ((\Mux8~17_combout  & (\Reg[15][23]~q )) # (!\Mux8~17_combout  & ((\Reg[14][23]~q ))))) # (!ifid_ifinstr_o_22 & (((\Mux8~17_combout ))))

	.dataa(\Reg[15][23]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[14][23]~q ),
	.datad(\Mux8~17_combout ),
	.cin(gnd),
	.combout(\Mux8~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~18 .lut_mask = 16'hBBC0;
defparam \Mux8~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y35_N9
dffeas \Reg[1][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][23] .is_wysiwyg = "true";
defparam \Reg[1][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N8
cycloneive_lcell_comb \Mux8~14 (
// Equation(s):
// \Mux8~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[3][23]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[1][23]~q )))))

	.dataa(\Reg[3][23]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[1][23]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux8~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~14 .lut_mask = 16'h88C0;
defparam \Mux8~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N4
cycloneive_lcell_comb \Mux8~15 (
// Equation(s):
// \Mux8~15_combout  = (\Mux8~14_combout ) # ((\Reg[2][23]~q  & (!ifid_ifinstr_o_21 & ifid_ifinstr_o_22)))

	.dataa(\Reg[2][23]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(ifid_ifinstr_o_22),
	.datad(\Mux8~14_combout ),
	.cin(gnd),
	.combout(\Mux8~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~15 .lut_mask = 16'hFF20;
defparam \Mux8~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N8
cycloneive_lcell_comb \Reg[6][23]~feeder (
// Equation(s):
// \Reg[6][23]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat26),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[6][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[6][23]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[6][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N9
dffeas \Reg[6][23] (
	.clk(!CLK),
	.d(\Reg[6][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][23] .is_wysiwyg = "true";
defparam \Reg[6][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N25
dffeas \Reg[7][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][23] .is_wysiwyg = "true";
defparam \Reg[7][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y39_N9
dffeas \Reg[5][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][23] .is_wysiwyg = "true";
defparam \Reg[5][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y39_N11
dffeas \Reg[4][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][23] .is_wysiwyg = "true";
defparam \Reg[4][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N10
cycloneive_lcell_comb \Mux8~12 (
// Equation(s):
// \Mux8~12_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[5][23]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[4][23]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[5][23]~q ),
	.datac(\Reg[4][23]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux8~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~12 .lut_mask = 16'hEE50;
defparam \Mux8~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N24
cycloneive_lcell_comb \Mux8~13 (
// Equation(s):
// \Mux8~13_combout  = (ifid_ifinstr_o_22 & ((\Mux8~12_combout  & ((\Reg[7][23]~q ))) # (!\Mux8~12_combout  & (\Reg[6][23]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux8~12_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[6][23]~q ),
	.datac(\Reg[7][23]~q ),
	.datad(\Mux8~12_combout ),
	.cin(gnd),
	.combout(\Mux8~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~13 .lut_mask = 16'hF588;
defparam \Mux8~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N20
cycloneive_lcell_comb \Mux8~16 (
// Equation(s):
// \Mux8~16_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Mux8~13_combout ))) # (!ifid_ifinstr_o_23 & (\Mux8~15_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux8~15_combout ),
	.datac(\Mux8~13_combout ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux8~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~16 .lut_mask = 16'hFA44;
defparam \Mux8~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N27
dffeas \Reg[11][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][23] .is_wysiwyg = "true";
defparam \Reg[11][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y33_N1
dffeas \Reg[9][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][23] .is_wysiwyg = "true";
defparam \Reg[9][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N1
dffeas \Reg[10][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][23] .is_wysiwyg = "true";
defparam \Reg[10][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N0
cycloneive_lcell_comb \Mux8~10 (
// Equation(s):
// \Mux8~10_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[10][23]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[8][23]~q ))))

	.dataa(\Reg[8][23]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[10][23]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux8~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~10 .lut_mask = 16'hFC22;
defparam \Mux8~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N0
cycloneive_lcell_comb \Mux8~11 (
// Equation(s):
// \Mux8~11_combout  = (ifid_ifinstr_o_21 & ((\Mux8~10_combout  & (\Reg[11][23]~q )) # (!\Mux8~10_combout  & ((\Reg[9][23]~q ))))) # (!ifid_ifinstr_o_21 & (((\Mux8~10_combout ))))

	.dataa(\Reg[11][23]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[9][23]~q ),
	.datad(\Mux8~10_combout ),
	.cin(gnd),
	.combout(\Mux8~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~11 .lut_mask = 16'hBBC0;
defparam \Mux8~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N11
dffeas \Reg[28][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][21] .is_wysiwyg = "true";
defparam \Reg[28][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y33_N25
dffeas \Reg[16][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][21] .is_wysiwyg = "true";
defparam \Reg[16][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N24
cycloneive_lcell_comb \Mux10~4 (
// Equation(s):
// \Mux10~4_combout  = (ifid_ifinstr_o_24 & ((\Reg[24][21]~q ) # ((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & (((\Reg[16][21]~q  & !ifid_ifinstr_o_23))))

	.dataa(\Reg[24][21]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[16][21]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~4 .lut_mask = 16'hCCB8;
defparam \Mux10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N10
cycloneive_lcell_comb \Mux10~5 (
// Equation(s):
// \Mux10~5_combout  = (ifid_ifinstr_o_23 & ((\Mux10~4_combout  & ((\Reg[28][21]~q ))) # (!\Mux10~4_combout  & (\Reg[20][21]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux10~4_combout ))))

	.dataa(\Reg[20][21]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[28][21]~q ),
	.datad(\Mux10~4_combout ),
	.cin(gnd),
	.combout(\Mux10~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~5 .lut_mask = 16'hF388;
defparam \Mux10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N21
dffeas \Reg[18][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][21] .is_wysiwyg = "true";
defparam \Reg[18][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N20
cycloneive_lcell_comb \Mux10~2 (
// Equation(s):
// \Mux10~2_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[26][21]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[18][21]~q )))))

	.dataa(\Reg[26][21]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[18][21]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~2 .lut_mask = 16'hEE30;
defparam \Mux10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N1
dffeas \Reg[22][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][21] .is_wysiwyg = "true";
defparam \Reg[22][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N0
cycloneive_lcell_comb \Mux10~3 (
// Equation(s):
// \Mux10~3_combout  = (ifid_ifinstr_o_23 & ((\Mux10~2_combout  & (\Reg[30][21]~q )) # (!\Mux10~2_combout  & ((\Reg[22][21]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux10~2_combout ))))

	.dataa(\Reg[30][21]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Mux10~2_combout ),
	.datad(\Reg[22][21]~q ),
	.cin(gnd),
	.combout(\Mux10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~3 .lut_mask = 16'hBCB0;
defparam \Mux10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N26
cycloneive_lcell_comb \Mux10~6 (
// Equation(s):
// \Mux10~6_combout  = (ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21) # ((\Mux10~3_combout )))) # (!ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & (\Mux10~5_combout )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux10~5_combout ),
	.datad(\Mux10~3_combout ),
	.cin(gnd),
	.combout(\Mux10~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~6 .lut_mask = 16'hBA98;
defparam \Mux10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N25
dffeas \Reg[27][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][21] .is_wysiwyg = "true";
defparam \Reg[27][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N3
dffeas \Reg[31][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][21] .is_wysiwyg = "true";
defparam \Reg[31][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N14
cycloneive_lcell_comb \Reg[23][21]~feeder (
// Equation(s):
// \Reg[23][21]~feeder_combout  = \wdat~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat27),
	.cin(gnd),
	.combout(\Reg[23][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[23][21]~feeder .lut_mask = 16'hFF00;
defparam \Reg[23][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N15
dffeas \Reg[23][21] (
	.clk(!CLK),
	.d(\Reg[23][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][21] .is_wysiwyg = "true";
defparam \Reg[23][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N5
dffeas \Reg[19][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][21] .is_wysiwyg = "true";
defparam \Reg[19][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N4
cycloneive_lcell_comb \Mux10~7 (
// Equation(s):
// \Mux10~7_combout  = (ifid_ifinstr_o_23 & ((\Reg[23][21]~q ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((\Reg[19][21]~q  & !ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[23][21]~q ),
	.datac(\Reg[19][21]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux10~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~7 .lut_mask = 16'hAAD8;
defparam \Mux10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N26
cycloneive_lcell_comb \Mux10~8 (
// Equation(s):
// \Mux10~8_combout  = (\Mux10~7_combout  & (((\Reg[31][21]~q ) # (!ifid_ifinstr_o_24)))) # (!\Mux10~7_combout  & (\Reg[27][21]~q  & ((ifid_ifinstr_o_24))))

	.dataa(\Reg[27][21]~q ),
	.datab(\Reg[31][21]~q ),
	.datac(\Mux10~7_combout ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux10~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~8 .lut_mask = 16'hCAF0;
defparam \Mux10~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N15
dffeas \Reg[17][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][21] .is_wysiwyg = "true";
defparam \Reg[17][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y37_N5
dffeas \Reg[21][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][21] .is_wysiwyg = "true";
defparam \Reg[21][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N14
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// \Mux10~0_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[21][21]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[17][21]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[17][21]~q ),
	.datad(\Reg[21][21]~q ),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hDC98;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y37_N19
dffeas \Reg[29][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][21] .is_wysiwyg = "true";
defparam \Reg[29][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N13
dffeas \Reg[25][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][21] .is_wysiwyg = "true";
defparam \Reg[25][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N18
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// \Mux10~1_combout  = (ifid_ifinstr_o_24 & ((\Mux10~0_combout  & (\Reg[29][21]~q )) # (!\Mux10~0_combout  & ((\Reg[25][21]~q ))))) # (!ifid_ifinstr_o_24 & (\Mux10~0_combout ))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux10~0_combout ),
	.datac(\Reg[29][21]~q ),
	.datad(\Reg[25][21]~q ),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'hE6C4;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y37_N25
dffeas \Reg[13][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][21] .is_wysiwyg = "true";
defparam \Reg[13][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y37_N3
dffeas \Reg[12][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][21] .is_wysiwyg = "true";
defparam \Reg[12][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y37_N24
cycloneive_lcell_comb \Mux10~17 (
// Equation(s):
// \Mux10~17_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[13][21]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[12][21]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[13][21]~q ),
	.datad(\Reg[12][21]~q ),
	.cin(gnd),
	.combout(\Mux10~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~17 .lut_mask = 16'hD9C8;
defparam \Mux10~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y37_N17
dffeas \Reg[14][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][21] .is_wysiwyg = "true";
defparam \Reg[14][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N8
cycloneive_lcell_comb \Reg[15][21]~feeder (
// Equation(s):
// \Reg[15][21]~feeder_combout  = \wdat~57_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat27),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[15][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[15][21]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[15][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y37_N9
dffeas \Reg[15][21] (
	.clk(!CLK),
	.d(\Reg[15][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][21] .is_wysiwyg = "true";
defparam \Reg[15][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N16
cycloneive_lcell_comb \Mux10~18 (
// Equation(s):
// \Mux10~18_combout  = (ifid_ifinstr_o_22 & ((\Mux10~17_combout  & ((\Reg[15][21]~q ))) # (!\Mux10~17_combout  & (\Reg[14][21]~q )))) # (!ifid_ifinstr_o_22 & (\Mux10~17_combout ))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Mux10~17_combout ),
	.datac(\Reg[14][21]~q ),
	.datad(\Reg[15][21]~q ),
	.cin(gnd),
	.combout(\Mux10~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~18 .lut_mask = 16'hEC64;
defparam \Mux10~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N29
dffeas \Reg[6][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][21] .is_wysiwyg = "true";
defparam \Reg[6][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y39_N19
dffeas \Reg[7][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][21] .is_wysiwyg = "true";
defparam \Reg[7][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N18
cycloneive_lcell_comb \Mux10~13 (
// Equation(s):
// \Mux10~13_combout  = (\Mux10~12_combout  & (((\Reg[7][21]~q ) # (!ifid_ifinstr_o_22)))) # (!\Mux10~12_combout  & (\Reg[6][21]~q  & ((ifid_ifinstr_o_22))))

	.dataa(\Mux10~12_combout ),
	.datab(\Reg[6][21]~q ),
	.datac(\Reg[7][21]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux10~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~13 .lut_mask = 16'hE4AA;
defparam \Mux10~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N7
dffeas \Reg[2][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][21] .is_wysiwyg = "true";
defparam \Reg[2][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N19
dffeas \Reg[3][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][21] .is_wysiwyg = "true";
defparam \Reg[3][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N17
dffeas \Reg[1][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][21] .is_wysiwyg = "true";
defparam \Reg[1][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N16
cycloneive_lcell_comb \Mux10~14 (
// Equation(s):
// \Mux10~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[3][21]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[1][21]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[3][21]~q ),
	.datac(\Reg[1][21]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux10~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~14 .lut_mask = 16'h88A0;
defparam \Mux10~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N10
cycloneive_lcell_comb \Mux10~15 (
// Equation(s):
// \Mux10~15_combout  = (\Mux10~14_combout ) # ((ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & \Reg[2][21]~q )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[2][21]~q ),
	.datad(\Mux10~14_combout ),
	.cin(gnd),
	.combout(\Mux10~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~15 .lut_mask = 16'hFF20;
defparam \Mux10~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N8
cycloneive_lcell_comb \Mux10~16 (
// Equation(s):
// \Mux10~16_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & (\Mux10~13_combout )) # (!ifid_ifinstr_o_23 & ((\Mux10~15_combout )))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Mux10~13_combout ),
	.datad(\Mux10~15_combout ),
	.cin(gnd),
	.combout(\Mux10~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~16 .lut_mask = 16'hD9C8;
defparam \Mux10~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N31
dffeas \Reg[11][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][21] .is_wysiwyg = "true";
defparam \Reg[11][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N15
dffeas \Reg[8][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][21] .is_wysiwyg = "true";
defparam \Reg[8][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N17
dffeas \Reg[10][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][21] .is_wysiwyg = "true";
defparam \Reg[10][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N16
cycloneive_lcell_comb \Mux10~10 (
// Equation(s):
// \Mux10~10_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[10][21]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[8][21]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[8][21]~q ),
	.datac(\Reg[10][21]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux10~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~10 .lut_mask = 16'hFA44;
defparam \Mux10~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N17
dffeas \Reg[9][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][21] .is_wysiwyg = "true";
defparam \Reg[9][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N16
cycloneive_lcell_comb \Mux10~11 (
// Equation(s):
// \Mux10~11_combout  = (\Mux10~10_combout  & ((\Reg[11][21]~q ) # ((!ifid_ifinstr_o_21)))) # (!\Mux10~10_combout  & (((\Reg[9][21]~q  & ifid_ifinstr_o_21))))

	.dataa(\Reg[11][21]~q ),
	.datab(\Mux10~10_combout ),
	.datac(\Reg[9][21]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux10~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~11 .lut_mask = 16'hB8CC;
defparam \Mux10~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N3
dffeas \Reg[30][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][20] .is_wysiwyg = "true";
defparam \Reg[30][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N15
dffeas \Reg[18][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][20] .is_wysiwyg = "true";
defparam \Reg[18][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N16
cycloneive_lcell_comb \Reg[22][20]~feeder (
// Equation(s):
// \Reg[22][20]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat28),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[22][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[22][20]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[22][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N17
dffeas \Reg[22][20] (
	.clk(!CLK),
	.d(\Reg[22][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][20] .is_wysiwyg = "true";
defparam \Reg[22][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N14
cycloneive_lcell_comb \Mux11~2 (
// Equation(s):
// \Mux11~2_combout  = (ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24) # ((\Reg[22][20]~q )))) # (!ifid_ifinstr_o_23 & (!ifid_ifinstr_o_24 & (\Reg[18][20]~q )))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[18][20]~q ),
	.datad(\Reg[22][20]~q ),
	.cin(gnd),
	.combout(\Mux11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~2 .lut_mask = 16'hBA98;
defparam \Mux11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y30_N5
dffeas \Reg[26][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][20] .is_wysiwyg = "true";
defparam \Reg[26][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N22
cycloneive_lcell_comb \Mux11~3 (
// Equation(s):
// \Mux11~3_combout  = (ifid_ifinstr_o_24 & ((\Mux11~2_combout  & (\Reg[30][20]~q )) # (!\Mux11~2_combout  & ((\Reg[26][20]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux11~2_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[30][20]~q ),
	.datac(\Mux11~2_combout ),
	.datad(\Reg[26][20]~q ),
	.cin(gnd),
	.combout(\Mux11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~3 .lut_mask = 16'hDAD0;
defparam \Mux11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y32_N9
dffeas \Reg[16][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][20] .is_wysiwyg = "true";
defparam \Reg[16][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N8
cycloneive_lcell_comb \Mux11~4 (
// Equation(s):
// \Mux11~4_combout  = (ifid_ifinstr_o_23 & ((\Reg[20][20]~q ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((\Reg[16][20]~q  & !ifid_ifinstr_o_24))))

	.dataa(\Reg[20][20]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[16][20]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~4 .lut_mask = 16'hCCB8;
defparam \Mux11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N17
dffeas \Reg[28][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][20] .is_wysiwyg = "true";
defparam \Reg[28][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N16
cycloneive_lcell_comb \Mux11~5 (
// Equation(s):
// \Mux11~5_combout  = (\Mux11~4_combout  & (((\Reg[28][20]~q ) # (!ifid_ifinstr_o_24)))) # (!\Mux11~4_combout  & (\Reg[24][20]~q  & ((ifid_ifinstr_o_24))))

	.dataa(\Reg[24][20]~q ),
	.datab(\Mux11~4_combout ),
	.datac(\Reg[28][20]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux11~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~5 .lut_mask = 16'hE2CC;
defparam \Mux11~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N12
cycloneive_lcell_comb \Mux11~6 (
// Equation(s):
// \Mux11~6_combout  = (ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21) # ((\Mux11~3_combout )))) # (!ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & ((\Mux11~5_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux11~3_combout ),
	.datad(\Mux11~5_combout ),
	.cin(gnd),
	.combout(\Mux11~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~6 .lut_mask = 16'hB9A8;
defparam \Mux11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N9
dffeas \Reg[23][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][20] .is_wysiwyg = "true";
defparam \Reg[23][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N24
cycloneive_lcell_comb \Reg[31][20]~feeder (
// Equation(s):
// \Reg[31][20]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat28),
	.cin(gnd),
	.combout(\Reg[31][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[31][20]~feeder .lut_mask = 16'hFF00;
defparam \Reg[31][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N25
dffeas \Reg[31][20] (
	.clk(!CLK),
	.d(\Reg[31][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][20] .is_wysiwyg = "true";
defparam \Reg[31][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N3
dffeas \Reg[19][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][20] .is_wysiwyg = "true";
defparam \Reg[19][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N10
cycloneive_lcell_comb \Reg[27][20]~feeder (
// Equation(s):
// \Reg[27][20]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat28),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[27][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[27][20]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[27][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N11
dffeas \Reg[27][20] (
	.clk(!CLK),
	.d(\Reg[27][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][20] .is_wysiwyg = "true";
defparam \Reg[27][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N2
cycloneive_lcell_comb \Mux11~7 (
// Equation(s):
// \Mux11~7_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Reg[27][20]~q ))) # (!ifid_ifinstr_o_24 & (\Reg[19][20]~q ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[19][20]~q ),
	.datad(\Reg[27][20]~q ),
	.cin(gnd),
	.combout(\Mux11~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~7 .lut_mask = 16'hDC98;
defparam \Mux11~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N10
cycloneive_lcell_comb \Mux11~8 (
// Equation(s):
// \Mux11~8_combout  = (\Mux11~7_combout  & (((\Reg[31][20]~q ) # (!ifid_ifinstr_o_23)))) # (!\Mux11~7_combout  & (\Reg[23][20]~q  & ((ifid_ifinstr_o_23))))

	.dataa(\Reg[23][20]~q ),
	.datab(\Reg[31][20]~q ),
	.datac(\Mux11~7_combout ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux11~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~8 .lut_mask = 16'hCAF0;
defparam \Mux11~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N28
cycloneive_lcell_comb \Reg[21][20]~feeder (
// Equation(s):
// \Reg[21][20]~feeder_combout  = \wdat~59_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat28),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[21][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[21][20]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[21][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N29
dffeas \Reg[21][20] (
	.clk(!CLK),
	.d(\Reg[21][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][20] .is_wysiwyg = "true";
defparam \Reg[21][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N25
dffeas \Reg[29][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][20] .is_wysiwyg = "true";
defparam \Reg[29][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N23
dffeas \Reg[17][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][20] .is_wysiwyg = "true";
defparam \Reg[17][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N22
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// \Mux11~0_combout  = (ifid_ifinstr_o_23 & (((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[25][20]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[17][20]~q )))))

	.dataa(\Reg[25][20]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[17][20]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hEE30;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N24
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// \Mux11~1_combout  = (ifid_ifinstr_o_23 & ((\Mux11~0_combout  & ((\Reg[29][20]~q ))) # (!\Mux11~0_combout  & (\Reg[21][20]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux11~0_combout ))))

	.dataa(\Reg[21][20]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[29][20]~q ),
	.datad(\Mux11~0_combout ),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'hF388;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N21
dffeas \Reg[14][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][20] .is_wysiwyg = "true";
defparam \Reg[14][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N15
dffeas \Reg[12][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][20] .is_wysiwyg = "true";
defparam \Reg[12][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N13
dffeas \Reg[13][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][20] .is_wysiwyg = "true";
defparam \Reg[13][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N12
cycloneive_lcell_comb \Mux11~17 (
// Equation(s):
// \Mux11~17_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[13][20]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[12][20]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[12][20]~q ),
	.datac(\Reg[13][20]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux11~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~17 .lut_mask = 16'hFA44;
defparam \Mux11~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N15
dffeas \Reg[15][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][20] .is_wysiwyg = "true";
defparam \Reg[15][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N14
cycloneive_lcell_comb \Mux11~18 (
// Equation(s):
// \Mux11~18_combout  = (\Mux11~17_combout  & (((\Reg[15][20]~q ) # (!ifid_ifinstr_o_22)))) # (!\Mux11~17_combout  & (\Reg[14][20]~q  & ((ifid_ifinstr_o_22))))

	.dataa(\Reg[14][20]~q ),
	.datab(\Mux11~17_combout ),
	.datac(\Reg[15][20]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux11~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~18 .lut_mask = 16'hE2CC;
defparam \Mux11~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N29
dffeas \Reg[7][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][20] .is_wysiwyg = "true";
defparam \Reg[7][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y38_N19
dffeas \Reg[6][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][20] .is_wysiwyg = "true";
defparam \Reg[6][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y39_N1
dffeas \Reg[5][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][20] .is_wysiwyg = "true";
defparam \Reg[5][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N0
cycloneive_lcell_comb \Mux11~10 (
// Equation(s):
// \Mux11~10_combout  = (ifid_ifinstr_o_21 & (((\Reg[5][20]~q ) # (ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & (\Reg[4][20]~q  & ((!ifid_ifinstr_o_22))))

	.dataa(\Reg[4][20]~q ),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[5][20]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux11~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~10 .lut_mask = 16'hCCE2;
defparam \Mux11~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N18
cycloneive_lcell_comb \Mux11~11 (
// Equation(s):
// \Mux11~11_combout  = (ifid_ifinstr_o_22 & ((\Mux11~10_combout  & (\Reg[7][20]~q )) # (!\Mux11~10_combout  & ((\Reg[6][20]~q ))))) # (!ifid_ifinstr_o_22 & (((\Mux11~10_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[7][20]~q ),
	.datac(\Reg[6][20]~q ),
	.datad(\Mux11~10_combout ),
	.cin(gnd),
	.combout(\Mux11~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~11 .lut_mask = 16'hDDA0;
defparam \Mux11~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N15
dffeas \Reg[2][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][20] .is_wysiwyg = "true";
defparam \Reg[2][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N4
cycloneive_lcell_comb \Mux11~15 (
// Equation(s):
// \Mux11~15_combout  = (\Mux11~14_combout ) # ((!ifid_ifinstr_o_21 & (ifid_ifinstr_o_22 & \Reg[2][20]~q )))

	.dataa(\Mux11~14_combout ),
	.datab(ifid_ifinstr_o_21),
	.datac(ifid_ifinstr_o_22),
	.datad(\Reg[2][20]~q ),
	.cin(gnd),
	.combout(\Mux11~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~15 .lut_mask = 16'hBAAA;
defparam \Mux11~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N15
dffeas \Reg[9][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][20] .is_wysiwyg = "true";
defparam \Reg[9][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y35_N5
dffeas \Reg[11][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][20] .is_wysiwyg = "true";
defparam \Reg[11][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N21
dffeas \Reg[10][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][20] .is_wysiwyg = "true";
defparam \Reg[10][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N19
dffeas \Reg[8][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][20] .is_wysiwyg = "true";
defparam \Reg[8][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N18
cycloneive_lcell_comb \Mux11~12 (
// Equation(s):
// \Mux11~12_combout  = (ifid_ifinstr_o_22 & ((\Reg[10][20]~q ) # ((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & (((\Reg[8][20]~q  & !ifid_ifinstr_o_21))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[10][20]~q ),
	.datac(\Reg[8][20]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux11~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~12 .lut_mask = 16'hAAD8;
defparam \Mux11~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N4
cycloneive_lcell_comb \Mux11~13 (
// Equation(s):
// \Mux11~13_combout  = (ifid_ifinstr_o_21 & ((\Mux11~12_combout  & ((\Reg[11][20]~q ))) # (!\Mux11~12_combout  & (\Reg[9][20]~q )))) # (!ifid_ifinstr_o_21 & (((\Mux11~12_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[9][20]~q ),
	.datac(\Reg[11][20]~q ),
	.datad(\Mux11~12_combout ),
	.cin(gnd),
	.combout(\Mux11~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~13 .lut_mask = 16'hF588;
defparam \Mux11~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N18
cycloneive_lcell_comb \Mux11~16 (
// Equation(s):
// \Mux11~16_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Mux11~13_combout )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & (\Mux11~15_combout )))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Mux11~15_combout ),
	.datad(\Mux11~13_combout ),
	.cin(gnd),
	.combout(\Mux11~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~16 .lut_mask = 16'hBA98;
defparam \Mux11~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y30_N19
dffeas \Reg[18][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][18] .is_wysiwyg = "true";
defparam \Reg[18][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N8
cycloneive_lcell_comb \Reg[22][18]~feeder (
// Equation(s):
// \Reg[22][18]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat29),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[22][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[22][18]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[22][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N9
dffeas \Reg[22][18] (
	.clk(!CLK),
	.d(\Reg[22][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][18] .is_wysiwyg = "true";
defparam \Reg[22][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N18
cycloneive_lcell_comb \Mux13~2 (
// Equation(s):
// \Mux13~2_combout  = (ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24) # ((\Reg[22][18]~q )))) # (!ifid_ifinstr_o_23 & (!ifid_ifinstr_o_24 & (\Reg[18][18]~q )))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[18][18]~q ),
	.datad(\Reg[22][18]~q ),
	.cin(gnd),
	.combout(\Mux13~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~2 .lut_mask = 16'hBA98;
defparam \Mux13~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N7
dffeas \Reg[30][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][18] .is_wysiwyg = "true";
defparam \Reg[30][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N17
dffeas \Reg[26][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][18] .is_wysiwyg = "true";
defparam \Reg[26][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N14
cycloneive_lcell_comb \Mux13~3 (
// Equation(s):
// \Mux13~3_combout  = (ifid_ifinstr_o_24 & ((\Mux13~2_combout  & (\Reg[30][18]~q )) # (!\Mux13~2_combout  & ((\Reg[26][18]~q ))))) # (!ifid_ifinstr_o_24 & (\Mux13~2_combout ))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux13~2_combout ),
	.datac(\Reg[30][18]~q ),
	.datad(\Reg[26][18]~q ),
	.cin(gnd),
	.combout(\Mux13~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~3 .lut_mask = 16'hE6C4;
defparam \Mux13~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y32_N27
dffeas \Reg[24][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][18] .is_wysiwyg = "true";
defparam \Reg[24][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N21
dffeas \Reg[28][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][18] .is_wysiwyg = "true";
defparam \Reg[28][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N20
cycloneive_lcell_comb \Mux13~5 (
// Equation(s):
// \Mux13~5_combout  = (\Mux13~4_combout  & (((\Reg[28][18]~q ) # (!ifid_ifinstr_o_24)))) # (!\Mux13~4_combout  & (\Reg[24][18]~q  & ((ifid_ifinstr_o_24))))

	.dataa(\Mux13~4_combout ),
	.datab(\Reg[24][18]~q ),
	.datac(\Reg[28][18]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux13~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~5 .lut_mask = 16'hE4AA;
defparam \Mux13~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N6
cycloneive_lcell_comb \Mux13~6 (
// Equation(s):
// \Mux13~6_combout  = (ifid_ifinstr_o_22 & ((\Mux13~3_combout ) # ((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & (((\Mux13~5_combout  & !ifid_ifinstr_o_21))))

	.dataa(\Mux13~3_combout ),
	.datab(\Mux13~5_combout ),
	.datac(ifid_ifinstr_o_22),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux13~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~6 .lut_mask = 16'hF0AC;
defparam \Mux13~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N20
cycloneive_lcell_comb \Reg[31][18]~feeder (
// Equation(s):
// \Reg[31][18]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat29),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[31][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[31][18]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[31][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y29_N21
dffeas \Reg[31][18] (
	.clk(!CLK),
	.d(\Reg[31][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][18] .is_wysiwyg = "true";
defparam \Reg[31][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N29
dffeas \Reg[23][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][18] .is_wysiwyg = "true";
defparam \Reg[23][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N7
dffeas \Reg[19][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][18] .is_wysiwyg = "true";
defparam \Reg[19][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N6
cycloneive_lcell_comb \Reg[27][18]~feeder (
// Equation(s):
// \Reg[27][18]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat29),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[27][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[27][18]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[27][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N7
dffeas \Reg[27][18] (
	.clk(!CLK),
	.d(\Reg[27][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][18] .is_wysiwyg = "true";
defparam \Reg[27][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N6
cycloneive_lcell_comb \Mux13~7 (
// Equation(s):
// \Mux13~7_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & ((\Reg[27][18]~q ))) # (!ifid_ifinstr_o_24 & (\Reg[19][18]~q ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[19][18]~q ),
	.datad(\Reg[27][18]~q ),
	.cin(gnd),
	.combout(\Mux13~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~7 .lut_mask = 16'hDC98;
defparam \Mux13~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N8
cycloneive_lcell_comb \Mux13~8 (
// Equation(s):
// \Mux13~8_combout  = (ifid_ifinstr_o_23 & ((\Mux13~7_combout  & (\Reg[31][18]~q )) # (!\Mux13~7_combout  & ((\Reg[23][18]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux13~7_combout ))))

	.dataa(\Reg[31][18]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[23][18]~q ),
	.datad(\Mux13~7_combout ),
	.cin(gnd),
	.combout(\Mux13~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~8 .lut_mask = 16'hBBC0;
defparam \Mux13~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N14
cycloneive_lcell_comb \Reg[21][18]~feeder (
// Equation(s):
// \Reg[21][18]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat29),
	.cin(gnd),
	.combout(\Reg[21][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[21][18]~feeder .lut_mask = 16'hFF00;
defparam \Reg[21][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y38_N15
dffeas \Reg[21][18] (
	.clk(!CLK),
	.d(\Reg[21][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][18] .is_wysiwyg = "true";
defparam \Reg[21][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N9
dffeas \Reg[29][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][18] .is_wysiwyg = "true";
defparam \Reg[29][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N16
cycloneive_lcell_comb \Reg[25][18]~feeder (
// Equation(s):
// \Reg[25][18]~feeder_combout  = \wdat~61_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat29),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[25][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][18]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[25][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y32_N17
dffeas \Reg[25][18] (
	.clk(!CLK),
	.d(\Reg[25][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][18] .is_wysiwyg = "true";
defparam \Reg[25][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N29
dffeas \Reg[17][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][18] .is_wysiwyg = "true";
defparam \Reg[17][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N6
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// \Mux13~0_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[25][18]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[17][18]~q )))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[25][18]~q ),
	.datad(\Reg[17][18]~q ),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hD9C8;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N8
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// \Mux13~1_combout  = (ifid_ifinstr_o_23 & ((\Mux13~0_combout  & ((\Reg[29][18]~q ))) # (!\Mux13~0_combout  & (\Reg[21][18]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux13~0_combout ))))

	.dataa(\Reg[21][18]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[29][18]~q ),
	.datad(\Mux13~0_combout ),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'hF388;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N13
dffeas \Reg[14][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][18] .is_wysiwyg = "true";
defparam \Reg[14][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N3
dffeas \Reg[15][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][18] .is_wysiwyg = "true";
defparam \Reg[15][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N25
dffeas \Reg[13][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][18] .is_wysiwyg = "true";
defparam \Reg[13][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N27
dffeas \Reg[12][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][18] .is_wysiwyg = "true";
defparam \Reg[12][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N26
cycloneive_lcell_comb \Mux13~17 (
// Equation(s):
// \Mux13~17_combout  = (ifid_ifinstr_o_22 & (((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & (\Reg[13][18]~q )) # (!ifid_ifinstr_o_21 & ((\Reg[12][18]~q )))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[13][18]~q ),
	.datac(\Reg[12][18]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux13~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~17 .lut_mask = 16'hEE50;
defparam \Mux13~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N2
cycloneive_lcell_comb \Mux13~18 (
// Equation(s):
// \Mux13~18_combout  = (ifid_ifinstr_o_22 & ((\Mux13~17_combout  & ((\Reg[15][18]~q ))) # (!\Mux13~17_combout  & (\Reg[14][18]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux13~17_combout ))))

	.dataa(\Reg[14][18]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[15][18]~q ),
	.datad(\Mux13~17_combout ),
	.cin(gnd),
	.combout(\Mux13~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~18 .lut_mask = 16'hF388;
defparam \Mux13~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N5
dffeas \Reg[5][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][18] .is_wysiwyg = "true";
defparam \Reg[5][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N3
dffeas \Reg[4][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][18] .is_wysiwyg = "true";
defparam \Reg[4][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N4
cycloneive_lcell_comb \Mux13~10 (
// Equation(s):
// \Mux13~10_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22) # ((\Reg[5][18]~q )))) # (!ifid_ifinstr_o_21 & (!ifid_ifinstr_o_22 & ((\Reg[4][18]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[5][18]~q ),
	.datad(\Reg[4][18]~q ),
	.cin(gnd),
	.combout(\Mux13~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~10 .lut_mask = 16'hB9A8;
defparam \Mux13~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N1
dffeas \Reg[6][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][18] .is_wysiwyg = "true";
defparam \Reg[6][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y39_N19
dffeas \Reg[7][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][18] .is_wysiwyg = "true";
defparam \Reg[7][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N0
cycloneive_lcell_comb \Mux13~11 (
// Equation(s):
// \Mux13~11_combout  = (\Mux13~10_combout  & (((\Reg[7][18]~q )) # (!ifid_ifinstr_o_22))) # (!\Mux13~10_combout  & (ifid_ifinstr_o_22 & (\Reg[6][18]~q )))

	.dataa(\Mux13~10_combout ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[6][18]~q ),
	.datad(\Reg[7][18]~q ),
	.cin(gnd),
	.combout(\Mux13~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~11 .lut_mask = 16'hEA62;
defparam \Mux13~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y32_N11
dffeas \Reg[9][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][18] .is_wysiwyg = "true";
defparam \Reg[9][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y36_N17
dffeas \Reg[11][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][18] .is_wysiwyg = "true";
defparam \Reg[11][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N9
dffeas \Reg[10][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][18] .is_wysiwyg = "true";
defparam \Reg[10][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N7
dffeas \Reg[8][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][18] .is_wysiwyg = "true";
defparam \Reg[8][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N6
cycloneive_lcell_comb \Mux13~12 (
// Equation(s):
// \Mux13~12_combout  = (ifid_ifinstr_o_22 & ((\Reg[10][18]~q ) # ((ifid_ifinstr_o_21)))) # (!ifid_ifinstr_o_22 & (((\Reg[8][18]~q  & !ifid_ifinstr_o_21))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[10][18]~q ),
	.datac(\Reg[8][18]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux13~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~12 .lut_mask = 16'hAAD8;
defparam \Mux13~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N16
cycloneive_lcell_comb \Mux13~13 (
// Equation(s):
// \Mux13~13_combout  = (ifid_ifinstr_o_21 & ((\Mux13~12_combout  & ((\Reg[11][18]~q ))) # (!\Mux13~12_combout  & (\Reg[9][18]~q )))) # (!ifid_ifinstr_o_21 & (((\Mux13~12_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[9][18]~q ),
	.datac(\Reg[11][18]~q ),
	.datad(\Mux13~12_combout ),
	.cin(gnd),
	.combout(\Mux13~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~13 .lut_mask = 16'hF588;
defparam \Mux13~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N31
dffeas \Reg[1][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][18] .is_wysiwyg = "true";
defparam \Reg[1][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N13
dffeas \Reg[3][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][18] .is_wysiwyg = "true";
defparam \Reg[3][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N30
cycloneive_lcell_comb \Mux13~14 (
// Equation(s):
// \Mux13~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][18]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][18]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[1][18]~q ),
	.datad(\Reg[3][18]~q ),
	.cin(gnd),
	.combout(\Mux13~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~14 .lut_mask = 16'hA820;
defparam \Mux13~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y36_N11
dffeas \Reg[2][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][18] .is_wysiwyg = "true";
defparam \Reg[2][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N10
cycloneive_lcell_comb \Mux13~15 (
// Equation(s):
// \Mux13~15_combout  = (\Mux13~14_combout ) # ((!ifid_ifinstr_o_21 & (\Reg[2][18]~q  & ifid_ifinstr_o_22)))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux13~14_combout ),
	.datac(\Reg[2][18]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux13~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~15 .lut_mask = 16'hDCCC;
defparam \Mux13~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N20
cycloneive_lcell_comb \Mux13~16 (
// Equation(s):
// \Mux13~16_combout  = (ifid_ifinstr_o_24 & ((\Mux13~13_combout ) # ((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & (((!ifid_ifinstr_o_23 & \Mux13~15_combout ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux13~13_combout ),
	.datac(ifid_ifinstr_o_23),
	.datad(\Mux13~15_combout ),
	.cin(gnd),
	.combout(\Mux13~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~16 .lut_mask = 16'hADA8;
defparam \Mux13~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y29_N7
dffeas \Reg[27][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][19] .is_wysiwyg = "true";
defparam \Reg[27][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y29_N13
dffeas \Reg[31][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][19] .is_wysiwyg = "true";
defparam \Reg[31][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N18
cycloneive_lcell_comb \Reg[23][19]~feeder (
// Equation(s):
// \Reg[23][19]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat30),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[23][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[23][19]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[23][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N19
dffeas \Reg[23][19] (
	.clk(!CLK),
	.d(\Reg[23][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][19] .is_wysiwyg = "true";
defparam \Reg[23][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N13
dffeas \Reg[19][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][19] .is_wysiwyg = "true";
defparam \Reg[19][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N12
cycloneive_lcell_comb \Mux12~7 (
// Equation(s):
// \Mux12~7_combout  = (ifid_ifinstr_o_23 & ((\Reg[23][19]~q ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((\Reg[19][19]~q  & !ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[23][19]~q ),
	.datac(\Reg[19][19]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux12~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~7 .lut_mask = 16'hAAD8;
defparam \Mux12~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N10
cycloneive_lcell_comb \Mux12~8 (
// Equation(s):
// \Mux12~8_combout  = (\Mux12~7_combout  & (((\Reg[31][19]~q ) # (!ifid_ifinstr_o_24)))) # (!\Mux12~7_combout  & (\Reg[27][19]~q  & ((ifid_ifinstr_o_24))))

	.dataa(\Reg[27][19]~q ),
	.datab(\Reg[31][19]~q ),
	.datac(\Mux12~7_combout ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux12~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~8 .lut_mask = 16'hCAF0;
defparam \Mux12~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N19
dffeas \Reg[17][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][19] .is_wysiwyg = "true";
defparam \Reg[17][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N11
dffeas \Reg[21][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][19] .is_wysiwyg = "true";
defparam \Reg[21][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N18
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (ifid_ifinstr_o_24 & (ifid_ifinstr_o_23)) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[21][19]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[17][19]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[17][19]~q ),
	.datad(\Reg[21][19]~q ),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hDC98;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y38_N1
dffeas \Reg[29][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][19] .is_wysiwyg = "true";
defparam \Reg[29][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N25
dffeas \Reg[25][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][19] .is_wysiwyg = "true";
defparam \Reg[25][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N0
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// \Mux12~1_combout  = (ifid_ifinstr_o_24 & ((\Mux12~0_combout  & (\Reg[29][19]~q )) # (!\Mux12~0_combout  & ((\Reg[25][19]~q ))))) # (!ifid_ifinstr_o_24 & (\Mux12~0_combout ))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Mux12~0_combout ),
	.datac(\Reg[29][19]~q ),
	.datad(\Reg[25][19]~q ),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hE6C4;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N25
dffeas \Reg[22][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][19] .is_wysiwyg = "true";
defparam \Reg[22][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N13
dffeas \Reg[26][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][19] .is_wysiwyg = "true";
defparam \Reg[26][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N12
cycloneive_lcell_comb \Mux12~2 (
// Equation(s):
// \Mux12~2_combout  = (ifid_ifinstr_o_24 & (((\Reg[26][19]~q ) # (ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & (\Reg[18][19]~q  & ((!ifid_ifinstr_o_23))))

	.dataa(\Reg[18][19]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[26][19]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux12~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~2 .lut_mask = 16'hCCE2;
defparam \Mux12~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N24
cycloneive_lcell_comb \Mux12~3 (
// Equation(s):
// \Mux12~3_combout  = (ifid_ifinstr_o_23 & ((\Mux12~2_combout  & (\Reg[30][19]~q )) # (!\Mux12~2_combout  & ((\Reg[22][19]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux12~2_combout ))))

	.dataa(\Reg[30][19]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[22][19]~q ),
	.datad(\Mux12~2_combout ),
	.cin(gnd),
	.combout(\Mux12~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~3 .lut_mask = 16'hBBC0;
defparam \Mux12~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y33_N7
dffeas \Reg[20][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][19] .is_wysiwyg = "true";
defparam \Reg[20][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y33_N1
dffeas \Reg[16][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][19] .is_wysiwyg = "true";
defparam \Reg[16][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N0
cycloneive_lcell_comb \Mux12~4 (
// Equation(s):
// \Mux12~4_combout  = (ifid_ifinstr_o_24 & ((\Reg[24][19]~q ) # ((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & (((\Reg[16][19]~q  & !ifid_ifinstr_o_23))))

	.dataa(\Reg[24][19]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[16][19]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux12~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~4 .lut_mask = 16'hCCB8;
defparam \Mux12~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y34_N12
cycloneive_lcell_comb \Mux12~5 (
// Equation(s):
// \Mux12~5_combout  = (ifid_ifinstr_o_23 & ((\Mux12~4_combout  & (\Reg[28][19]~q )) # (!\Mux12~4_combout  & ((\Reg[20][19]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux12~4_combout ))))

	.dataa(\Reg[28][19]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[20][19]~q ),
	.datad(\Mux12~4_combout ),
	.cin(gnd),
	.combout(\Mux12~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~5 .lut_mask = 16'hBBC0;
defparam \Mux12~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N20
cycloneive_lcell_comb \Mux12~6 (
// Equation(s):
// \Mux12~6_combout  = (ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21) # ((\Mux12~3_combout )))) # (!ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & ((\Mux12~5_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux12~3_combout ),
	.datad(\Mux12~5_combout ),
	.cin(gnd),
	.combout(\Mux12~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~6 .lut_mask = 16'hB9A8;
defparam \Mux12~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N27
dffeas \Reg[11][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][19] .is_wysiwyg = "true";
defparam \Reg[11][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N3
dffeas \Reg[8][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][19] .is_wysiwyg = "true";
defparam \Reg[8][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N13
dffeas \Reg[10][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][19] .is_wysiwyg = "true";
defparam \Reg[10][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N12
cycloneive_lcell_comb \Mux12~10 (
// Equation(s):
// \Mux12~10_combout  = (ifid_ifinstr_o_21 & (((ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[10][19]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[8][19]~q ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[8][19]~q ),
	.datac(\Reg[10][19]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux12~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~10 .lut_mask = 16'hFA44;
defparam \Mux12~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N1
dffeas \Reg[9][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][19] .is_wysiwyg = "true";
defparam \Reg[9][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N0
cycloneive_lcell_comb \Mux12~11 (
// Equation(s):
// \Mux12~11_combout  = (\Mux12~10_combout  & ((\Reg[11][19]~q ) # ((!ifid_ifinstr_o_21)))) # (!\Mux12~10_combout  & (((\Reg[9][19]~q  & ifid_ifinstr_o_21))))

	.dataa(\Reg[11][19]~q ),
	.datab(\Mux12~10_combout ),
	.datac(\Reg[9][19]~q ),
	.datad(ifid_ifinstr_o_21),
	.cin(gnd),
	.combout(\Mux12~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~11 .lut_mask = 16'hB8CC;
defparam \Mux12~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y34_N23
dffeas \Reg[12][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][19] .is_wysiwyg = "true";
defparam \Reg[12][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y34_N29
dffeas \Reg[13][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][19] .is_wysiwyg = "true";
defparam \Reg[13][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N22
cycloneive_lcell_comb \Mux12~17 (
// Equation(s):
// \Mux12~17_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[13][19]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[12][19]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[12][19]~q ),
	.datad(\Reg[13][19]~q ),
	.cin(gnd),
	.combout(\Mux12~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~17 .lut_mask = 16'hDC98;
defparam \Mux12~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N18
cycloneive_lcell_comb \Reg[15][19]~feeder (
// Equation(s):
// \Reg[15][19]~feeder_combout  = \wdat~63_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat30),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[15][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[15][19]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[15][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N19
dffeas \Reg[15][19] (
	.clk(!CLK),
	.d(\Reg[15][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][19] .is_wysiwyg = "true";
defparam \Reg[15][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N5
dffeas \Reg[14][19] (
	.clk(!CLK),
	.d(wdat30),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][19] .is_wysiwyg = "true";
defparam \Reg[14][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N8
cycloneive_lcell_comb \Mux12~18 (
// Equation(s):
// \Mux12~18_combout  = (\Mux12~17_combout  & ((\Reg[15][19]~q ) # ((!ifid_ifinstr_o_22)))) # (!\Mux12~17_combout  & (((\Reg[14][19]~q  & ifid_ifinstr_o_22))))

	.dataa(\Mux12~17_combout ),
	.datab(\Reg[15][19]~q ),
	.datac(\Reg[14][19]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux12~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~18 .lut_mask = 16'hD8AA;
defparam \Mux12~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N5
dffeas \Reg[6][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][19] .is_wysiwyg = "true";
defparam \Reg[6][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y39_N15
dffeas \Reg[7][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][19] .is_wysiwyg = "true";
defparam \Reg[7][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y39_N19
dffeas \Reg[4][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][19] .is_wysiwyg = "true";
defparam \Reg[4][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y39_N17
dffeas \Reg[5][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][19] .is_wysiwyg = "true";
defparam \Reg[5][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N18
cycloneive_lcell_comb \Mux12~12 (
// Equation(s):
// \Mux12~12_combout  = (ifid_ifinstr_o_22 & (ifid_ifinstr_o_21)) # (!ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21 & ((\Reg[5][19]~q ))) # (!ifid_ifinstr_o_21 & (\Reg[4][19]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[4][19]~q ),
	.datad(\Reg[5][19]~q ),
	.cin(gnd),
	.combout(\Mux12~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~12 .lut_mask = 16'hDC98;
defparam \Mux12~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N14
cycloneive_lcell_comb \Mux12~13 (
// Equation(s):
// \Mux12~13_combout  = (ifid_ifinstr_o_22 & ((\Mux12~12_combout  & ((\Reg[7][19]~q ))) # (!\Mux12~12_combout  & (\Reg[6][19]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux12~12_combout ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(\Reg[6][19]~q ),
	.datac(\Reg[7][19]~q ),
	.datad(\Mux12~12_combout ),
	.cin(gnd),
	.combout(\Mux12~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~13 .lut_mask = 16'hF588;
defparam \Mux12~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y35_N5
dffeas \Reg[1][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][19] .is_wysiwyg = "true";
defparam \Reg[1][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N3
dffeas \Reg[3][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][19] .is_wysiwyg = "true";
defparam \Reg[3][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N4
cycloneive_lcell_comb \Mux12~14 (
// Equation(s):
// \Mux12~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][19]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][19]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[1][19]~q ),
	.datad(\Reg[3][19]~q ),
	.cin(gnd),
	.combout(\Mux12~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~14 .lut_mask = 16'hC840;
defparam \Mux12~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y36_N31
dffeas \Reg[2][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][19] .is_wysiwyg = "true";
defparam \Reg[2][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y36_N30
cycloneive_lcell_comb \Mux12~15 (
// Equation(s):
// \Mux12~15_combout  = (\Mux12~14_combout ) # ((!ifid_ifinstr_o_21 & (\Reg[2][19]~q  & ifid_ifinstr_o_22)))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Mux12~14_combout ),
	.datac(\Reg[2][19]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux12~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~15 .lut_mask = 16'hDCCC;
defparam \Mux12~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N24
cycloneive_lcell_comb \Mux12~16 (
// Equation(s):
// \Mux12~16_combout  = (ifid_ifinstr_o_23 & ((\Mux12~13_combout ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((!ifid_ifinstr_o_24 & \Mux12~15_combout ))))

	.dataa(\Mux12~13_combout ),
	.datab(ifid_ifinstr_o_23),
	.datac(ifid_ifinstr_o_24),
	.datad(\Mux12~15_combout ),
	.cin(gnd),
	.combout(\Mux12~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~16 .lut_mask = 16'hCBC8;
defparam \Mux12~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N7
dffeas \Reg[31][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[31][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[31][17] .is_wysiwyg = "true";
defparam \Reg[31][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N2
cycloneive_lcell_comb \Reg[23][17]~feeder (
// Equation(s):
// \Reg[23][17]~feeder_combout  = \wdat~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat31),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[23][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[23][17]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[23][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N3
dffeas \Reg[23][17] (
	.clk(!CLK),
	.d(\Reg[23][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[23][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[23][17] .is_wysiwyg = "true";
defparam \Reg[23][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N17
dffeas \Reg[19][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][17] .is_wysiwyg = "true";
defparam \Reg[19][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N16
cycloneive_lcell_comb \Mux14~7 (
// Equation(s):
// \Mux14~7_combout  = (ifid_ifinstr_o_23 & ((\Reg[23][17]~q ) # ((ifid_ifinstr_o_24)))) # (!ifid_ifinstr_o_23 & (((\Reg[19][17]~q  & !ifid_ifinstr_o_24))))

	.dataa(ifid_ifinstr_o_23),
	.datab(\Reg[23][17]~q ),
	.datac(\Reg[19][17]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux14~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~7 .lut_mask = 16'hAAD8;
defparam \Mux14~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N17
dffeas \Reg[27][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][17] .is_wysiwyg = "true";
defparam \Reg[27][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N26
cycloneive_lcell_comb \Mux14~8 (
// Equation(s):
// \Mux14~8_combout  = (\Mux14~7_combout  & ((\Reg[31][17]~q ) # ((!ifid_ifinstr_o_24)))) # (!\Mux14~7_combout  & (((\Reg[27][17]~q  & ifid_ifinstr_o_24))))

	.dataa(\Reg[31][17]~q ),
	.datab(\Mux14~7_combout ),
	.datac(\Reg[27][17]~q ),
	.datad(ifid_ifinstr_o_24),
	.cin(gnd),
	.combout(\Mux14~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~8 .lut_mask = 16'hB8CC;
defparam \Mux14~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N5
dffeas \Reg[28][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][17] .is_wysiwyg = "true";
defparam \Reg[28][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y32_N3
dffeas \Reg[24][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][17] .is_wysiwyg = "true";
defparam \Reg[24][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y32_N21
dffeas \Reg[16][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][17] .is_wysiwyg = "true";
defparam \Reg[16][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N2
cycloneive_lcell_comb \Mux14~4 (
// Equation(s):
// \Mux14~4_combout  = (ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23) # ((\Reg[24][17]~q )))) # (!ifid_ifinstr_o_24 & (!ifid_ifinstr_o_23 & ((\Reg[16][17]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[24][17]~q ),
	.datad(\Reg[16][17]~q ),
	.cin(gnd),
	.combout(\Mux14~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~4 .lut_mask = 16'hB9A8;
defparam \Mux14~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N4
cycloneive_lcell_comb \Mux14~5 (
// Equation(s):
// \Mux14~5_combout  = (ifid_ifinstr_o_23 & ((\Mux14~4_combout  & ((\Reg[28][17]~q ))) # (!\Mux14~4_combout  & (\Reg[20][17]~q )))) # (!ifid_ifinstr_o_23 & (((\Mux14~4_combout ))))

	.dataa(\Reg[20][17]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[28][17]~q ),
	.datad(\Mux14~4_combout ),
	.cin(gnd),
	.combout(\Mux14~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~5 .lut_mask = 16'hF388;
defparam \Mux14~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N9
dffeas \Reg[22][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][17] .is_wysiwyg = "true";
defparam \Reg[22][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N1
dffeas \Reg[26][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[26][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[26][17] .is_wysiwyg = "true";
defparam \Reg[26][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N11
dffeas \Reg[18][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][17] .is_wysiwyg = "true";
defparam \Reg[18][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N0
cycloneive_lcell_comb \Mux14~2 (
// Equation(s):
// \Mux14~2_combout  = (ifid_ifinstr_o_23 & (ifid_ifinstr_o_24)) # (!ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24 & (\Reg[26][17]~q )) # (!ifid_ifinstr_o_24 & ((\Reg[18][17]~q )))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[26][17]~q ),
	.datad(\Reg[18][17]~q ),
	.cin(gnd),
	.combout(\Mux14~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~2 .lut_mask = 16'hD9C8;
defparam \Mux14~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N8
cycloneive_lcell_comb \Mux14~3 (
// Equation(s):
// \Mux14~3_combout  = (ifid_ifinstr_o_23 & ((\Mux14~2_combout  & (\Reg[30][17]~q )) # (!\Mux14~2_combout  & ((\Reg[22][17]~q ))))) # (!ifid_ifinstr_o_23 & (((\Mux14~2_combout ))))

	.dataa(\Reg[30][17]~q ),
	.datab(ifid_ifinstr_o_23),
	.datac(\Reg[22][17]~q ),
	.datad(\Mux14~2_combout ),
	.cin(gnd),
	.combout(\Mux14~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~3 .lut_mask = 16'hBBC0;
defparam \Mux14~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N2
cycloneive_lcell_comb \Mux14~6 (
// Equation(s):
// \Mux14~6_combout  = (ifid_ifinstr_o_22 & ((ifid_ifinstr_o_21) # ((\Mux14~3_combout )))) # (!ifid_ifinstr_o_22 & (!ifid_ifinstr_o_21 & (\Mux14~5_combout )))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Mux14~5_combout ),
	.datad(\Mux14~3_combout ),
	.cin(gnd),
	.combout(\Mux14~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~6 .lut_mask = 16'hBA98;
defparam \Mux14~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y38_N5
dffeas \Reg[29][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[29][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[29][17] .is_wysiwyg = "true";
defparam \Reg[29][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y37_N11
dffeas \Reg[25][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][17] .is_wysiwyg = "true";
defparam \Reg[25][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y38_N29
dffeas \Reg[17][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][17] .is_wysiwyg = "true";
defparam \Reg[17][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y38_N31
dffeas \Reg[21][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][17] .is_wysiwyg = "true";
defparam \Reg[21][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N30
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// \Mux14~0_combout  = (ifid_ifinstr_o_24 & (((ifid_ifinstr_o_23)))) # (!ifid_ifinstr_o_24 & ((ifid_ifinstr_o_23 & ((\Reg[21][17]~q ))) # (!ifid_ifinstr_o_23 & (\Reg[17][17]~q ))))

	.dataa(ifid_ifinstr_o_24),
	.datab(\Reg[17][17]~q ),
	.datac(\Reg[21][17]~q ),
	.datad(ifid_ifinstr_o_23),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hFA44;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N10
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// \Mux14~1_combout  = (ifid_ifinstr_o_24 & ((\Mux14~0_combout  & (\Reg[29][17]~q )) # (!\Mux14~0_combout  & ((\Reg[25][17]~q ))))) # (!ifid_ifinstr_o_24 & (((\Mux14~0_combout ))))

	.dataa(\Reg[29][17]~q ),
	.datab(ifid_ifinstr_o_24),
	.datac(\Reg[25][17]~q ),
	.datad(\Mux14~0_combout ),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hBBC0;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N9
dffeas \Reg[6][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][17] .is_wysiwyg = "true";
defparam \Reg[6][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y39_N11
dffeas \Reg[7][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[7][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[7][17] .is_wysiwyg = "true";
defparam \Reg[7][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N10
cycloneive_lcell_comb \Mux14~13 (
// Equation(s):
// \Mux14~13_combout  = (\Mux14~12_combout  & (((\Reg[7][17]~q ) # (!ifid_ifinstr_o_22)))) # (!\Mux14~12_combout  & (\Reg[6][17]~q  & ((ifid_ifinstr_o_22))))

	.dataa(\Mux14~12_combout ),
	.datab(\Reg[6][17]~q ),
	.datac(\Reg[7][17]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux14~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~13 .lut_mask = 16'hE4AA;
defparam \Mux14~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y35_N25
dffeas \Reg[1][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][17] .is_wysiwyg = "true";
defparam \Reg[1][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y35_N11
dffeas \Reg[3][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[3][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[3][17] .is_wysiwyg = "true";
defparam \Reg[3][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N24
cycloneive_lcell_comb \Mux14~14 (
// Equation(s):
// \Mux14~14_combout  = (ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & ((\Reg[3][17]~q ))) # (!ifid_ifinstr_o_22 & (\Reg[1][17]~q ))))

	.dataa(ifid_ifinstr_o_22),
	.datab(ifid_ifinstr_o_21),
	.datac(\Reg[1][17]~q ),
	.datad(\Reg[3][17]~q ),
	.cin(gnd),
	.combout(\Mux14~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~14 .lut_mask = 16'hC840;
defparam \Mux14~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N21
dffeas \Reg[2][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][17] .is_wysiwyg = "true";
defparam \Reg[2][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N2
cycloneive_lcell_comb \Mux14~15 (
// Equation(s):
// \Mux14~15_combout  = (\Mux14~14_combout ) # ((!ifid_ifinstr_o_21 & (ifid_ifinstr_o_22 & \Reg[2][17]~q )))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Mux14~14_combout ),
	.datad(\Reg[2][17]~q ),
	.cin(gnd),
	.combout(\Mux14~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~15 .lut_mask = 16'hF4F0;
defparam \Mux14~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N24
cycloneive_lcell_comb \Mux14~16 (
// Equation(s):
// \Mux14~16_combout  = (ifid_ifinstr_o_23 & ((ifid_ifinstr_o_24) # ((\Mux14~13_combout )))) # (!ifid_ifinstr_o_23 & (!ifid_ifinstr_o_24 & ((\Mux14~15_combout ))))

	.dataa(ifid_ifinstr_o_23),
	.datab(ifid_ifinstr_o_24),
	.datac(\Mux14~13_combout ),
	.datad(\Mux14~15_combout ),
	.cin(gnd),
	.combout(\Mux14~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~16 .lut_mask = 16'hB9A8;
defparam \Mux14~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N29
dffeas \Reg[11][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[11][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[11][17] .is_wysiwyg = "true";
defparam \Reg[11][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y35_N11
dffeas \Reg[9][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][17] .is_wysiwyg = "true";
defparam \Reg[9][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N25
dffeas \Reg[10][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][17] .is_wysiwyg = "true";
defparam \Reg[10][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N3
dffeas \Reg[8][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][17] .is_wysiwyg = "true";
defparam \Reg[8][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N24
cycloneive_lcell_comb \Mux14~10 (
// Equation(s):
// \Mux14~10_combout  = (ifid_ifinstr_o_21 & (ifid_ifinstr_o_22)) # (!ifid_ifinstr_o_21 & ((ifid_ifinstr_o_22 & (\Reg[10][17]~q )) # (!ifid_ifinstr_o_22 & ((\Reg[8][17]~q )))))

	.dataa(ifid_ifinstr_o_21),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[10][17]~q ),
	.datad(\Reg[8][17]~q ),
	.cin(gnd),
	.combout(\Mux14~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~10 .lut_mask = 16'hD9C8;
defparam \Mux14~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N10
cycloneive_lcell_comb \Mux14~11 (
// Equation(s):
// \Mux14~11_combout  = (ifid_ifinstr_o_21 & ((\Mux14~10_combout  & (\Reg[11][17]~q )) # (!\Mux14~10_combout  & ((\Reg[9][17]~q ))))) # (!ifid_ifinstr_o_21 & (((\Mux14~10_combout ))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[11][17]~q ),
	.datac(\Reg[9][17]~q ),
	.datad(\Mux14~10_combout ),
	.cin(gnd),
	.combout(\Mux14~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~11 .lut_mask = 16'hDDA0;
defparam \Mux14~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N30
cycloneive_lcell_comb \Reg[14][17]~feeder (
// Equation(s):
// \Reg[14][17]~feeder_combout  = \wdat~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat31),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[14][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[14][17]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[14][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N31
dffeas \Reg[14][17] (
	.clk(!CLK),
	.d(\Reg[14][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[14][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[14][17] .is_wysiwyg = "true";
defparam \Reg[14][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N16
cycloneive_lcell_comb \Reg[15][17]~feeder (
// Equation(s):
// \Reg[15][17]~feeder_combout  = \wdat~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat31),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[15][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[15][17]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[15][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N17
dffeas \Reg[15][17] (
	.clk(!CLK),
	.d(\Reg[15][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[15][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[15][17] .is_wysiwyg = "true";
defparam \Reg[15][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N19
dffeas \Reg[12][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][17] .is_wysiwyg = "true";
defparam \Reg[12][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N17
dffeas \Reg[13][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][17] .is_wysiwyg = "true";
defparam \Reg[13][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N16
cycloneive_lcell_comb \Mux14~17 (
// Equation(s):
// \Mux14~17_combout  = (ifid_ifinstr_o_21 & (((\Reg[13][17]~q ) # (ifid_ifinstr_o_22)))) # (!ifid_ifinstr_o_21 & (\Reg[12][17]~q  & ((!ifid_ifinstr_o_22))))

	.dataa(ifid_ifinstr_o_21),
	.datab(\Reg[12][17]~q ),
	.datac(\Reg[13][17]~q ),
	.datad(ifid_ifinstr_o_22),
	.cin(gnd),
	.combout(\Mux14~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~17 .lut_mask = 16'hAAE4;
defparam \Mux14~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N14
cycloneive_lcell_comb \Mux14~18 (
// Equation(s):
// \Mux14~18_combout  = (ifid_ifinstr_o_22 & ((\Mux14~17_combout  & ((\Reg[15][17]~q ))) # (!\Mux14~17_combout  & (\Reg[14][17]~q )))) # (!ifid_ifinstr_o_22 & (((\Mux14~17_combout ))))

	.dataa(\Reg[14][17]~q ),
	.datab(ifid_ifinstr_o_22),
	.datac(\Reg[15][17]~q ),
	.datad(\Mux14~17_combout ),
	.cin(gnd),
	.combout(\Mux14~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~18 .lut_mask = 16'hF388;
defparam \Mux14~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N26
cycloneive_lcell_comb \Mux32~0 (
// Equation(s):
// \Mux32~0_combout  = (ifid_ifinstr_o_19 & ((\Reg[25][31]~q ) # ((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & (((!ifid_ifinstr_o_18 & \Reg[17][31]~q ))))

	.dataa(\Reg[25][31]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(ifid_ifinstr_o_18),
	.datad(\Reg[17][31]~q ),
	.cin(gnd),
	.combout(\Mux32~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~0 .lut_mask = 16'hCBC8;
defparam \Mux32~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N24
cycloneive_lcell_comb \Mux32~1 (
// Equation(s):
// \Mux32~1_combout  = (\Mux32~0_combout  & (((\Reg[29][31]~q )) # (!ifid_ifinstr_o_18))) # (!\Mux32~0_combout  & (ifid_ifinstr_o_18 & (\Reg[21][31]~q )))

	.dataa(\Mux32~0_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[21][31]~q ),
	.datad(\Reg[29][31]~q ),
	.cin(gnd),
	.combout(\Mux32~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~1 .lut_mask = 16'hEA62;
defparam \Mux32~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y34_N27
dffeas \Reg[30][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][31] .is_wysiwyg = "true";
defparam \Reg[30][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N26
cycloneive_lcell_comb \Mux32~3 (
// Equation(s):
// \Mux32~3_combout  = (\Mux32~2_combout  & (((\Reg[30][31]~q ) # (!ifid_ifinstr_o_19)))) # (!\Mux32~2_combout  & (\Reg[26][31]~q  & ((ifid_ifinstr_o_19))))

	.dataa(\Mux32~2_combout ),
	.datab(\Reg[26][31]~q ),
	.datac(\Reg[30][31]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux32~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~3 .lut_mask = 16'hE4AA;
defparam \Mux32~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y32_N19
dffeas \Reg[16][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][31] .is_wysiwyg = "true";
defparam \Reg[16][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N18
cycloneive_lcell_comb \Mux32~4 (
// Equation(s):
// \Mux32~4_combout  = (ifid_ifinstr_o_18 & ((\Reg[20][31]~q ) # ((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (((\Reg[16][31]~q  & !ifid_ifinstr_o_19))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[20][31]~q ),
	.datac(\Reg[16][31]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux32~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~4 .lut_mask = 16'hAAD8;
defparam \Mux32~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N18
cycloneive_lcell_comb \Mux32~5 (
// Equation(s):
// \Mux32~5_combout  = (ifid_ifinstr_o_19 & ((\Mux32~4_combout  & ((\Reg[28][31]~q ))) # (!\Mux32~4_combout  & (\Reg[24][31]~q )))) # (!ifid_ifinstr_o_19 & (((\Mux32~4_combout ))))

	.dataa(\Reg[24][31]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[28][31]~q ),
	.datad(\Mux32~4_combout ),
	.cin(gnd),
	.combout(\Mux32~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~5 .lut_mask = 16'hF388;
defparam \Mux32~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N22
cycloneive_lcell_comb \Mux32~6 (
// Equation(s):
// \Mux32~6_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Mux32~3_combout )) # (!ifid_ifinstr_o_17 & ((\Mux32~5_combout )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux32~3_combout ),
	.datad(\Mux32~5_combout ),
	.cin(gnd),
	.combout(\Mux32~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~6 .lut_mask = 16'hD9C8;
defparam \Mux32~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N11
dffeas \Reg[19][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat17),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][31] .is_wysiwyg = "true";
defparam \Reg[19][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N10
cycloneive_lcell_comb \Mux32~7 (
// Equation(s):
// \Mux32~7_combout  = (ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18) # ((\Reg[27][31]~q )))) # (!ifid_ifinstr_o_19 & (!ifid_ifinstr_o_18 & (\Reg[19][31]~q )))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[19][31]~q ),
	.datad(\Reg[27][31]~q ),
	.cin(gnd),
	.combout(\Mux32~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~7 .lut_mask = 16'hBA98;
defparam \Mux32~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N22
cycloneive_lcell_comb \Mux32~8 (
// Equation(s):
// \Mux32~8_combout  = (ifid_ifinstr_o_18 & ((\Mux32~7_combout  & (\Reg[31][31]~q )) # (!\Mux32~7_combout  & ((\Reg[23][31]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux32~7_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[31][31]~q ),
	.datac(\Reg[23][31]~q ),
	.datad(\Mux32~7_combout ),
	.cin(gnd),
	.combout(\Mux32~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~8 .lut_mask = 16'hDDA0;
defparam \Mux32~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N4
cycloneive_lcell_comb \Mux32~17 (
// Equation(s):
// \Mux32~17_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[13][31]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[12][31]~q )))))

	.dataa(\Reg[13][31]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[12][31]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux32~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~17 .lut_mask = 16'hEE30;
defparam \Mux32~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N30
cycloneive_lcell_comb \Mux32~18 (
// Equation(s):
// \Mux32~18_combout  = (\Mux32~17_combout  & (((\Reg[15][31]~q ) # (!ifid_ifinstr_o_17)))) # (!\Mux32~17_combout  & (\Reg[14][31]~q  & ((ifid_ifinstr_o_17))))

	.dataa(\Mux32~17_combout ),
	.datab(\Reg[14][31]~q ),
	.datac(\Reg[15][31]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux32~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~18 .lut_mask = 16'hE4AA;
defparam \Mux32~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N0
cycloneive_lcell_comb \Mux32~10 (
// Equation(s):
// \Mux32~10_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17) # ((\Reg[5][31]~q )))) # (!ifid_ifinstr_o_16 & (!ifid_ifinstr_o_17 & ((\Reg[4][31]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[5][31]~q ),
	.datad(\Reg[4][31]~q ),
	.cin(gnd),
	.combout(\Mux32~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~10 .lut_mask = 16'hB9A8;
defparam \Mux32~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N24
cycloneive_lcell_comb \Mux32~11 (
// Equation(s):
// \Mux32~11_combout  = (\Mux32~10_combout  & ((\Reg[7][31]~q ) # ((!ifid_ifinstr_o_17)))) # (!\Mux32~10_combout  & (((\Reg[6][31]~q  & ifid_ifinstr_o_17))))

	.dataa(\Reg[7][31]~q ),
	.datab(\Mux32~10_combout ),
	.datac(\Reg[6][31]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux32~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~11 .lut_mask = 16'hB8CC;
defparam \Mux32~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N30
cycloneive_lcell_comb \Mux32~15 (
// Equation(s):
// \Mux32~15_combout  = (\Mux32~14_combout ) # ((ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & \Reg[2][31]~q )))

	.dataa(\Mux32~14_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(ifid_ifinstr_o_16),
	.datad(\Reg[2][31]~q ),
	.cin(gnd),
	.combout(\Mux32~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~15 .lut_mask = 16'hAEAA;
defparam \Mux32~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N10
cycloneive_lcell_comb \Mux32~13 (
// Equation(s):
// \Mux32~13_combout  = (\Mux32~12_combout  & (((\Reg[11][31]~q ) # (!ifid_ifinstr_o_16)))) # (!\Mux32~12_combout  & (\Reg[9][31]~q  & ((ifid_ifinstr_o_16))))

	.dataa(\Mux32~12_combout ),
	.datab(\Reg[9][31]~q ),
	.datac(\Reg[11][31]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux32~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~13 .lut_mask = 16'hE4AA;
defparam \Mux32~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N0
cycloneive_lcell_comb \Mux32~16 (
// Equation(s):
// \Mux32~16_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Mux32~13_combout ))) # (!ifid_ifinstr_o_19 & (\Mux32~15_combout ))))

	.dataa(\Mux32~15_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux32~13_combout ),
	.cin(gnd),
	.combout(\Mux32~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~16 .lut_mask = 16'hF2C2;
defparam \Mux32~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y30_N23
dffeas \Reg[18][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][16] .is_wysiwyg = "true";
defparam \Reg[18][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N22
cycloneive_lcell_comb \Mux47~2 (
// Equation(s):
// \Mux47~2_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[26][16]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[18][16]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[18][16]~q ),
	.datad(\Reg[26][16]~q ),
	.cin(gnd),
	.combout(\Mux47~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~2 .lut_mask = 16'hDC98;
defparam \Mux47~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N3
dffeas \Reg[22][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][16] .is_wysiwyg = "true";
defparam \Reg[22][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N24
cycloneive_lcell_comb \Mux47~3 (
// Equation(s):
// \Mux47~3_combout  = (ifid_ifinstr_o_18 & ((\Mux47~2_combout  & (\Reg[30][16]~q )) # (!\Mux47~2_combout  & ((\Reg[22][16]~q ))))) # (!ifid_ifinstr_o_18 & (\Mux47~2_combout ))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux47~2_combout ),
	.datac(\Reg[30][16]~q ),
	.datad(\Reg[22][16]~q ),
	.cin(gnd),
	.combout(\Mux47~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~3 .lut_mask = 16'hE6C4;
defparam \Mux47~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N25
dffeas \Reg[20][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat9),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][16] .is_wysiwyg = "true";
defparam \Reg[20][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N4
cycloneive_lcell_comb \Mux47~4 (
// Equation(s):
// \Mux47~4_combout  = (ifid_ifinstr_o_19 & (((\Reg[24][16]~q ) # (ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & (\Reg[16][16]~q  & ((!ifid_ifinstr_o_18))))

	.dataa(\Reg[16][16]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[24][16]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux47~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~4 .lut_mask = 16'hCCE2;
defparam \Mux47~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N24
cycloneive_lcell_comb \Mux47~5 (
// Equation(s):
// \Mux47~5_combout  = (ifid_ifinstr_o_18 & ((\Mux47~4_combout  & (\Reg[28][16]~q )) # (!\Mux47~4_combout  & ((\Reg[20][16]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux47~4_combout ))))

	.dataa(\Reg[28][16]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[20][16]~q ),
	.datad(\Mux47~4_combout ),
	.cin(gnd),
	.combout(\Mux47~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~5 .lut_mask = 16'hBBC0;
defparam \Mux47~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N26
cycloneive_lcell_comb \Mux47~6 (
// Equation(s):
// \Mux47~6_combout  = (ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16) # ((\Mux47~3_combout )))) # (!ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & ((\Mux47~5_combout ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux47~3_combout ),
	.datad(\Mux47~5_combout ),
	.cin(gnd),
	.combout(\Mux47~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~6 .lut_mask = 16'hB9A8;
defparam \Mux47~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N30
cycloneive_lcell_comb \Mux47~7 (
// Equation(s):
// \Mux47~7_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Reg[23][16]~q ))) # (!ifid_ifinstr_o_18 & (\Reg[19][16]~q ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[19][16]~q ),
	.datad(\Reg[23][16]~q ),
	.cin(gnd),
	.combout(\Mux47~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~7 .lut_mask = 16'hDC98;
defparam \Mux47~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N14
cycloneive_lcell_comb \Mux47~8 (
// Equation(s):
// \Mux47~8_combout  = (ifid_ifinstr_o_19 & ((\Mux47~7_combout  & ((\Reg[31][16]~q ))) # (!\Mux47~7_combout  & (\Reg[27][16]~q )))) # (!ifid_ifinstr_o_19 & (((\Mux47~7_combout ))))

	.dataa(\Reg[27][16]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[31][16]~q ),
	.datad(\Mux47~7_combout ),
	.cin(gnd),
	.combout(\Mux47~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~8 .lut_mask = 16'hF388;
defparam \Mux47~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N26
cycloneive_lcell_comb \Mux47~0 (
// Equation(s):
// \Mux47~0_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[21][16]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[17][16]~q )))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[21][16]~q ),
	.datad(\Reg[17][16]~q ),
	.cin(gnd),
	.combout(\Mux47~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~0 .lut_mask = 16'hD9C8;
defparam \Mux47~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N8
cycloneive_lcell_comb \Mux47~1 (
// Equation(s):
// \Mux47~1_combout  = (ifid_ifinstr_o_19 & ((\Mux47~0_combout  & (\Reg[29][16]~q )) # (!\Mux47~0_combout  & ((\Reg[25][16]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux47~0_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[29][16]~q ),
	.datac(\Mux47~0_combout ),
	.datad(\Reg[25][16]~q ),
	.cin(gnd),
	.combout(\Mux47~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~1 .lut_mask = 16'hDAD0;
defparam \Mux47~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N2
cycloneive_lcell_comb \Mux47~17 (
// Equation(s):
// \Mux47~17_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17) # ((\Reg[13][16]~q )))) # (!ifid_ifinstr_o_16 & (!ifid_ifinstr_o_17 & ((\Reg[12][16]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[13][16]~q ),
	.datad(\Reg[12][16]~q ),
	.cin(gnd),
	.combout(\Mux47~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~17 .lut_mask = 16'hB9A8;
defparam \Mux47~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N22
cycloneive_lcell_comb \Mux47~18 (
// Equation(s):
// \Mux47~18_combout  = (ifid_ifinstr_o_17 & ((\Mux47~17_combout  & ((\Reg[15][16]~q ))) # (!\Mux47~17_combout  & (\Reg[14][16]~q )))) # (!ifid_ifinstr_o_17 & (((\Mux47~17_combout ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[14][16]~q ),
	.datac(\Reg[15][16]~q ),
	.datad(\Mux47~17_combout ),
	.cin(gnd),
	.combout(\Mux47~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~18 .lut_mask = 16'hF588;
defparam \Mux47~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N20
cycloneive_lcell_comb \Mux47~10 (
// Equation(s):
// \Mux47~10_combout  = (ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16) # ((\Reg[10][16]~q )))) # (!ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & ((\Reg[8][16]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[10][16]~q ),
	.datad(\Reg[8][16]~q ),
	.cin(gnd),
	.combout(\Mux47~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~10 .lut_mask = 16'hB9A8;
defparam \Mux47~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N2
cycloneive_lcell_comb \Mux47~11 (
// Equation(s):
// \Mux47~11_combout  = (\Mux47~10_combout  & ((\Reg[11][16]~q ) # ((!ifid_ifinstr_o_16)))) # (!\Mux47~10_combout  & (((\Reg[9][16]~q  & ifid_ifinstr_o_16))))

	.dataa(\Mux47~10_combout ),
	.datab(\Reg[11][16]~q ),
	.datac(\Reg[9][16]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux47~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~11 .lut_mask = 16'hD8AA;
defparam \Mux47~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N20
cycloneive_lcell_comb \Mux47~14 (
// Equation(s):
// \Mux47~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][16]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][16]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[3][16]~q ),
	.datad(\Reg[1][16]~q ),
	.cin(gnd),
	.combout(\Mux47~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~14 .lut_mask = 16'hA280;
defparam \Mux47~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N14
cycloneive_lcell_comb \Mux47~15 (
// Equation(s):
// \Mux47~15_combout  = (\Mux47~14_combout ) # ((ifid_ifinstr_o_17 & (\Reg[2][16]~q  & !ifid_ifinstr_o_16)))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[2][16]~q ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux47~14_combout ),
	.cin(gnd),
	.combout(\Mux47~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~15 .lut_mask = 16'hFF08;
defparam \Mux47~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N22
cycloneive_lcell_comb \Mux47~13 (
// Equation(s):
// \Mux47~13_combout  = (\Mux47~12_combout  & (((\Reg[7][16]~q )) # (!ifid_ifinstr_o_17))) # (!\Mux47~12_combout  & (ifid_ifinstr_o_17 & ((\Reg[6][16]~q ))))

	.dataa(\Mux47~12_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[7][16]~q ),
	.datad(\Reg[6][16]~q ),
	.cin(gnd),
	.combout(\Mux47~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~13 .lut_mask = 16'hE6A2;
defparam \Mux47~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N0
cycloneive_lcell_comb \Mux47~16 (
// Equation(s):
// \Mux47~16_combout  = (ifid_ifinstr_o_19 & (((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Mux47~13_combout ))) # (!ifid_ifinstr_o_18 & (\Mux47~15_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Mux47~15_combout ),
	.datac(ifid_ifinstr_o_18),
	.datad(\Mux47~13_combout ),
	.cin(gnd),
	.combout(\Mux47~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~16 .lut_mask = 16'hF4A4;
defparam \Mux47~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N16
cycloneive_lcell_comb \Mux46~7 (
// Equation(s):
// \Mux46~7_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[27][17]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[19][17]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[19][17]~q ),
	.datac(\Reg[27][17]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux46~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~7 .lut_mask = 16'hFA44;
defparam \Mux46~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N6
cycloneive_lcell_comb \Mux46~8 (
// Equation(s):
// \Mux46~8_combout  = (ifid_ifinstr_o_18 & ((\Mux46~7_combout  & (\Reg[31][17]~q )) # (!\Mux46~7_combout  & ((\Reg[23][17]~q ))))) # (!ifid_ifinstr_o_18 & (\Mux46~7_combout ))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux46~7_combout ),
	.datac(\Reg[31][17]~q ),
	.datad(\Reg[23][17]~q ),
	.cin(gnd),
	.combout(\Mux46~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~8 .lut_mask = 16'hE6C4;
defparam \Mux46~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N28
cycloneive_lcell_comb \Mux46~0 (
// Equation(s):
// \Mux46~0_combout  = (ifid_ifinstr_o_19 & ((\Reg[25][17]~q ) # ((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & (((\Reg[17][17]~q  & !ifid_ifinstr_o_18))))

	.dataa(\Reg[25][17]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[17][17]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux46~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~0 .lut_mask = 16'hCCB8;
defparam \Mux46~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N4
cycloneive_lcell_comb \Mux46~1 (
// Equation(s):
// \Mux46~1_combout  = (ifid_ifinstr_o_18 & ((\Mux46~0_combout  & ((\Reg[29][17]~q ))) # (!\Mux46~0_combout  & (\Reg[21][17]~q )))) # (!ifid_ifinstr_o_18 & (((\Mux46~0_combout ))))

	.dataa(\Reg[21][17]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[29][17]~q ),
	.datad(\Mux46~0_combout ),
	.cin(gnd),
	.combout(\Mux46~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~1 .lut_mask = 16'hF388;
defparam \Mux46~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N18
cycloneive_lcell_comb \Reg[20][17]~feeder (
// Equation(s):
// \Reg[20][17]~feeder_combout  = \wdat~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat31),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[20][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[20][17]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[20][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N19
dffeas \Reg[20][17] (
	.clk(!CLK),
	.d(\Reg[20][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][17] .is_wysiwyg = "true";
defparam \Reg[20][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N20
cycloneive_lcell_comb \Mux46~4 (
// Equation(s):
// \Mux46~4_combout  = (ifid_ifinstr_o_18 & ((\Reg[20][17]~q ) # ((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (((\Reg[16][17]~q  & !ifid_ifinstr_o_19))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[20][17]~q ),
	.datac(\Reg[16][17]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux46~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~4 .lut_mask = 16'hAAD8;
defparam \Mux46~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N6
cycloneive_lcell_comb \Mux46~5 (
// Equation(s):
// \Mux46~5_combout  = (ifid_ifinstr_o_19 & ((\Mux46~4_combout  & (\Reg[28][17]~q )) # (!\Mux46~4_combout  & ((\Reg[24][17]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux46~4_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[28][17]~q ),
	.datac(\Mux46~4_combout ),
	.datad(\Reg[24][17]~q ),
	.cin(gnd),
	.combout(\Mux46~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~5 .lut_mask = 16'hDAD0;
defparam \Mux46~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N16
cycloneive_lcell_comb \Reg[30][17]~feeder (
// Equation(s):
// \Reg[30][17]~feeder_combout  = \wdat~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat31),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[30][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[30][17]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[30][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N17
dffeas \Reg[30][17] (
	.clk(!CLK),
	.d(\Reg[30][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][17] .is_wysiwyg = "true";
defparam \Reg[30][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N10
cycloneive_lcell_comb \Mux46~2 (
// Equation(s):
// \Mux46~2_combout  = (ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19) # ((\Reg[22][17]~q )))) # (!ifid_ifinstr_o_18 & (!ifid_ifinstr_o_19 & (\Reg[18][17]~q )))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[18][17]~q ),
	.datad(\Reg[22][17]~q ),
	.cin(gnd),
	.combout(\Mux46~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~2 .lut_mask = 16'hBA98;
defparam \Mux46~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N12
cycloneive_lcell_comb \Mux46~3 (
// Equation(s):
// \Mux46~3_combout  = (ifid_ifinstr_o_19 & ((\Mux46~2_combout  & (\Reg[30][17]~q )) # (!\Mux46~2_combout  & ((\Reg[26][17]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux46~2_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[30][17]~q ),
	.datac(\Reg[26][17]~q ),
	.datad(\Mux46~2_combout ),
	.cin(gnd),
	.combout(\Mux46~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~3 .lut_mask = 16'hDDA0;
defparam \Mux46~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N10
cycloneive_lcell_comb \Mux46~6 (
// Equation(s):
// \Mux46~6_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Mux46~3_combout ))) # (!ifid_ifinstr_o_17 & (\Mux46~5_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux46~5_combout ),
	.datad(\Mux46~3_combout ),
	.cin(gnd),
	.combout(\Mux46~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~6 .lut_mask = 16'hDC98;
defparam \Mux46~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N18
cycloneive_lcell_comb \Mux46~17 (
// Equation(s):
// \Mux46~17_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[13][17]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[12][17]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[13][17]~q ),
	.datac(\Reg[12][17]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux46~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~17 .lut_mask = 16'hEE50;
defparam \Mux46~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N6
cycloneive_lcell_comb \Mux46~18 (
// Equation(s):
// \Mux46~18_combout  = (\Mux46~17_combout  & (((\Reg[15][17]~q ) # (!ifid_ifinstr_o_17)))) # (!\Mux46~17_combout  & (\Reg[14][17]~q  & ((ifid_ifinstr_o_17))))

	.dataa(\Reg[14][17]~q ),
	.datab(\Reg[15][17]~q ),
	.datac(\Mux46~17_combout ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux46~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~18 .lut_mask = 16'hCAF0;
defparam \Mux46~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N20
cycloneive_lcell_comb \Mux46~15 (
// Equation(s):
// \Mux46~15_combout  = (\Mux46~14_combout ) # ((!ifid_ifinstr_o_16 & (\Reg[2][17]~q  & ifid_ifinstr_o_17)))

	.dataa(\Mux46~14_combout ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[2][17]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux46~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~15 .lut_mask = 16'hBAAA;
defparam \Mux46~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N2
cycloneive_lcell_comb \Mux46~12 (
// Equation(s):
// \Mux46~12_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[10][17]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[8][17]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[8][17]~q ),
	.datad(\Reg[10][17]~q ),
	.cin(gnd),
	.combout(\Mux46~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~12 .lut_mask = 16'hDC98;
defparam \Mux46~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N28
cycloneive_lcell_comb \Mux46~13 (
// Equation(s):
// \Mux46~13_combout  = (ifid_ifinstr_o_16 & ((\Mux46~12_combout  & ((\Reg[11][17]~q ))) # (!\Mux46~12_combout  & (\Reg[9][17]~q )))) # (!ifid_ifinstr_o_16 & (((\Mux46~12_combout ))))

	.dataa(\Reg[9][17]~q ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[11][17]~q ),
	.datad(\Mux46~12_combout ),
	.cin(gnd),
	.combout(\Mux46~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~13 .lut_mask = 16'hF388;
defparam \Mux46~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N22
cycloneive_lcell_comb \Mux46~16 (
// Equation(s):
// \Mux46~16_combout  = (ifid_ifinstr_o_19 & (((ifid_ifinstr_o_18) # (\Mux46~13_combout )))) # (!ifid_ifinstr_o_19 & (\Mux46~15_combout  & (!ifid_ifinstr_o_18)))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Mux46~15_combout ),
	.datac(ifid_ifinstr_o_18),
	.datad(\Mux46~13_combout ),
	.cin(gnd),
	.combout(\Mux46~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~16 .lut_mask = 16'hAEA4;
defparam \Mux46~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y39_N13
dffeas \Reg[5][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][17] .is_wysiwyg = "true";
defparam \Reg[5][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y39_N3
dffeas \Reg[4][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat31),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][17] .is_wysiwyg = "true";
defparam \Reg[4][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N12
cycloneive_lcell_comb \Mux46~10 (
// Equation(s):
// \Mux46~10_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[5][17]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[4][17]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[5][17]~q ),
	.datad(\Reg[4][17]~q ),
	.cin(gnd),
	.combout(\Mux46~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~10 .lut_mask = 16'hD9C8;
defparam \Mux46~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N8
cycloneive_lcell_comb \Mux46~11 (
// Equation(s):
// \Mux46~11_combout  = (\Mux46~10_combout  & ((\Reg[7][17]~q ) # ((!ifid_ifinstr_o_17)))) # (!\Mux46~10_combout  & (((\Reg[6][17]~q  & ifid_ifinstr_o_17))))

	.dataa(\Reg[7][17]~q ),
	.datab(\Mux46~10_combout ),
	.datac(\Reg[6][17]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux46~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~11 .lut_mask = 16'hB8CC;
defparam \Mux46~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N3
dffeas \Reg[20][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][18] .is_wysiwyg = "true";
defparam \Reg[20][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y32_N29
dffeas \Reg[16][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat29),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][18] .is_wysiwyg = "true";
defparam \Reg[16][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N26
cycloneive_lcell_comb \Mux45~4 (
// Equation(s):
// \Mux45~4_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[24][18]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[16][18]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[16][18]~q ),
	.datac(\Reg[24][18]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux45~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~4 .lut_mask = 16'hFA44;
defparam \Mux45~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N2
cycloneive_lcell_comb \Mux45~5 (
// Equation(s):
// \Mux45~5_combout  = (ifid_ifinstr_o_18 & ((\Mux45~4_combout  & (\Reg[28][18]~q )) # (!\Mux45~4_combout  & ((\Reg[20][18]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux45~4_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[28][18]~q ),
	.datac(\Reg[20][18]~q ),
	.datad(\Mux45~4_combout ),
	.cin(gnd),
	.combout(\Mux45~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~5 .lut_mask = 16'hDDA0;
defparam \Mux45~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N16
cycloneive_lcell_comb \Mux45~2 (
// Equation(s):
// \Mux45~2_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[26][18]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[18][18]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[18][18]~q ),
	.datac(\Reg[26][18]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux45~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~2 .lut_mask = 16'hFA44;
defparam \Mux45~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N6
cycloneive_lcell_comb \Mux45~3 (
// Equation(s):
// \Mux45~3_combout  = (ifid_ifinstr_o_18 & ((\Mux45~2_combout  & ((\Reg[30][18]~q ))) # (!\Mux45~2_combout  & (\Reg[22][18]~q )))) # (!ifid_ifinstr_o_18 & (((\Mux45~2_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[22][18]~q ),
	.datac(\Reg[30][18]~q ),
	.datad(\Mux45~2_combout ),
	.cin(gnd),
	.combout(\Mux45~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~3 .lut_mask = 16'hF588;
defparam \Mux45~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N6
cycloneive_lcell_comb \Mux45~6 (
// Equation(s):
// \Mux45~6_combout  = (ifid_ifinstr_o_17 & (((\Mux45~3_combout ) # (ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & (\Mux45~5_combout  & ((!ifid_ifinstr_o_16))))

	.dataa(\Mux45~5_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux45~3_combout ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux45~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~6 .lut_mask = 16'hCCE2;
defparam \Mux45~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N28
cycloneive_lcell_comb \Mux45~7 (
// Equation(s):
// \Mux45~7_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[23][18]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[19][18]~q )))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[23][18]~q ),
	.datad(\Reg[19][18]~q ),
	.cin(gnd),
	.combout(\Mux45~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~7 .lut_mask = 16'hD9C8;
defparam \Mux45~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N30
cycloneive_lcell_comb \Mux45~8 (
// Equation(s):
// \Mux45~8_combout  = (\Mux45~7_combout  & ((\Reg[31][18]~q ) # ((!ifid_ifinstr_o_19)))) # (!\Mux45~7_combout  & (((ifid_ifinstr_o_19 & \Reg[27][18]~q ))))

	.dataa(\Mux45~7_combout ),
	.datab(\Reg[31][18]~q ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Reg[27][18]~q ),
	.cin(gnd),
	.combout(\Mux45~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~8 .lut_mask = 16'hDA8A;
defparam \Mux45~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N28
cycloneive_lcell_comb \Mux45~0 (
// Equation(s):
// \Mux45~0_combout  = (ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19) # ((\Reg[21][18]~q )))) # (!ifid_ifinstr_o_18 & (!ifid_ifinstr_o_19 & (\Reg[17][18]~q )))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[17][18]~q ),
	.datad(\Reg[21][18]~q ),
	.cin(gnd),
	.combout(\Mux45~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~0 .lut_mask = 16'hBA98;
defparam \Mux45~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N20
cycloneive_lcell_comb \Mux45~1 (
// Equation(s):
// \Mux45~1_combout  = (ifid_ifinstr_o_19 & ((\Mux45~0_combout  & ((\Reg[29][18]~q ))) # (!\Mux45~0_combout  & (\Reg[25][18]~q )))) # (!ifid_ifinstr_o_19 & (((\Mux45~0_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[25][18]~q ),
	.datac(\Reg[29][18]~q ),
	.datad(\Mux45~0_combout ),
	.cin(gnd),
	.combout(\Mux45~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~1 .lut_mask = 16'hF588;
defparam \Mux45~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N8
cycloneive_lcell_comb \Mux45~10 (
// Equation(s):
// \Mux45~10_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[10][18]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[8][18]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[10][18]~q ),
	.datad(\Reg[8][18]~q ),
	.cin(gnd),
	.combout(\Mux45~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~10 .lut_mask = 16'hD9C8;
defparam \Mux45~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N10
cycloneive_lcell_comb \Mux45~11 (
// Equation(s):
// \Mux45~11_combout  = (\Mux45~10_combout  & ((\Reg[11][18]~q ) # ((!ifid_ifinstr_o_16)))) # (!\Mux45~10_combout  & (((\Reg[9][18]~q  & ifid_ifinstr_o_16))))

	.dataa(\Reg[11][18]~q ),
	.datab(\Mux45~10_combout ),
	.datac(\Reg[9][18]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux45~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~11 .lut_mask = 16'hB8CC;
defparam \Mux45~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N24
cycloneive_lcell_comb \Mux45~17 (
// Equation(s):
// \Mux45~17_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[13][18]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[12][18]~q ))))

	.dataa(\Reg[12][18]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[13][18]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux45~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~17 .lut_mask = 16'hFC22;
defparam \Mux45~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N12
cycloneive_lcell_comb \Mux45~18 (
// Equation(s):
// \Mux45~18_combout  = (ifid_ifinstr_o_17 & ((\Mux45~17_combout  & ((\Reg[15][18]~q ))) # (!\Mux45~17_combout  & (\Reg[14][18]~q )))) # (!ifid_ifinstr_o_17 & (\Mux45~17_combout ))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux45~17_combout ),
	.datac(\Reg[14][18]~q ),
	.datad(\Reg[15][18]~q ),
	.cin(gnd),
	.combout(\Mux45~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~18 .lut_mask = 16'hEC64;
defparam \Mux45~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N18
cycloneive_lcell_comb \Mux45~13 (
// Equation(s):
// \Mux45~13_combout  = (\Mux45~12_combout  & (((\Reg[7][18]~q ) # (!ifid_ifinstr_o_17)))) # (!\Mux45~12_combout  & (\Reg[6][18]~q  & ((ifid_ifinstr_o_17))))

	.dataa(\Mux45~12_combout ),
	.datab(\Reg[6][18]~q ),
	.datac(\Reg[7][18]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux45~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~13 .lut_mask = 16'hE4AA;
defparam \Mux45~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N30
cycloneive_lcell_comb \Mux45~15 (
// Equation(s):
// \Mux45~15_combout  = (\Mux45~14_combout ) # ((ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & \Reg[2][18]~q )))

	.dataa(\Mux45~14_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(ifid_ifinstr_o_16),
	.datad(\Reg[2][18]~q ),
	.cin(gnd),
	.combout(\Mux45~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~15 .lut_mask = 16'hAEAA;
defparam \Mux45~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N18
cycloneive_lcell_comb \Mux45~16 (
// Equation(s):
// \Mux45~16_combout  = (ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19) # ((\Mux45~13_combout )))) # (!ifid_ifinstr_o_18 & (!ifid_ifinstr_o_19 & ((\Mux45~15_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Mux45~13_combout ),
	.datad(\Mux45~15_combout ),
	.cin(gnd),
	.combout(\Mux45~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~16 .lut_mask = 16'hB9A8;
defparam \Mux45~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N24
cycloneive_lcell_comb \Mux44~0 (
// Equation(s):
// \Mux44~0_combout  = (ifid_ifinstr_o_19 & (((\Reg[25][19]~q ) # (ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & (\Reg[17][19]~q  & ((!ifid_ifinstr_o_18))))

	.dataa(\Reg[17][19]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[25][19]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux44~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~0 .lut_mask = 16'hCCE2;
defparam \Mux44~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N10
cycloneive_lcell_comb \Mux44~1 (
// Equation(s):
// \Mux44~1_combout  = (\Mux44~0_combout  & (((\Reg[29][19]~q )) # (!ifid_ifinstr_o_18))) # (!\Mux44~0_combout  & (ifid_ifinstr_o_18 & (\Reg[21][19]~q )))

	.dataa(\Mux44~0_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[21][19]~q ),
	.datad(\Reg[29][19]~q ),
	.cin(gnd),
	.combout(\Mux44~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~1 .lut_mask = 16'hEA62;
defparam \Mux44~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N6
cycloneive_lcell_comb \Mux44~7 (
// Equation(s):
// \Mux44~7_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[27][19]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[19][19]~q ))))

	.dataa(\Reg[19][19]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[27][19]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux44~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~7 .lut_mask = 16'hFC22;
defparam \Mux44~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N12
cycloneive_lcell_comb \Mux44~8 (
// Equation(s):
// \Mux44~8_combout  = (ifid_ifinstr_o_18 & ((\Mux44~7_combout  & ((\Reg[31][19]~q ))) # (!\Mux44~7_combout  & (\Reg[23][19]~q )))) # (!ifid_ifinstr_o_18 & (((\Mux44~7_combout ))))

	.dataa(\Reg[23][19]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[31][19]~q ),
	.datad(\Mux44~7_combout ),
	.cin(gnd),
	.combout(\Mux44~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~8 .lut_mask = 16'hF388;
defparam \Mux44~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N1
dffeas \Reg[24][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][19] .is_wysiwyg = "true";
defparam \Reg[24][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N6
cycloneive_lcell_comb \Mux44~4 (
// Equation(s):
// \Mux44~4_combout  = (ifid_ifinstr_o_19 & (((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Reg[20][19]~q ))) # (!ifid_ifinstr_o_18 & (\Reg[16][19]~q ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[16][19]~q ),
	.datac(\Reg[20][19]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux44~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~4 .lut_mask = 16'hFA44;
defparam \Mux44~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N0
cycloneive_lcell_comb \Mux44~5 (
// Equation(s):
// \Mux44~5_combout  = (ifid_ifinstr_o_19 & ((\Mux44~4_combout  & (\Reg[28][19]~q )) # (!\Mux44~4_combout  & ((\Reg[24][19]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux44~4_combout ))))

	.dataa(\Reg[28][19]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[24][19]~q ),
	.datad(\Mux44~4_combout ),
	.cin(gnd),
	.combout(\Mux44~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~5 .lut_mask = 16'hBBC0;
defparam \Mux44~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N11
dffeas \Reg[30][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][19] .is_wysiwyg = "true";
defparam \Reg[30][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N31
dffeas \Reg[18][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat30),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][19] .is_wysiwyg = "true";
defparam \Reg[18][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N30
cycloneive_lcell_comb \Mux44~2 (
// Equation(s):
// \Mux44~2_combout  = (ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19) # ((\Reg[22][19]~q )))) # (!ifid_ifinstr_o_18 & (!ifid_ifinstr_o_19 & (\Reg[18][19]~q )))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[18][19]~q ),
	.datad(\Reg[22][19]~q ),
	.cin(gnd),
	.combout(\Mux44~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~2 .lut_mask = 16'hBA98;
defparam \Mux44~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N10
cycloneive_lcell_comb \Mux44~3 (
// Equation(s):
// \Mux44~3_combout  = (ifid_ifinstr_o_19 & ((\Mux44~2_combout  & ((\Reg[30][19]~q ))) # (!\Mux44~2_combout  & (\Reg[26][19]~q )))) # (!ifid_ifinstr_o_19 & (((\Mux44~2_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[26][19]~q ),
	.datac(\Reg[30][19]~q ),
	.datad(\Mux44~2_combout ),
	.cin(gnd),
	.combout(\Mux44~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~3 .lut_mask = 16'hF588;
defparam \Mux44~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N18
cycloneive_lcell_comb \Mux44~6 (
// Equation(s):
// \Mux44~6_combout  = (ifid_ifinstr_o_16 & (((ifid_ifinstr_o_17)))) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Mux44~3_combout ))) # (!ifid_ifinstr_o_17 & (\Mux44~5_combout ))))

	.dataa(\Mux44~5_combout ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux44~3_combout ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux44~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~6 .lut_mask = 16'hFC22;
defparam \Mux44~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N2
cycloneive_lcell_comb \Mux44~12 (
// Equation(s):
// \Mux44~12_combout  = (ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16) # ((\Reg[10][19]~q )))) # (!ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & (\Reg[8][19]~q )))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[8][19]~q ),
	.datad(\Reg[10][19]~q ),
	.cin(gnd),
	.combout(\Mux44~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~12 .lut_mask = 16'hBA98;
defparam \Mux44~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N26
cycloneive_lcell_comb \Mux44~13 (
// Equation(s):
// \Mux44~13_combout  = (ifid_ifinstr_o_16 & ((\Mux44~12_combout  & ((\Reg[11][19]~q ))) # (!\Mux44~12_combout  & (\Reg[9][19]~q )))) # (!ifid_ifinstr_o_16 & (((\Mux44~12_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[9][19]~q ),
	.datac(\Reg[11][19]~q ),
	.datad(\Mux44~12_combout ),
	.cin(gnd),
	.combout(\Mux44~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~13 .lut_mask = 16'hF588;
defparam \Mux44~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N2
cycloneive_lcell_comb \Mux44~14 (
// Equation(s):
// \Mux44~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][19]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][19]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[3][19]~q ),
	.datad(\Reg[1][19]~q ),
	.cin(gnd),
	.combout(\Mux44~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~14 .lut_mask = 16'hA280;
defparam \Mux44~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N6
cycloneive_lcell_comb \Mux44~15 (
// Equation(s):
// \Mux44~15_combout  = (\Mux44~14_combout ) # ((\Reg[2][19]~q  & (ifid_ifinstr_o_17 & !ifid_ifinstr_o_16)))

	.dataa(\Reg[2][19]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux44~14_combout ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux44~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~15 .lut_mask = 16'hF0F8;
defparam \Mux44~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N2
cycloneive_lcell_comb \Mux44~16 (
// Equation(s):
// \Mux44~16_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Mux44~13_combout )) # (!ifid_ifinstr_o_19 & ((\Mux44~15_combout )))))

	.dataa(\Mux44~13_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Mux44~15_combout ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux44~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~16 .lut_mask = 16'hEE30;
defparam \Mux44~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N28
cycloneive_lcell_comb \Mux44~17 (
// Equation(s):
// \Mux44~17_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[13][19]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[12][19]~q ))))

	.dataa(\Reg[12][19]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[13][19]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux44~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~17 .lut_mask = 16'hFC22;
defparam \Mux44~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N0
cycloneive_lcell_comb \Mux44~18 (
// Equation(s):
// \Mux44~18_combout  = (\Mux44~17_combout  & (((\Reg[15][19]~q ) # (!ifid_ifinstr_o_17)))) # (!\Mux44~17_combout  & (\Reg[14][19]~q  & (ifid_ifinstr_o_17)))

	.dataa(\Mux44~17_combout ),
	.datab(\Reg[14][19]~q ),
	.datac(ifid_ifinstr_o_17),
	.datad(\Reg[15][19]~q ),
	.cin(gnd),
	.combout(\Mux44~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~18 .lut_mask = 16'hEA4A;
defparam \Mux44~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N16
cycloneive_lcell_comb \Mux44~10 (
// Equation(s):
// \Mux44~10_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[5][19]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[4][19]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[5][19]~q ),
	.datad(\Reg[4][19]~q ),
	.cin(gnd),
	.combout(\Mux44~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~10 .lut_mask = 16'hD9C8;
defparam \Mux44~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N4
cycloneive_lcell_comb \Mux44~11 (
// Equation(s):
// \Mux44~11_combout  = (ifid_ifinstr_o_17 & ((\Mux44~10_combout  & (\Reg[7][19]~q )) # (!\Mux44~10_combout  & ((\Reg[6][19]~q ))))) # (!ifid_ifinstr_o_17 & (((\Mux44~10_combout ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[7][19]~q ),
	.datac(\Reg[6][19]~q ),
	.datad(\Mux44~10_combout ),
	.cin(gnd),
	.combout(\Mux44~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~11 .lut_mask = 16'hDDA0;
defparam \Mux44~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N8
cycloneive_lcell_comb \Mux43~7 (
// Equation(s):
// \Mux43~7_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[23][20]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[19][20]~q )))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[23][20]~q ),
	.datad(\Reg[19][20]~q ),
	.cin(gnd),
	.combout(\Mux43~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~7 .lut_mask = 16'hD9C8;
defparam \Mux43~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N4
cycloneive_lcell_comb \Mux43~8 (
// Equation(s):
// \Mux43~8_combout  = (\Mux43~7_combout  & (((\Reg[31][20]~q ) # (!ifid_ifinstr_o_19)))) # (!\Mux43~7_combout  & (\Reg[27][20]~q  & (ifid_ifinstr_o_19)))

	.dataa(\Reg[27][20]~q ),
	.datab(\Mux43~7_combout ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Reg[31][20]~q ),
	.cin(gnd),
	.combout(\Mux43~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~8 .lut_mask = 16'hEC2C;
defparam \Mux43~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N26
cycloneive_lcell_comb \Mux43~0 (
// Equation(s):
// \Mux43~0_combout  = (ifid_ifinstr_o_18 & ((\Reg[21][20]~q ) # ((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (((\Reg[17][20]~q  & !ifid_ifinstr_o_19))))

	.dataa(\Reg[21][20]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[17][20]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux43~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~0 .lut_mask = 16'hCCB8;
defparam \Mux43~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y38_N19
dffeas \Reg[25][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][20] .is_wysiwyg = "true";
defparam \Reg[25][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N18
cycloneive_lcell_comb \Mux43~1 (
// Equation(s):
// \Mux43~1_combout  = (\Mux43~0_combout  & ((\Reg[29][20]~q ) # ((!ifid_ifinstr_o_19)))) # (!\Mux43~0_combout  & (((\Reg[25][20]~q  & ifid_ifinstr_o_19))))

	.dataa(\Reg[29][20]~q ),
	.datab(\Mux43~0_combout ),
	.datac(\Reg[25][20]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux43~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~1 .lut_mask = 16'hB8CC;
defparam \Mux43~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N4
cycloneive_lcell_comb \Mux43~2 (
// Equation(s):
// \Mux43~2_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[26][20]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[18][20]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[18][20]~q ),
	.datac(\Reg[26][20]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux43~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~2 .lut_mask = 16'hFA44;
defparam \Mux43~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N2
cycloneive_lcell_comb \Mux43~3 (
// Equation(s):
// \Mux43~3_combout  = (ifid_ifinstr_o_18 & ((\Mux43~2_combout  & (\Reg[30][20]~q )) # (!\Mux43~2_combout  & ((\Reg[22][20]~q ))))) # (!ifid_ifinstr_o_18 & (\Mux43~2_combout ))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux43~2_combout ),
	.datac(\Reg[30][20]~q ),
	.datad(\Reg[22][20]~q ),
	.cin(gnd),
	.combout(\Mux43~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~3 .lut_mask = 16'hE6C4;
defparam \Mux43~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y32_N11
dffeas \Reg[24][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][20] .is_wysiwyg = "true";
defparam \Reg[24][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N10
cycloneive_lcell_comb \Mux43~4 (
// Equation(s):
// \Mux43~4_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[24][20]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[16][20]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[16][20]~q ),
	.datac(\Reg[24][20]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux43~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~4 .lut_mask = 16'hFA44;
defparam \Mux43~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N15
dffeas \Reg[20][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat28),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][20] .is_wysiwyg = "true";
defparam \Reg[20][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N14
cycloneive_lcell_comb \Mux43~5 (
// Equation(s):
// \Mux43~5_combout  = (ifid_ifinstr_o_18 & ((\Mux43~4_combout  & ((\Reg[28][20]~q ))) # (!\Mux43~4_combout  & (\Reg[20][20]~q )))) # (!ifid_ifinstr_o_18 & (\Mux43~4_combout ))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux43~4_combout ),
	.datac(\Reg[20][20]~q ),
	.datad(\Reg[28][20]~q ),
	.cin(gnd),
	.combout(\Mux43~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~5 .lut_mask = 16'hEC64;
defparam \Mux43~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N12
cycloneive_lcell_comb \Mux43~6 (
// Equation(s):
// \Mux43~6_combout  = (ifid_ifinstr_o_16 & (((ifid_ifinstr_o_17)))) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Mux43~3_combout )) # (!ifid_ifinstr_o_17 & ((\Mux43~5_combout )))))

	.dataa(\Mux43~3_combout ),
	.datab(\Mux43~5_combout ),
	.datac(ifid_ifinstr_o_16),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux43~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~6 .lut_mask = 16'hFA0C;
defparam \Mux43~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N14
cycloneive_lcell_comb \Mux43~17 (
// Equation(s):
// \Mux43~17_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[13][20]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[12][20]~q )))))

	.dataa(\Reg[13][20]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[12][20]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux43~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~17 .lut_mask = 16'hEE30;
defparam \Mux43~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N20
cycloneive_lcell_comb \Mux43~18 (
// Equation(s):
// \Mux43~18_combout  = (\Mux43~17_combout  & ((\Reg[15][20]~q ) # ((!ifid_ifinstr_o_17)))) # (!\Mux43~17_combout  & (((\Reg[14][20]~q  & ifid_ifinstr_o_17))))

	.dataa(\Mux43~17_combout ),
	.datab(\Reg[15][20]~q ),
	.datac(\Reg[14][20]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux43~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~18 .lut_mask = 16'hD8AA;
defparam \Mux43~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N20
cycloneive_lcell_comb \Mux43~10 (
// Equation(s):
// \Mux43~10_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[10][20]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[8][20]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[10][20]~q ),
	.datad(\Reg[8][20]~q ),
	.cin(gnd),
	.combout(\Mux43~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~10 .lut_mask = 16'hD9C8;
defparam \Mux43~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N14
cycloneive_lcell_comb \Mux43~11 (
// Equation(s):
// \Mux43~11_combout  = (\Mux43~10_combout  & ((\Reg[11][20]~q ) # ((!ifid_ifinstr_o_16)))) # (!\Mux43~10_combout  & (((\Reg[9][20]~q  & ifid_ifinstr_o_16))))

	.dataa(\Mux43~10_combout ),
	.datab(\Reg[11][20]~q ),
	.datac(\Reg[9][20]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux43~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~11 .lut_mask = 16'hD8AA;
defparam \Mux43~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N14
cycloneive_lcell_comb \Mux43~15 (
// Equation(s):
// \Mux43~15_combout  = (\Mux43~14_combout ) # ((!ifid_ifinstr_o_16 & (\Reg[2][20]~q  & ifid_ifinstr_o_17)))

	.dataa(\Mux43~14_combout ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[2][20]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux43~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~15 .lut_mask = 16'hBAAA;
defparam \Mux43~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N28
cycloneive_lcell_comb \Mux43~13 (
// Equation(s):
// \Mux43~13_combout  = (\Mux43~12_combout  & (((\Reg[7][20]~q ) # (!ifid_ifinstr_o_17)))) # (!\Mux43~12_combout  & (\Reg[6][20]~q  & ((ifid_ifinstr_o_17))))

	.dataa(\Mux43~12_combout ),
	.datab(\Reg[6][20]~q ),
	.datac(\Reg[7][20]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux43~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~13 .lut_mask = 16'hE4AA;
defparam \Mux43~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N24
cycloneive_lcell_comb \Mux43~16 (
// Equation(s):
// \Mux43~16_combout  = (ifid_ifinstr_o_18 & (((\Mux43~13_combout ) # (ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (\Mux43~15_combout  & ((!ifid_ifinstr_o_19))))

	.dataa(\Mux43~15_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Mux43~13_combout ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux43~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~16 .lut_mask = 16'hCCE2;
defparam \Mux43~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N24
cycloneive_lcell_comb \Mux42~7 (
// Equation(s):
// \Mux42~7_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Reg[27][21]~q )) # (!ifid_ifinstr_o_19 & ((\Reg[19][21]~q )))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[27][21]~q ),
	.datad(\Reg[19][21]~q ),
	.cin(gnd),
	.combout(\Mux42~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~7 .lut_mask = 16'hD9C8;
defparam \Mux42~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N2
cycloneive_lcell_comb \Mux42~8 (
// Equation(s):
// \Mux42~8_combout  = (ifid_ifinstr_o_18 & ((\Mux42~7_combout  & ((\Reg[31][21]~q ))) # (!\Mux42~7_combout  & (\Reg[23][21]~q )))) # (!ifid_ifinstr_o_18 & (((\Mux42~7_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[23][21]~q ),
	.datac(\Reg[31][21]~q ),
	.datad(\Mux42~7_combout ),
	.cin(gnd),
	.combout(\Mux42~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~8 .lut_mask = 16'hF588;
defparam \Mux42~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N12
cycloneive_lcell_comb \Mux42~0 (
// Equation(s):
// \Mux42~0_combout  = (ifid_ifinstr_o_19 & (((\Reg[25][21]~q ) # (ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & (\Reg[17][21]~q  & ((!ifid_ifinstr_o_18))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[17][21]~q ),
	.datac(\Reg[25][21]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux42~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~0 .lut_mask = 16'hAAE4;
defparam \Mux42~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N4
cycloneive_lcell_comb \Mux42~1 (
// Equation(s):
// \Mux42~1_combout  = (ifid_ifinstr_o_18 & ((\Mux42~0_combout  & (\Reg[29][21]~q )) # (!\Mux42~0_combout  & ((\Reg[21][21]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux42~0_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[29][21]~q ),
	.datac(\Reg[21][21]~q ),
	.datad(\Mux42~0_combout ),
	.cin(gnd),
	.combout(\Mux42~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~1 .lut_mask = 16'hDDA0;
defparam \Mux42~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y33_N3
dffeas \Reg[20][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][21] .is_wysiwyg = "true";
defparam \Reg[20][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N2
cycloneive_lcell_comb \Mux42~4 (
// Equation(s):
// \Mux42~4_combout  = (ifid_ifinstr_o_19 & (((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Reg[20][21]~q ))) # (!ifid_ifinstr_o_18 & (\Reg[16][21]~q ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[16][21]~q ),
	.datac(\Reg[20][21]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux42~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~4 .lut_mask = 16'hFA44;
defparam \Mux42~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N17
dffeas \Reg[24][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][21] .is_wysiwyg = "true";
defparam \Reg[24][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N16
cycloneive_lcell_comb \Mux42~5 (
// Equation(s):
// \Mux42~5_combout  = (\Mux42~4_combout  & ((\Reg[28][21]~q ) # ((!ifid_ifinstr_o_19)))) # (!\Mux42~4_combout  & (((\Reg[24][21]~q  & ifid_ifinstr_o_19))))

	.dataa(\Reg[28][21]~q ),
	.datab(\Mux42~4_combout ),
	.datac(\Reg[24][21]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux42~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~5 .lut_mask = 16'hB8CC;
defparam \Mux42~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N23
dffeas \Reg[30][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][21] .is_wysiwyg = "true";
defparam \Reg[30][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N0
cycloneive_lcell_comb \Mux42~2 (
// Equation(s):
// \Mux42~2_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[22][21]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[18][21]~q )))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[22][21]~q ),
	.datad(\Reg[18][21]~q ),
	.cin(gnd),
	.combout(\Mux42~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~2 .lut_mask = 16'hD9C8;
defparam \Mux42~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N22
cycloneive_lcell_comb \Mux42~3 (
// Equation(s):
// \Mux42~3_combout  = (ifid_ifinstr_o_19 & ((\Mux42~2_combout  & ((\Reg[30][21]~q ))) # (!\Mux42~2_combout  & (\Reg[26][21]~q )))) # (!ifid_ifinstr_o_19 & (((\Mux42~2_combout ))))

	.dataa(\Reg[26][21]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[30][21]~q ),
	.datad(\Mux42~2_combout ),
	.cin(gnd),
	.combout(\Mux42~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~3 .lut_mask = 16'hF388;
defparam \Mux42~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N20
cycloneive_lcell_comb \Mux42~6 (
// Equation(s):
// \Mux42~6_combout  = (ifid_ifinstr_o_17 & (((\Mux42~3_combout ) # (ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & (\Mux42~5_combout  & ((!ifid_ifinstr_o_16))))

	.dataa(\Mux42~5_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux42~3_combout ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux42~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~6 .lut_mask = 16'hCCE2;
defparam \Mux42~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y37_N2
cycloneive_lcell_comb \Mux42~17 (
// Equation(s):
// \Mux42~17_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[13][21]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[12][21]~q )))))

	.dataa(\Reg[13][21]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[12][21]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux42~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~17 .lut_mask = 16'hEE30;
defparam \Mux42~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N6
cycloneive_lcell_comb \Mux42~18 (
// Equation(s):
// \Mux42~18_combout  = (ifid_ifinstr_o_17 & ((\Mux42~17_combout  & (\Reg[15][21]~q )) # (!\Mux42~17_combout  & ((\Reg[14][21]~q ))))) # (!ifid_ifinstr_o_17 & (((\Mux42~17_combout ))))

	.dataa(\Reg[15][21]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux42~17_combout ),
	.datad(\Reg[14][21]~q ),
	.cin(gnd),
	.combout(\Mux42~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~18 .lut_mask = 16'hBCB0;
defparam \Mux42~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y39_N29
dffeas \Reg[5][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat27),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][21] .is_wysiwyg = "true";
defparam \Reg[5][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N28
cycloneive_lcell_comb \Mux42~10 (
// Equation(s):
// \Mux42~10_combout  = (ifid_ifinstr_o_16 & (((\Reg[5][21]~q ) # (ifid_ifinstr_o_17)))) # (!ifid_ifinstr_o_16 & (\Reg[4][21]~q  & ((!ifid_ifinstr_o_17))))

	.dataa(\Reg[4][21]~q ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[5][21]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux42~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~10 .lut_mask = 16'hCCE2;
defparam \Mux42~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N28
cycloneive_lcell_comb \Mux42~11 (
// Equation(s):
// \Mux42~11_combout  = (ifid_ifinstr_o_17 & ((\Mux42~10_combout  & ((\Reg[7][21]~q ))) # (!\Mux42~10_combout  & (\Reg[6][21]~q )))) # (!ifid_ifinstr_o_17 & (\Mux42~10_combout ))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux42~10_combout ),
	.datac(\Reg[6][21]~q ),
	.datad(\Reg[7][21]~q ),
	.cin(gnd),
	.combout(\Mux42~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~11 .lut_mask = 16'hEC64;
defparam \Mux42~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N6
cycloneive_lcell_comb \Mux42~15 (
// Equation(s):
// \Mux42~15_combout  = (\Mux42~14_combout ) # ((!ifid_ifinstr_o_16 & (\Reg[2][21]~q  & ifid_ifinstr_o_17)))

	.dataa(\Mux42~14_combout ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[2][21]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux42~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~15 .lut_mask = 16'hBAAA;
defparam \Mux42~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N14
cycloneive_lcell_comb \Mux42~12 (
// Equation(s):
// \Mux42~12_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[10][21]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[8][21]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[8][21]~q ),
	.datad(\Reg[10][21]~q ),
	.cin(gnd),
	.combout(\Mux42~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~12 .lut_mask = 16'hDC98;
defparam \Mux42~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N30
cycloneive_lcell_comb \Mux42~13 (
// Equation(s):
// \Mux42~13_combout  = (ifid_ifinstr_o_16 & ((\Mux42~12_combout  & ((\Reg[11][21]~q ))) # (!\Mux42~12_combout  & (\Reg[9][21]~q )))) # (!ifid_ifinstr_o_16 & (((\Mux42~12_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[9][21]~q ),
	.datac(\Reg[11][21]~q ),
	.datad(\Mux42~12_combout ),
	.cin(gnd),
	.combout(\Mux42~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~13 .lut_mask = 16'hF588;
defparam \Mux42~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N28
cycloneive_lcell_comb \Mux42~16 (
// Equation(s):
// \Mux42~16_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Mux42~13_combout ))) # (!ifid_ifinstr_o_19 & (\Mux42~15_combout ))))

	.dataa(\Mux42~15_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Mux42~13_combout ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux42~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~16 .lut_mask = 16'hFC22;
defparam \Mux42~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N14
cycloneive_lcell_comb \Reg[20][22]~feeder (
// Equation(s):
// \Reg[20][22]~feeder_combout  = \wdat~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat25),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[20][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[20][22]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[20][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N15
dffeas \Reg[20][22] (
	.clk(!CLK),
	.d(\Reg[20][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][22] .is_wysiwyg = "true";
defparam \Reg[20][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N16
cycloneive_lcell_comb \Mux41~4 (
// Equation(s):
// \Mux41~4_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[24][22]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[16][22]~q ))))

	.dataa(\Reg[16][22]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[24][22]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux41~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~4 .lut_mask = 16'hFC22;
defparam \Mux41~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N8
cycloneive_lcell_comb \Mux41~5 (
// Equation(s):
// \Mux41~5_combout  = (ifid_ifinstr_o_18 & ((\Mux41~4_combout  & ((\Reg[28][22]~q ))) # (!\Mux41~4_combout  & (\Reg[20][22]~q )))) # (!ifid_ifinstr_o_18 & (((\Mux41~4_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[20][22]~q ),
	.datac(\Reg[28][22]~q ),
	.datad(\Mux41~4_combout ),
	.cin(gnd),
	.combout(\Mux41~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~5 .lut_mask = 16'hF588;
defparam \Mux41~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N22
cycloneive_lcell_comb \Mux41~2 (
// Equation(s):
// \Mux41~2_combout  = (ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18) # ((\Reg[26][22]~q )))) # (!ifid_ifinstr_o_19 & (!ifid_ifinstr_o_18 & ((\Reg[18][22]~q ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[26][22]~q ),
	.datad(\Reg[18][22]~q ),
	.cin(gnd),
	.combout(\Mux41~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~2 .lut_mask = 16'hB9A8;
defparam \Mux41~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N2
cycloneive_lcell_comb \Mux41~3 (
// Equation(s):
// \Mux41~3_combout  = (ifid_ifinstr_o_18 & ((\Mux41~2_combout  & ((\Reg[30][22]~q ))) # (!\Mux41~2_combout  & (\Reg[22][22]~q )))) # (!ifid_ifinstr_o_18 & (\Mux41~2_combout ))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux41~2_combout ),
	.datac(\Reg[22][22]~q ),
	.datad(\Reg[30][22]~q ),
	.cin(gnd),
	.combout(\Mux41~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~3 .lut_mask = 16'hEC64;
defparam \Mux41~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N12
cycloneive_lcell_comb \Mux41~6 (
// Equation(s):
// \Mux41~6_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Mux41~3_combout ))) # (!ifid_ifinstr_o_17 & (\Mux41~5_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux41~5_combout ),
	.datad(\Mux41~3_combout ),
	.cin(gnd),
	.combout(\Mux41~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~6 .lut_mask = 16'hDC98;
defparam \Mux41~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N14
cycloneive_lcell_comb \Mux41~7 (
// Equation(s):
// \Mux41~7_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Reg[23][22]~q ))) # (!ifid_ifinstr_o_18 & (\Reg[19][22]~q ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[19][22]~q ),
	.datad(\Reg[23][22]~q ),
	.cin(gnd),
	.combout(\Mux41~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~7 .lut_mask = 16'hDC98;
defparam \Mux41~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N10
cycloneive_lcell_comb \Mux41~8 (
// Equation(s):
// \Mux41~8_combout  = (\Mux41~7_combout  & (((\Reg[31][22]~q )) # (!ifid_ifinstr_o_19))) # (!\Mux41~7_combout  & (ifid_ifinstr_o_19 & ((\Reg[27][22]~q ))))

	.dataa(\Mux41~7_combout ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[31][22]~q ),
	.datad(\Reg[27][22]~q ),
	.cin(gnd),
	.combout(\Mux41~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~8 .lut_mask = 16'hE6A2;
defparam \Mux41~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N16
cycloneive_lcell_comb \Mux41~0 (
// Equation(s):
// \Mux41~0_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[21][22]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[17][22]~q )))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[21][22]~q ),
	.datad(\Reg[17][22]~q ),
	.cin(gnd),
	.combout(\Mux41~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~0 .lut_mask = 16'hD9C8;
defparam \Mux41~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y38_N31
dffeas \Reg[25][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat25),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][22] .is_wysiwyg = "true";
defparam \Reg[25][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N30
cycloneive_lcell_comb \Mux41~1 (
// Equation(s):
// \Mux41~1_combout  = (\Mux41~0_combout  & ((\Reg[29][22]~q ) # ((!ifid_ifinstr_o_19)))) # (!\Mux41~0_combout  & (((\Reg[25][22]~q  & ifid_ifinstr_o_19))))

	.dataa(\Reg[29][22]~q ),
	.datab(\Mux41~0_combout ),
	.datac(\Reg[25][22]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux41~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~1 .lut_mask = 16'hB8CC;
defparam \Mux41~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N12
cycloneive_lcell_comb \Mux41~14 (
// Equation(s):
// \Mux41~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[3][22]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[1][22]~q ))))

	.dataa(\Reg[1][22]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[3][22]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux41~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~14 .lut_mask = 16'hE200;
defparam \Mux41~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y35_N20
cycloneive_lcell_comb \Mux41~15 (
// Equation(s):
// \Mux41~15_combout  = (\Mux41~14_combout ) # ((!ifid_ifinstr_o_16 & (ifid_ifinstr_o_17 & \Reg[2][22]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[2][22]~q ),
	.datad(\Mux41~14_combout ),
	.cin(gnd),
	.combout(\Mux41~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~15 .lut_mask = 16'hFF40;
defparam \Mux41~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N14
cycloneive_lcell_comb \Mux41~12 (
// Equation(s):
// \Mux41~12_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[5][22]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[4][22]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[4][22]~q ),
	.datad(\Reg[5][22]~q ),
	.cin(gnd),
	.combout(\Mux41~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~12 .lut_mask = 16'hDC98;
defparam \Mux41~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N30
cycloneive_lcell_comb \Mux41~13 (
// Equation(s):
// \Mux41~13_combout  = (ifid_ifinstr_o_17 & ((\Mux41~12_combout  & ((\Reg[7][22]~q ))) # (!\Mux41~12_combout  & (\Reg[6][22]~q )))) # (!ifid_ifinstr_o_17 & (((\Mux41~12_combout ))))

	.dataa(\Reg[6][22]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[7][22]~q ),
	.datad(\Mux41~12_combout ),
	.cin(gnd),
	.combout(\Mux41~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~13 .lut_mask = 16'hF388;
defparam \Mux41~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N20
cycloneive_lcell_comb \Mux41~16 (
// Equation(s):
// \Mux41~16_combout  = (ifid_ifinstr_o_19 & (((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Mux41~13_combout ))) # (!ifid_ifinstr_o_18 & (\Mux41~15_combout ))))

	.dataa(\Mux41~15_combout ),
	.datab(ifid_ifinstr_o_19),
	.datac(ifid_ifinstr_o_18),
	.datad(\Mux41~13_combout ),
	.cin(gnd),
	.combout(\Mux41~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~16 .lut_mask = 16'hF2C2;
defparam \Mux41~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N30
cycloneive_lcell_comb \Reg[9][22]~feeder (
// Equation(s):
// \Reg[9][22]~feeder_combout  = \wdat~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat25),
	.cin(gnd),
	.combout(\Reg[9][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[9][22]~feeder .lut_mask = 16'hFF00;
defparam \Reg[9][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y32_N31
dffeas \Reg[9][22] (
	.clk(!CLK),
	.d(\Reg[9][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][22] .is_wysiwyg = "true";
defparam \Reg[9][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N4
cycloneive_lcell_comb \Mux41~10 (
// Equation(s):
// \Mux41~10_combout  = (ifid_ifinstr_o_17 & (((\Reg[10][22]~q ) # (ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & (\Reg[8][22]~q  & ((!ifid_ifinstr_o_16))))

	.dataa(\Reg[8][22]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[10][22]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux41~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~10 .lut_mask = 16'hCCE2;
defparam \Mux41~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N18
cycloneive_lcell_comb \Mux41~11 (
// Equation(s):
// \Mux41~11_combout  = (ifid_ifinstr_o_16 & ((\Mux41~10_combout  & ((\Reg[11][22]~q ))) # (!\Mux41~10_combout  & (\Reg[9][22]~q )))) # (!ifid_ifinstr_o_16 & (((\Mux41~10_combout ))))

	.dataa(\Reg[9][22]~q ),
	.datab(\Reg[11][22]~q ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux41~10_combout ),
	.cin(gnd),
	.combout(\Mux41~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~11 .lut_mask = 16'hCFA0;
defparam \Mux41~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y37_N28
cycloneive_lcell_comb \Mux41~17 (
// Equation(s):
// \Mux41~17_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[13][22]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[12][22]~q ))))

	.dataa(\Reg[12][22]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[13][22]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux41~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~17 .lut_mask = 16'hFC22;
defparam \Mux41~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N10
cycloneive_lcell_comb \Mux41~18 (
// Equation(s):
// \Mux41~18_combout  = (ifid_ifinstr_o_17 & ((\Mux41~17_combout  & ((\Reg[15][22]~q ))) # (!\Mux41~17_combout  & (\Reg[14][22]~q )))) # (!ifid_ifinstr_o_17 & (\Mux41~17_combout ))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux41~17_combout ),
	.datac(\Reg[14][22]~q ),
	.datad(\Reg[15][22]~q ),
	.cin(gnd),
	.combout(\Mux41~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~18 .lut_mask = 16'hEC64;
defparam \Mux41~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N14
cycloneive_lcell_comb \Reg[21][23]~feeder (
// Equation(s):
// \Reg[21][23]~feeder_combout  = \wdat~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat26),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[21][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[21][23]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[21][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N15
dffeas \Reg[21][23] (
	.clk(!CLK),
	.d(\Reg[21][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][23] .is_wysiwyg = "true";
defparam \Reg[21][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N16
cycloneive_lcell_comb \Mux40~0 (
// Equation(s):
// \Mux40~0_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Reg[25][23]~q )) # (!ifid_ifinstr_o_19 & ((\Reg[17][23]~q )))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[25][23]~q ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Reg[17][23]~q ),
	.cin(gnd),
	.combout(\Mux40~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~0 .lut_mask = 16'hE5E0;
defparam \Mux40~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N30
cycloneive_lcell_comb \Mux40~1 (
// Equation(s):
// \Mux40~1_combout  = (\Mux40~0_combout  & (((\Reg[29][23]~q ) # (!ifid_ifinstr_o_18)))) # (!\Mux40~0_combout  & (\Reg[21][23]~q  & ((ifid_ifinstr_o_18))))

	.dataa(\Reg[21][23]~q ),
	.datab(\Mux40~0_combout ),
	.datac(\Reg[29][23]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux40~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~1 .lut_mask = 16'hE2CC;
defparam \Mux40~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N26
cycloneive_lcell_comb \Mux40~7 (
// Equation(s):
// \Mux40~7_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[27][23]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[19][23]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[19][23]~q ),
	.datad(\Reg[27][23]~q ),
	.cin(gnd),
	.combout(\Mux40~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~7 .lut_mask = 16'hDC98;
defparam \Mux40~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N22
cycloneive_lcell_comb \Mux40~8 (
// Equation(s):
// \Mux40~8_combout  = (\Mux40~7_combout  & (((\Reg[31][23]~q ) # (!ifid_ifinstr_o_18)))) # (!\Mux40~7_combout  & (\Reg[23][23]~q  & ((ifid_ifinstr_o_18))))

	.dataa(\Mux40~7_combout ),
	.datab(\Reg[23][23]~q ),
	.datac(\Reg[31][23]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux40~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~8 .lut_mask = 16'hE4AA;
defparam \Mux40~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N7
dffeas \Reg[30][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][23] .is_wysiwyg = "true";
defparam \Reg[30][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N6
cycloneive_lcell_comb \Mux40~2 (
// Equation(s):
// \Mux40~2_combout  = (ifid_ifinstr_o_18 & ((\Reg[22][23]~q ) # ((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (((\Reg[18][23]~q  & !ifid_ifinstr_o_19))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[22][23]~q ),
	.datac(\Reg[18][23]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux40~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~2 .lut_mask = 16'hAAD8;
defparam \Mux40~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N6
cycloneive_lcell_comb \Mux40~3 (
// Equation(s):
// \Mux40~3_combout  = (ifid_ifinstr_o_19 & ((\Mux40~2_combout  & ((\Reg[30][23]~q ))) # (!\Mux40~2_combout  & (\Reg[26][23]~q )))) # (!ifid_ifinstr_o_19 & (((\Mux40~2_combout ))))

	.dataa(\Reg[26][23]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[30][23]~q ),
	.datad(\Mux40~2_combout ),
	.cin(gnd),
	.combout(\Mux40~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~3 .lut_mask = 16'hF388;
defparam \Mux40~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N6
cycloneive_lcell_comb \Mux40~5 (
// Equation(s):
// \Mux40~5_combout  = (\Mux40~4_combout  & (((\Reg[28][23]~q ) # (!ifid_ifinstr_o_19)))) # (!\Mux40~4_combout  & (\Reg[24][23]~q  & ((ifid_ifinstr_o_19))))

	.dataa(\Mux40~4_combout ),
	.datab(\Reg[24][23]~q ),
	.datac(\Reg[28][23]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux40~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~5 .lut_mask = 16'hE4AA;
defparam \Mux40~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N22
cycloneive_lcell_comb \Mux40~6 (
// Equation(s):
// \Mux40~6_combout  = (ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16) # ((\Mux40~3_combout )))) # (!ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & ((\Mux40~5_combout ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux40~3_combout ),
	.datad(\Mux40~5_combout ),
	.cin(gnd),
	.combout(\Mux40~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~6 .lut_mask = 16'hB9A8;
defparam \Mux40~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N8
cycloneive_lcell_comb \Mux40~10 (
// Equation(s):
// \Mux40~10_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[5][23]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[4][23]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[5][23]~q ),
	.datad(\Reg[4][23]~q ),
	.cin(gnd),
	.combout(\Mux40~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~10 .lut_mask = 16'hD9C8;
defparam \Mux40~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N0
cycloneive_lcell_comb \Mux40~11 (
// Equation(s):
// \Mux40~11_combout  = (\Mux40~10_combout  & ((\Reg[7][23]~q ) # ((!ifid_ifinstr_o_17)))) # (!\Mux40~10_combout  & (((\Reg[6][23]~q  & ifid_ifinstr_o_17))))

	.dataa(\Reg[7][23]~q ),
	.datab(\Reg[6][23]~q ),
	.datac(\Mux40~10_combout ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux40~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~11 .lut_mask = 16'hACF0;
defparam \Mux40~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N11
dffeas \Reg[2][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[2][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[2][23] .is_wysiwyg = "true";
defparam \Reg[2][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N10
cycloneive_lcell_comb \Mux40~15 (
// Equation(s):
// \Mux40~15_combout  = (\Mux40~14_combout ) # ((!ifid_ifinstr_o_16 & (\Reg[2][23]~q  & ifid_ifinstr_o_17)))

	.dataa(\Mux40~14_combout ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[2][23]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux40~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~15 .lut_mask = 16'hBAAA;
defparam \Mux40~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y32_N23
dffeas \Reg[8][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat26),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][23] .is_wysiwyg = "true";
defparam \Reg[8][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N22
cycloneive_lcell_comb \Mux40~12 (
// Equation(s):
// \Mux40~12_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[10][23]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[8][23]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[8][23]~q ),
	.datad(\Reg[10][23]~q ),
	.cin(gnd),
	.combout(\Mux40~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~12 .lut_mask = 16'hDC98;
defparam \Mux40~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N26
cycloneive_lcell_comb \Mux40~13 (
// Equation(s):
// \Mux40~13_combout  = (ifid_ifinstr_o_16 & ((\Mux40~12_combout  & ((\Reg[11][23]~q ))) # (!\Mux40~12_combout  & (\Reg[9][23]~q )))) # (!ifid_ifinstr_o_16 & (((\Mux40~12_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[9][23]~q ),
	.datac(\Reg[11][23]~q ),
	.datad(\Mux40~12_combout ),
	.cin(gnd),
	.combout(\Mux40~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~13 .lut_mask = 16'hF588;
defparam \Mux40~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N26
cycloneive_lcell_comb \Mux40~16 (
// Equation(s):
// \Mux40~16_combout  = (ifid_ifinstr_o_19 & (((\Mux40~13_combout ) # (ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & (\Mux40~15_combout  & ((!ifid_ifinstr_o_18))))

	.dataa(\Mux40~15_combout ),
	.datab(\Mux40~13_combout ),
	.datac(ifid_ifinstr_o_19),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux40~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~16 .lut_mask = 16'hF0CA;
defparam \Mux40~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y37_N4
cycloneive_lcell_comb \Mux40~17 (
// Equation(s):
// \Mux40~17_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[13][23]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[12][23]~q ))))

	.dataa(\Reg[12][23]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[13][23]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux40~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~17 .lut_mask = 16'hFC22;
defparam \Mux40~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N14
cycloneive_lcell_comb \Mux40~18 (
// Equation(s):
// \Mux40~18_combout  = (ifid_ifinstr_o_17 & ((\Mux40~17_combout  & (\Reg[15][23]~q )) # (!\Mux40~17_combout  & ((\Reg[14][23]~q ))))) # (!ifid_ifinstr_o_17 & (\Mux40~17_combout ))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux40~17_combout ),
	.datac(\Reg[15][23]~q ),
	.datad(\Reg[14][23]~q ),
	.cin(gnd),
	.combout(\Mux40~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~18 .lut_mask = 16'hE6C4;
defparam \Mux40~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N2
cycloneive_lcell_comb \Mux39~7 (
// Equation(s):
// \Mux39~7_combout  = (ifid_ifinstr_o_18 & ((\Reg[23][24]~q ) # ((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (((\Reg[19][24]~q  & !ifid_ifinstr_o_19))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[23][24]~q ),
	.datac(\Reg[19][24]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux39~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~7 .lut_mask = 16'hAAD8;
defparam \Mux39~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N10
cycloneive_lcell_comb \Mux39~8 (
// Equation(s):
// \Mux39~8_combout  = (ifid_ifinstr_o_19 & ((\Mux39~7_combout  & ((\Reg[31][24]~q ))) # (!\Mux39~7_combout  & (\Reg[27][24]~q )))) # (!ifid_ifinstr_o_19 & (((\Mux39~7_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[27][24]~q ),
	.datac(\Reg[31][24]~q ),
	.datad(\Mux39~7_combout ),
	.cin(gnd),
	.combout(\Mux39~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~8 .lut_mask = 16'hF588;
defparam \Mux39~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N30
cycloneive_lcell_comb \Mux39~4 (
// Equation(s):
// \Mux39~4_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Reg[24][24]~q )) # (!ifid_ifinstr_o_19 & ((\Reg[16][24]~q )))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[24][24]~q ),
	.datac(\Reg[16][24]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux39~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~4 .lut_mask = 16'hEE50;
defparam \Mux39~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N9
dffeas \Reg[28][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][24] .is_wysiwyg = "true";
defparam \Reg[28][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N30
cycloneive_lcell_comb \Reg[20][24]~feeder (
// Equation(s):
// \Reg[20][24]~feeder_combout  = \wdat~51_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat24),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[20][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[20][24]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[20][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y34_N31
dffeas \Reg[20][24] (
	.clk(!CLK),
	.d(\Reg[20][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][24] .is_wysiwyg = "true";
defparam \Reg[20][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N8
cycloneive_lcell_comb \Mux39~5 (
// Equation(s):
// \Mux39~5_combout  = (ifid_ifinstr_o_18 & ((\Mux39~4_combout  & (\Reg[28][24]~q )) # (!\Mux39~4_combout  & ((\Reg[20][24]~q ))))) # (!ifid_ifinstr_o_18 & (\Mux39~4_combout ))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux39~4_combout ),
	.datac(\Reg[28][24]~q ),
	.datad(\Reg[20][24]~q ),
	.cin(gnd),
	.combout(\Mux39~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~5 .lut_mask = 16'hE6C4;
defparam \Mux39~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N4
cycloneive_lcell_comb \Mux39~2 (
// Equation(s):
// \Mux39~2_combout  = (ifid_ifinstr_o_19 & (((\Reg[26][24]~q ) # (ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & (\Reg[18][24]~q  & ((!ifid_ifinstr_o_18))))

	.dataa(\Reg[18][24]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[26][24]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux39~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~2 .lut_mask = 16'hCCE2;
defparam \Mux39~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N10
cycloneive_lcell_comb \Mux39~3 (
// Equation(s):
// \Mux39~3_combout  = (ifid_ifinstr_o_18 & ((\Mux39~2_combout  & (\Reg[30][24]~q )) # (!\Mux39~2_combout  & ((\Reg[22][24]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux39~2_combout ))))

	.dataa(\Reg[30][24]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[22][24]~q ),
	.datad(\Mux39~2_combout ),
	.cin(gnd),
	.combout(\Mux39~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~3 .lut_mask = 16'hBBC0;
defparam \Mux39~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N24
cycloneive_lcell_comb \Mux39~6 (
// Equation(s):
// \Mux39~6_combout  = (ifid_ifinstr_o_17 & (((\Mux39~3_combout ) # (ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & (\Mux39~5_combout  & ((!ifid_ifinstr_o_16))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux39~5_combout ),
	.datac(\Mux39~3_combout ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux39~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~6 .lut_mask = 16'hAAE4;
defparam \Mux39~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N14
cycloneive_lcell_comb \Mux39~0 (
// Equation(s):
// \Mux39~0_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[21][24]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[17][24]~q )))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[21][24]~q ),
	.datad(\Reg[17][24]~q ),
	.cin(gnd),
	.combout(\Mux39~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~0 .lut_mask = 16'hD9C8;
defparam \Mux39~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N6
cycloneive_lcell_comb \Mux39~1 (
// Equation(s):
// \Mux39~1_combout  = (\Mux39~0_combout  & ((\Reg[29][24]~q ) # ((!ifid_ifinstr_o_19)))) # (!\Mux39~0_combout  & (((\Reg[25][24]~q  & ifid_ifinstr_o_19))))

	.dataa(\Mux39~0_combout ),
	.datab(\Reg[29][24]~q ),
	.datac(\Reg[25][24]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux39~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~1 .lut_mask = 16'hD8AA;
defparam \Mux39~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y37_N20
cycloneive_lcell_comb \Mux39~17 (
// Equation(s):
// \Mux39~17_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17) # ((\Reg[13][24]~q )))) # (!ifid_ifinstr_o_16 & (!ifid_ifinstr_o_17 & ((\Reg[12][24]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[13][24]~q ),
	.datad(\Reg[12][24]~q ),
	.cin(gnd),
	.combout(\Mux39~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~17 .lut_mask = 16'hB9A8;
defparam \Mux39~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N30
cycloneive_lcell_comb \Mux39~18 (
// Equation(s):
// \Mux39~18_combout  = (\Mux39~17_combout  & ((\Reg[15][24]~q ) # ((!ifid_ifinstr_o_17)))) # (!\Mux39~17_combout  & (((\Reg[14][24]~q  & ifid_ifinstr_o_17))))

	.dataa(\Mux39~17_combout ),
	.datab(\Reg[15][24]~q ),
	.datac(\Reg[14][24]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux39~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~18 .lut_mask = 16'hD8AA;
defparam \Mux39~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N26
cycloneive_lcell_comb \Mux39~15 (
// Equation(s):
// \Mux39~15_combout  = (\Mux39~14_combout ) # ((ifid_ifinstr_o_17 & (\Reg[2][24]~q  & !ifid_ifinstr_o_16)))

	.dataa(\Mux39~14_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[2][24]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux39~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~15 .lut_mask = 16'hAAEA;
defparam \Mux39~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y39_N31
dffeas \Reg[4][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][24] .is_wysiwyg = "true";
defparam \Reg[4][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N30
cycloneive_lcell_comb \Mux39~12 (
// Equation(s):
// \Mux39~12_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[5][24]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[4][24]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[4][24]~q ),
	.datad(\Reg[5][24]~q ),
	.cin(gnd),
	.combout(\Mux39~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~12 .lut_mask = 16'hDC98;
defparam \Mux39~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N20
cycloneive_lcell_comb \Mux39~13 (
// Equation(s):
// \Mux39~13_combout  = (ifid_ifinstr_o_17 & ((\Mux39~12_combout  & ((\Reg[7][24]~q ))) # (!\Mux39~12_combout  & (\Reg[6][24]~q )))) # (!ifid_ifinstr_o_17 & (((\Mux39~12_combout ))))

	.dataa(\Reg[6][24]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[7][24]~q ),
	.datad(\Mux39~12_combout ),
	.cin(gnd),
	.combout(\Mux39~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~13 .lut_mask = 16'hF388;
defparam \Mux39~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N28
cycloneive_lcell_comb \Mux39~16 (
// Equation(s):
// \Mux39~16_combout  = (ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19) # ((\Mux39~13_combout )))) # (!ifid_ifinstr_o_18 & (!ifid_ifinstr_o_19 & (\Mux39~15_combout )))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Mux39~15_combout ),
	.datad(\Mux39~13_combout ),
	.cin(gnd),
	.combout(\Mux39~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~16 .lut_mask = 16'hBA98;
defparam \Mux39~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N28
cycloneive_lcell_comb \Mux39~10 (
// Equation(s):
// \Mux39~10_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[10][24]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[8][24]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[10][24]~q ),
	.datad(\Reg[8][24]~q ),
	.cin(gnd),
	.combout(\Mux39~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~10 .lut_mask = 16'hD9C8;
defparam \Mux39~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N13
dffeas \Reg[9][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat24),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][24] .is_wysiwyg = "true";
defparam \Reg[9][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N12
cycloneive_lcell_comb \Mux39~11 (
// Equation(s):
// \Mux39~11_combout  = (\Mux39~10_combout  & ((\Reg[11][24]~q ) # ((!ifid_ifinstr_o_16)))) # (!\Mux39~10_combout  & (((\Reg[9][24]~q  & ifid_ifinstr_o_16))))

	.dataa(\Mux39~10_combout ),
	.datab(\Reg[11][24]~q ),
	.datac(\Reg[9][24]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux39~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~11 .lut_mask = 16'hD8AA;
defparam \Mux39~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N6
cycloneive_lcell_comb \Mux38~7 (
// Equation(s):
// \Mux38~7_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Reg[27][25]~q )) # (!ifid_ifinstr_o_19 & ((\Reg[19][25]~q )))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[27][25]~q ),
	.datac(\Reg[19][25]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux38~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~7 .lut_mask = 16'hEE50;
defparam \Mux38~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N0
cycloneive_lcell_comb \Mux38~8 (
// Equation(s):
// \Mux38~8_combout  = (ifid_ifinstr_o_18 & ((\Mux38~7_combout  & (\Reg[31][25]~q )) # (!\Mux38~7_combout  & ((\Reg[23][25]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux38~7_combout ))))

	.dataa(\Reg[31][25]~q ),
	.datab(\Reg[23][25]~q ),
	.datac(ifid_ifinstr_o_18),
	.datad(\Mux38~7_combout ),
	.cin(gnd),
	.combout(\Mux38~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~8 .lut_mask = 16'hAFC0;
defparam \Mux38~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y33_N31
dffeas \Reg[16][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][25] .is_wysiwyg = "true";
defparam \Reg[16][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N30
cycloneive_lcell_comb \Mux38~4 (
// Equation(s):
// \Mux38~4_combout  = (ifid_ifinstr_o_19 & (((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[20][25]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[16][25]~q )))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[20][25]~q ),
	.datac(\Reg[16][25]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux38~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~4 .lut_mask = 16'hEE50;
defparam \Mux38~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N4
cycloneive_lcell_comb \Mux38~5 (
// Equation(s):
// \Mux38~5_combout  = (ifid_ifinstr_o_19 & ((\Mux38~4_combout  & ((\Reg[28][25]~q ))) # (!\Mux38~4_combout  & (\Reg[24][25]~q )))) # (!ifid_ifinstr_o_19 & (((\Mux38~4_combout ))))

	.dataa(\Reg[24][25]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[28][25]~q ),
	.datad(\Mux38~4_combout ),
	.cin(gnd),
	.combout(\Mux38~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~5 .lut_mask = 16'hF388;
defparam \Mux38~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N4
cycloneive_lcell_comb \Mux38~2 (
// Equation(s):
// \Mux38~2_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[22][25]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[18][25]~q )))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[22][25]~q ),
	.datad(\Reg[18][25]~q ),
	.cin(gnd),
	.combout(\Mux38~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~2 .lut_mask = 16'hD9C8;
defparam \Mux38~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N18
cycloneive_lcell_comb \Mux38~3 (
// Equation(s):
// \Mux38~3_combout  = (ifid_ifinstr_o_19 & ((\Mux38~2_combout  & (\Reg[30][25]~q )) # (!\Mux38~2_combout  & ((\Reg[26][25]~q ))))) # (!ifid_ifinstr_o_19 & (\Mux38~2_combout ))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Mux38~2_combout ),
	.datac(\Reg[30][25]~q ),
	.datad(\Reg[26][25]~q ),
	.cin(gnd),
	.combout(\Mux38~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~3 .lut_mask = 16'hE6C4;
defparam \Mux38~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N26
cycloneive_lcell_comb \Mux38~6 (
// Equation(s):
// \Mux38~6_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16) # (\Mux38~3_combout )))) # (!ifid_ifinstr_o_17 & (\Mux38~5_combout  & (!ifid_ifinstr_o_16)))

	.dataa(\Mux38~5_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux38~3_combout ),
	.cin(gnd),
	.combout(\Mux38~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~6 .lut_mask = 16'hCEC2;
defparam \Mux38~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N8
cycloneive_lcell_comb \Mux38~0 (
// Equation(s):
// \Mux38~0_combout  = (ifid_ifinstr_o_19 & (((\Reg[25][25]~q ) # (ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & (\Reg[17][25]~q  & ((!ifid_ifinstr_o_18))))

	.dataa(\Reg[17][25]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[25][25]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux38~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~0 .lut_mask = 16'hCCE2;
defparam \Mux38~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N12
cycloneive_lcell_comb \Mux38~1 (
// Equation(s):
// \Mux38~1_combout  = (ifid_ifinstr_o_18 & ((\Mux38~0_combout  & (\Reg[29][25]~q )) # (!\Mux38~0_combout  & ((\Reg[21][25]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux38~0_combout ))))

	.dataa(\Reg[29][25]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[21][25]~q ),
	.datad(\Mux38~0_combout ),
	.cin(gnd),
	.combout(\Mux38~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~1 .lut_mask = 16'hBBC0;
defparam \Mux38~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y37_N12
cycloneive_lcell_comb \Mux38~17 (
// Equation(s):
// \Mux38~17_combout  = (ifid_ifinstr_o_16 & (((\Reg[13][25]~q ) # (ifid_ifinstr_o_17)))) # (!ifid_ifinstr_o_16 & (\Reg[12][25]~q  & ((!ifid_ifinstr_o_17))))

	.dataa(\Reg[12][25]~q ),
	.datab(\Reg[13][25]~q ),
	.datac(ifid_ifinstr_o_16),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux38~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~17 .lut_mask = 16'hF0CA;
defparam \Mux38~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N24
cycloneive_lcell_comb \Mux38~18 (
// Equation(s):
// \Mux38~18_combout  = (ifid_ifinstr_o_17 & ((\Mux38~17_combout  & (\Reg[15][25]~q )) # (!\Mux38~17_combout  & ((\Reg[14][25]~q ))))) # (!ifid_ifinstr_o_17 & (((\Mux38~17_combout ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[15][25]~q ),
	.datac(\Reg[14][25]~q ),
	.datad(\Mux38~17_combout ),
	.cin(gnd),
	.combout(\Mux38~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~18 .lut_mask = 16'hDDA0;
defparam \Mux38~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N31
dffeas \Reg[6][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][25] .is_wysiwyg = "true";
defparam \Reg[6][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y39_N4
cycloneive_lcell_comb \Mux38~10 (
// Equation(s):
// \Mux38~10_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[5][25]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[4][25]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[5][25]~q ),
	.datad(\Reg[4][25]~q ),
	.cin(gnd),
	.combout(\Mux38~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~10 .lut_mask = 16'hD9C8;
defparam \Mux38~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N30
cycloneive_lcell_comb \Mux38~11 (
// Equation(s):
// \Mux38~11_combout  = (ifid_ifinstr_o_17 & ((\Mux38~10_combout  & (\Reg[7][25]~q )) # (!\Mux38~10_combout  & ((\Reg[6][25]~q ))))) # (!ifid_ifinstr_o_17 & (((\Mux38~10_combout ))))

	.dataa(\Reg[7][25]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[6][25]~q ),
	.datad(\Mux38~10_combout ),
	.cin(gnd),
	.combout(\Mux38~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~11 .lut_mask = 16'hBBC0;
defparam \Mux38~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y32_N27
dffeas \Reg[8][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat23),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][25] .is_wysiwyg = "true";
defparam \Reg[8][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N26
cycloneive_lcell_comb \Mux38~12 (
// Equation(s):
// \Mux38~12_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[10][25]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[8][25]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[8][25]~q ),
	.datad(\Reg[10][25]~q ),
	.cin(gnd),
	.combout(\Mux38~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~12 .lut_mask = 16'hDC98;
defparam \Mux38~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N6
cycloneive_lcell_comb \Mux38~13 (
// Equation(s):
// \Mux38~13_combout  = (ifid_ifinstr_o_16 & ((\Mux38~12_combout  & (\Reg[11][25]~q )) # (!\Mux38~12_combout  & ((\Reg[9][25]~q ))))) # (!ifid_ifinstr_o_16 & (\Mux38~12_combout ))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux38~12_combout ),
	.datac(\Reg[11][25]~q ),
	.datad(\Reg[9][25]~q ),
	.cin(gnd),
	.combout(\Mux38~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~13 .lut_mask = 16'hE6C4;
defparam \Mux38~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N28
cycloneive_lcell_comb \Mux38~14 (
// Equation(s):
// \Mux38~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[3][25]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[1][25]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[1][25]~q ),
	.datad(\Reg[3][25]~q ),
	.cin(gnd),
	.combout(\Mux38~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~14 .lut_mask = 16'hA820;
defparam \Mux38~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N20
cycloneive_lcell_comb \Mux38~15 (
// Equation(s):
// \Mux38~15_combout  = (\Mux38~14_combout ) # ((!ifid_ifinstr_o_16 & (ifid_ifinstr_o_17 & \Reg[2][25]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[2][25]~q ),
	.datad(\Mux38~14_combout ),
	.cin(gnd),
	.combout(\Mux38~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~15 .lut_mask = 16'hFF40;
defparam \Mux38~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N2
cycloneive_lcell_comb \Mux38~16 (
// Equation(s):
// \Mux38~16_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Mux38~13_combout )) # (!ifid_ifinstr_o_19 & ((\Mux38~15_combout )))))

	.dataa(\Mux38~13_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux38~15_combout ),
	.cin(gnd),
	.combout(\Mux38~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~16 .lut_mask = 16'hE3E0;
defparam \Mux38~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N10
cycloneive_lcell_comb \Mux37~0 (
// Equation(s):
// \Mux37~0_combout  = (ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19) # ((\Reg[21][26]~q )))) # (!ifid_ifinstr_o_18 & (!ifid_ifinstr_o_19 & (\Reg[17][26]~q )))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[17][26]~q ),
	.datad(\Reg[21][26]~q ),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~0 .lut_mask = 16'hBA98;
defparam \Mux37~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N28
cycloneive_lcell_comb \Mux37~1 (
// Equation(s):
// \Mux37~1_combout  = (\Mux37~0_combout  & (((\Reg[29][26]~q ) # (!ifid_ifinstr_o_19)))) # (!\Mux37~0_combout  & (\Reg[25][26]~q  & ((ifid_ifinstr_o_19))))

	.dataa(\Mux37~0_combout ),
	.datab(\Reg[25][26]~q ),
	.datac(\Reg[29][26]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux37~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~1 .lut_mask = 16'hE4AA;
defparam \Mux37~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N30
cycloneive_lcell_comb \Reg[27][26]~feeder (
// Equation(s):
// \Reg[27][26]~feeder_combout  = \wdat~45_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat21),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[27][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[27][26]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[27][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N31
dffeas \Reg[27][26] (
	.clk(!CLK),
	.d(\Reg[27][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][26] .is_wysiwyg = "true";
defparam \Reg[27][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N4
cycloneive_lcell_comb \Mux37~7 (
// Equation(s):
// \Mux37~7_combout  = (ifid_ifinstr_o_18 & (((\Reg[23][26]~q ) # (ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (\Reg[19][26]~q  & ((!ifid_ifinstr_o_19))))

	.dataa(\Reg[19][26]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[23][26]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux37~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~7 .lut_mask = 16'hCCE2;
defparam \Mux37~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N30
cycloneive_lcell_comb \Mux37~8 (
// Equation(s):
// \Mux37~8_combout  = (ifid_ifinstr_o_19 & ((\Mux37~7_combout  & ((\Reg[31][26]~q ))) # (!\Mux37~7_combout  & (\Reg[27][26]~q )))) # (!ifid_ifinstr_o_19 & (((\Mux37~7_combout ))))

	.dataa(\Reg[27][26]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[31][26]~q ),
	.datad(\Mux37~7_combout ),
	.cin(gnd),
	.combout(\Mux37~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~8 .lut_mask = 16'hF388;
defparam \Mux37~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N0
cycloneive_lcell_comb \Mux37~4 (
// Equation(s):
// \Mux37~4_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Reg[24][26]~q )) # (!ifid_ifinstr_o_19 & ((\Reg[16][26]~q )))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[24][26]~q ),
	.datad(\Reg[16][26]~q ),
	.cin(gnd),
	.combout(\Mux37~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~4 .lut_mask = 16'hD9C8;
defparam \Mux37~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N4
cycloneive_lcell_comb \Mux37~5 (
// Equation(s):
// \Mux37~5_combout  = (ifid_ifinstr_o_18 & ((\Mux37~4_combout  & (\Reg[28][26]~q )) # (!\Mux37~4_combout  & ((\Reg[20][26]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux37~4_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[28][26]~q ),
	.datac(\Reg[20][26]~q ),
	.datad(\Mux37~4_combout ),
	.cin(gnd),
	.combout(\Mux37~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~5 .lut_mask = 16'hDDA0;
defparam \Mux37~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N14
cycloneive_lcell_comb \Mux37~2 (
// Equation(s):
// \Mux37~2_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Reg[26][26]~q )) # (!ifid_ifinstr_o_19 & ((\Reg[18][26]~q )))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[26][26]~q ),
	.datad(\Reg[18][26]~q ),
	.cin(gnd),
	.combout(\Mux37~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~2 .lut_mask = 16'hD9C8;
defparam \Mux37~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N20
cycloneive_lcell_comb \Mux37~3 (
// Equation(s):
// \Mux37~3_combout  = (\Mux37~2_combout  & ((\Reg[30][26]~q ) # ((!ifid_ifinstr_o_18)))) # (!\Mux37~2_combout  & (((\Reg[22][26]~q  & ifid_ifinstr_o_18))))

	.dataa(\Reg[30][26]~q ),
	.datab(\Mux37~2_combout ),
	.datac(\Reg[22][26]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux37~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~3 .lut_mask = 16'hB8CC;
defparam \Mux37~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N22
cycloneive_lcell_comb \Mux37~6 (
// Equation(s):
// \Mux37~6_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16) # (\Mux37~3_combout )))) # (!ifid_ifinstr_o_17 & (\Mux37~5_combout  & (!ifid_ifinstr_o_16)))

	.dataa(\Mux37~5_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux37~3_combout ),
	.cin(gnd),
	.combout(\Mux37~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~6 .lut_mask = 16'hCEC2;
defparam \Mux37~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N18
cycloneive_lcell_comb \Mux37~14 (
// Equation(s):
// \Mux37~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[3][26]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[1][26]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[1][26]~q ),
	.datad(\Reg[3][26]~q ),
	.cin(gnd),
	.combout(\Mux37~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~14 .lut_mask = 16'hA820;
defparam \Mux37~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N16
cycloneive_lcell_comb \Mux37~15 (
// Equation(s):
// \Mux37~15_combout  = (\Mux37~14_combout ) # ((!ifid_ifinstr_o_16 & (\Reg[2][26]~q  & ifid_ifinstr_o_17)))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux37~14_combout ),
	.datac(\Reg[2][26]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux37~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~15 .lut_mask = 16'hDCCC;
defparam \Mux37~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N14
cycloneive_lcell_comb \Mux37~13 (
// Equation(s):
// \Mux37~13_combout  = (\Mux37~12_combout  & (((\Reg[7][26]~q )) # (!ifid_ifinstr_o_17))) # (!\Mux37~12_combout  & (ifid_ifinstr_o_17 & ((\Reg[6][26]~q ))))

	.dataa(\Mux37~12_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[7][26]~q ),
	.datad(\Reg[6][26]~q ),
	.cin(gnd),
	.combout(\Mux37~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~13 .lut_mask = 16'hE6A2;
defparam \Mux37~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N26
cycloneive_lcell_comb \Mux37~16 (
// Equation(s):
// \Mux37~16_combout  = (ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19) # ((\Mux37~13_combout )))) # (!ifid_ifinstr_o_18 & (!ifid_ifinstr_o_19 & (\Mux37~15_combout )))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Mux37~15_combout ),
	.datad(\Mux37~13_combout ),
	.cin(gnd),
	.combout(\Mux37~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~16 .lut_mask = 16'hBA98;
defparam \Mux37~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N12
cycloneive_lcell_comb \Mux37~10 (
// Equation(s):
// \Mux37~10_combout  = (ifid_ifinstr_o_17 & (((\Reg[10][26]~q ) # (ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & (\Reg[8][26]~q  & ((!ifid_ifinstr_o_16))))

	.dataa(\Reg[8][26]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[10][26]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux37~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~10 .lut_mask = 16'hCCE2;
defparam \Mux37~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N8
cycloneive_lcell_comb \Mux37~11 (
// Equation(s):
// \Mux37~11_combout  = (ifid_ifinstr_o_16 & ((\Mux37~10_combout  & (\Reg[11][26]~q )) # (!\Mux37~10_combout  & ((\Reg[9][26]~q ))))) # (!ifid_ifinstr_o_16 & (((\Mux37~10_combout ))))

	.dataa(\Reg[11][26]~q ),
	.datab(\Reg[9][26]~q ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux37~10_combout ),
	.cin(gnd),
	.combout(\Mux37~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~11 .lut_mask = 16'hAFC0;
defparam \Mux37~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y37_N10
cycloneive_lcell_comb \Mux37~17 (
// Equation(s):
// \Mux37~17_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17) # ((\Reg[13][26]~q )))) # (!ifid_ifinstr_o_16 & (!ifid_ifinstr_o_17 & (\Reg[12][26]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[12][26]~q ),
	.datad(\Reg[13][26]~q ),
	.cin(gnd),
	.combout(\Mux37~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~17 .lut_mask = 16'hBA98;
defparam \Mux37~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N24
cycloneive_lcell_comb \Mux37~18 (
// Equation(s):
// \Mux37~18_combout  = (\Mux37~17_combout  & ((\Reg[15][26]~q ) # ((!ifid_ifinstr_o_17)))) # (!\Mux37~17_combout  & (((\Reg[14][26]~q  & ifid_ifinstr_o_17))))

	.dataa(\Mux37~17_combout ),
	.datab(\Reg[15][26]~q ),
	.datac(\Reg[14][26]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux37~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~18 .lut_mask = 16'hD8AA;
defparam \Mux37~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N15
dffeas \Reg[19][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][5] .is_wysiwyg = "true";
defparam \Reg[19][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N14
cycloneive_lcell_comb \Mux58~7 (
// Equation(s):
// \Mux58~7_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Reg[27][5]~q )) # (!ifid_ifinstr_o_19 & ((\Reg[19][5]~q )))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[27][5]~q ),
	.datac(\Reg[19][5]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux58~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~7 .lut_mask = 16'hEE50;
defparam \Mux58~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N24
cycloneive_lcell_comb \Mux58~8 (
// Equation(s):
// \Mux58~8_combout  = (ifid_ifinstr_o_18 & ((\Mux58~7_combout  & ((\Reg[31][5]~q ))) # (!\Mux58~7_combout  & (\Reg[23][5]~q )))) # (!ifid_ifinstr_o_18 & (((\Mux58~7_combout ))))

	.dataa(\Reg[23][5]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Mux58~7_combout ),
	.datad(\Reg[31][5]~q ),
	.cin(gnd),
	.combout(\Mux58~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~8 .lut_mask = 16'hF838;
defparam \Mux58~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N0
cycloneive_lcell_comb \Mux58~0 (
// Equation(s):
// \Mux58~0_combout  = (ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18) # ((\Reg[25][5]~q )))) # (!ifid_ifinstr_o_19 & (!ifid_ifinstr_o_18 & (\Reg[17][5]~q )))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[17][5]~q ),
	.datad(\Reg[25][5]~q ),
	.cin(gnd),
	.combout(\Mux58~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~0 .lut_mask = 16'hBA98;
defparam \Mux58~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N6
cycloneive_lcell_comb \Mux58~1 (
// Equation(s):
// \Mux58~1_combout  = (\Mux58~0_combout  & (((\Reg[29][5]~q ) # (!ifid_ifinstr_o_18)))) # (!\Mux58~0_combout  & (\Reg[21][5]~q  & ((ifid_ifinstr_o_18))))

	.dataa(\Reg[21][5]~q ),
	.datab(\Mux58~0_combout ),
	.datac(\Reg[29][5]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux58~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~1 .lut_mask = 16'hE2CC;
defparam \Mux58~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N10
cycloneive_lcell_comb \Mux58~3 (
// Equation(s):
// \Mux58~3_combout  = (\Mux58~2_combout  & ((\Reg[30][5]~q ) # ((!ifid_ifinstr_o_19)))) # (!\Mux58~2_combout  & (((\Reg[26][5]~q  & ifid_ifinstr_o_19))))

	.dataa(\Mux58~2_combout ),
	.datab(\Reg[30][5]~q ),
	.datac(\Reg[26][5]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux58~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~3 .lut_mask = 16'hD8AA;
defparam \Mux58~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N18
cycloneive_lcell_comb \Mux58~4 (
// Equation(s):
// \Mux58~4_combout  = (ifid_ifinstr_o_19 & (((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Reg[20][5]~q ))) # (!ifid_ifinstr_o_18 & (\Reg[16][5]~q ))))

	.dataa(\Reg[16][5]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[20][5]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux58~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~4 .lut_mask = 16'hFC22;
defparam \Mux58~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N12
cycloneive_lcell_comb \Mux58~5 (
// Equation(s):
// \Mux58~5_combout  = (\Mux58~4_combout  & ((\Reg[28][5]~q ) # ((!ifid_ifinstr_o_19)))) # (!\Mux58~4_combout  & (((\Reg[24][5]~q  & ifid_ifinstr_o_19))))

	.dataa(\Reg[28][5]~q ),
	.datab(\Mux58~4_combout ),
	.datac(\Reg[24][5]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux58~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~5 .lut_mask = 16'hB8CC;
defparam \Mux58~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N18
cycloneive_lcell_comb \Mux58~6 (
// Equation(s):
// \Mux58~6_combout  = (ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16) # ((\Mux58~3_combout )))) # (!ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & ((\Mux58~5_combout ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux58~3_combout ),
	.datad(\Mux58~5_combout ),
	.cin(gnd),
	.combout(\Mux58~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~6 .lut_mask = 16'hB9A8;
defparam \Mux58~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N20
cycloneive_lcell_comb \Mux58~10 (
// Equation(s):
// \Mux58~10_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[5][5]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[4][5]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[4][5]~q ),
	.datac(\Reg[5][5]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux58~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~10 .lut_mask = 16'hFA44;
defparam \Mux58~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N13
dffeas \Reg[6][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[6][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[6][5] .is_wysiwyg = "true";
defparam \Reg[6][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N4
cycloneive_lcell_comb \Mux58~11 (
// Equation(s):
// \Mux58~11_combout  = (ifid_ifinstr_o_17 & ((\Mux58~10_combout  & (\Reg[7][5]~q )) # (!\Mux58~10_combout  & ((\Reg[6][5]~q ))))) # (!ifid_ifinstr_o_17 & (((\Mux58~10_combout ))))

	.dataa(\Reg[7][5]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux58~10_combout ),
	.datad(\Reg[6][5]~q ),
	.cin(gnd),
	.combout(\Mux58~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~11 .lut_mask = 16'hBCB0;
defparam \Mux58~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y34_N31
dffeas \Reg[12][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][5] .is_wysiwyg = "true";
defparam \Reg[12][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N30
cycloneive_lcell_comb \Mux58~17 (
// Equation(s):
// \Mux58~17_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17) # ((\Reg[13][5]~q )))) # (!ifid_ifinstr_o_16 & (!ifid_ifinstr_o_17 & (\Reg[12][5]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[12][5]~q ),
	.datad(\Reg[13][5]~q ),
	.cin(gnd),
	.combout(\Mux58~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~17 .lut_mask = 16'hBA98;
defparam \Mux58~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N26
cycloneive_lcell_comb \Mux58~18 (
// Equation(s):
// \Mux58~18_combout  = (\Mux58~17_combout  & (((\Reg[15][5]~q )) # (!ifid_ifinstr_o_17))) # (!\Mux58~17_combout  & (ifid_ifinstr_o_17 & ((\Reg[14][5]~q ))))

	.dataa(\Mux58~17_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[15][5]~q ),
	.datad(\Reg[14][5]~q ),
	.cin(gnd),
	.combout(\Mux58~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~18 .lut_mask = 16'hE6A2;
defparam \Mux58~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y35_N6
cycloneive_lcell_comb \Mux58~14 (
// Equation(s):
// \Mux58~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[3][5]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[1][5]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[1][5]~q ),
	.datad(\Reg[3][5]~q ),
	.cin(gnd),
	.combout(\Mux58~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~14 .lut_mask = 16'hA820;
defparam \Mux58~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N14
cycloneive_lcell_comb \Mux58~15 (
// Equation(s):
// \Mux58~15_combout  = (\Mux58~14_combout ) # ((!ifid_ifinstr_o_16 & (ifid_ifinstr_o_17 & \Reg[2][5]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[2][5]~q ),
	.datad(\Mux58~14_combout ),
	.cin(gnd),
	.combout(\Mux58~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~15 .lut_mask = 16'hFF40;
defparam \Mux58~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y31_N11
dffeas \Reg[8][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat8),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][5] .is_wysiwyg = "true";
defparam \Reg[8][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N10
cycloneive_lcell_comb \Mux58~12 (
// Equation(s):
// \Mux58~12_combout  = (ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16) # ((\Reg[10][5]~q )))) # (!ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & (\Reg[8][5]~q )))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[8][5]~q ),
	.datad(\Reg[10][5]~q ),
	.cin(gnd),
	.combout(\Mux58~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~12 .lut_mask = 16'hBA98;
defparam \Mux58~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N26
cycloneive_lcell_comb \Mux58~13 (
// Equation(s):
// \Mux58~13_combout  = (ifid_ifinstr_o_16 & ((\Mux58~12_combout  & ((\Reg[11][5]~q ))) # (!\Mux58~12_combout  & (\Reg[9][5]~q )))) # (!ifid_ifinstr_o_16 & (((\Mux58~12_combout ))))

	.dataa(\Reg[9][5]~q ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[11][5]~q ),
	.datad(\Mux58~12_combout ),
	.cin(gnd),
	.combout(\Mux58~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~13 .lut_mask = 16'hF388;
defparam \Mux58~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N0
cycloneive_lcell_comb \Mux58~16 (
// Equation(s):
// \Mux58~16_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Mux58~13_combout ))) # (!ifid_ifinstr_o_19 & (\Mux58~15_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux58~15_combout ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux58~13_combout ),
	.cin(gnd),
	.combout(\Mux58~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~16 .lut_mask = 16'hF4A4;
defparam \Mux58~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N2
cycloneive_lcell_comb \Mux57~7 (
// Equation(s):
// \Mux57~7_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[23][6]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[19][6]~q )))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[23][6]~q ),
	.datad(\Reg[19][6]~q ),
	.cin(gnd),
	.combout(\Mux57~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~7 .lut_mask = 16'hD9C8;
defparam \Mux57~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N8
cycloneive_lcell_comb \Mux57~8 (
// Equation(s):
// \Mux57~8_combout  = (ifid_ifinstr_o_19 & ((\Mux57~7_combout  & (\Reg[31][6]~q )) # (!\Mux57~7_combout  & ((\Reg[27][6]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux57~7_combout ))))

	.dataa(\Reg[31][6]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[27][6]~q ),
	.datad(\Mux57~7_combout ),
	.cin(gnd),
	.combout(\Mux57~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~8 .lut_mask = 16'hBBC0;
defparam \Mux57~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y38_N31
dffeas \Reg[17][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~3_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[17][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[17][6] .is_wysiwyg = "true";
defparam \Reg[17][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N30
cycloneive_lcell_comb \Mux57~0 (
// Equation(s):
// \Mux57~0_combout  = (ifid_ifinstr_o_19 & (((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[21][6]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[17][6]~q )))))

	.dataa(\Reg[21][6]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[17][6]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux57~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~0 .lut_mask = 16'hEE30;
defparam \Mux57~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N20
cycloneive_lcell_comb \Mux57~1 (
// Equation(s):
// \Mux57~1_combout  = (ifid_ifinstr_o_19 & ((\Mux57~0_combout  & ((\Reg[29][6]~q ))) # (!\Mux57~0_combout  & (\Reg[25][6]~q )))) # (!ifid_ifinstr_o_19 & (((\Mux57~0_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[25][6]~q ),
	.datac(\Mux57~0_combout ),
	.datad(\Reg[29][6]~q ),
	.cin(gnd),
	.combout(\Mux57~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~1 .lut_mask = 16'hF858;
defparam \Mux57~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N8
cycloneive_lcell_comb \Mux57~4 (
// Equation(s):
// \Mux57~4_combout  = (ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18) # ((\Reg[24][6]~q )))) # (!ifid_ifinstr_o_19 & (!ifid_ifinstr_o_18 & (\Reg[16][6]~q )))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[16][6]~q ),
	.datad(\Reg[24][6]~q ),
	.cin(gnd),
	.combout(\Mux57~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~4 .lut_mask = 16'hBA98;
defparam \Mux57~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N14
cycloneive_lcell_comb \Mux57~5 (
// Equation(s):
// \Mux57~5_combout  = (\Mux57~4_combout  & (((\Reg[28][6]~q ) # (!ifid_ifinstr_o_18)))) # (!\Mux57~4_combout  & (\Reg[20][6]~q  & ((ifid_ifinstr_o_18))))

	.dataa(\Reg[20][6]~q ),
	.datab(\Reg[28][6]~q ),
	.datac(\Mux57~4_combout ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux57~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~5 .lut_mask = 16'hCAF0;
defparam \Mux57~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N19
dffeas \Reg[30][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][6] .is_wysiwyg = "true";
defparam \Reg[30][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N2
cycloneive_lcell_comb \Mux57~2 (
// Equation(s):
// \Mux57~2_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[26][6]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[18][6]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[18][6]~q ),
	.datac(\Reg[26][6]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux57~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~2 .lut_mask = 16'hFA44;
defparam \Mux57~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N18
cycloneive_lcell_comb \Mux57~3 (
// Equation(s):
// \Mux57~3_combout  = (ifid_ifinstr_o_18 & ((\Mux57~2_combout  & ((\Reg[30][6]~q ))) # (!\Mux57~2_combout  & (\Reg[22][6]~q )))) # (!ifid_ifinstr_o_18 & (((\Mux57~2_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[22][6]~q ),
	.datac(\Reg[30][6]~q ),
	.datad(\Mux57~2_combout ),
	.cin(gnd),
	.combout(\Mux57~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~3 .lut_mask = 16'hF588;
defparam \Mux57~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N10
cycloneive_lcell_comb \Mux57~6 (
// Equation(s):
// \Mux57~6_combout  = (ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16) # ((\Mux57~3_combout )))) # (!ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & (\Mux57~5_combout )))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux57~5_combout ),
	.datad(\Mux57~3_combout ),
	.cin(gnd),
	.combout(\Mux57~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~6 .lut_mask = 16'hBA98;
defparam \Mux57~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N20
cycloneive_lcell_comb \Mux57~10 (
// Equation(s):
// \Mux57~10_combout  = (ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16) # ((\Reg[10][6]~q )))) # (!ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & ((\Reg[8][6]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[10][6]~q ),
	.datad(\Reg[8][6]~q ),
	.cin(gnd),
	.combout(\Mux57~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~10 .lut_mask = 16'hB9A8;
defparam \Mux57~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N16
cycloneive_lcell_comb \Mux57~11 (
// Equation(s):
// \Mux57~11_combout  = (ifid_ifinstr_o_16 & ((\Mux57~10_combout  & ((\Reg[11][6]~q ))) # (!\Mux57~10_combout  & (\Reg[9][6]~q )))) # (!ifid_ifinstr_o_16 & (\Mux57~10_combout ))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux57~10_combout ),
	.datac(\Reg[9][6]~q ),
	.datad(\Reg[11][6]~q ),
	.cin(gnd),
	.combout(\Mux57~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~11 .lut_mask = 16'hEC64;
defparam \Mux57~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y37_N8
cycloneive_lcell_comb \Mux57~17 (
// Equation(s):
// \Mux57~17_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[13][6]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[12][6]~q ))))

	.dataa(\Reg[12][6]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[13][6]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux57~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~17 .lut_mask = 16'hFC22;
defparam \Mux57~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N4
cycloneive_lcell_comb \Mux57~18 (
// Equation(s):
// \Mux57~18_combout  = (ifid_ifinstr_o_17 & ((\Mux57~17_combout  & (\Reg[15][6]~q )) # (!\Mux57~17_combout  & ((\Reg[14][6]~q ))))) # (!ifid_ifinstr_o_17 & (((\Mux57~17_combout ))))

	.dataa(\Reg[15][6]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[14][6]~q ),
	.datad(\Mux57~17_combout ),
	.cin(gnd),
	.combout(\Mux57~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~18 .lut_mask = 16'hBBC0;
defparam \Mux57~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N18
cycloneive_lcell_comb \Mux57~12 (
// Equation(s):
// \Mux57~12_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[5][6]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[4][6]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[5][6]~q ),
	.datac(\Reg[4][6]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux57~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~12 .lut_mask = 16'hEE50;
defparam \Mux57~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N10
cycloneive_lcell_comb \Mux57~13 (
// Equation(s):
// \Mux57~13_combout  = (ifid_ifinstr_o_17 & ((\Mux57~12_combout  & (\Reg[7][6]~q )) # (!\Mux57~12_combout  & ((\Reg[6][6]~q ))))) # (!ifid_ifinstr_o_17 & (\Mux57~12_combout ))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux57~12_combout ),
	.datac(\Reg[7][6]~q ),
	.datad(\Reg[6][6]~q ),
	.cin(gnd),
	.combout(\Mux57~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~13 .lut_mask = 16'hE6C4;
defparam \Mux57~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N7
dffeas \Reg[1][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat7),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][6] .is_wysiwyg = "true";
defparam \Reg[1][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N6
cycloneive_lcell_comb \Mux57~14 (
// Equation(s):
// \Mux57~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][6]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][6]~q )))))

	.dataa(\Reg[3][6]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[1][6]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux57~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~14 .lut_mask = 16'hB800;
defparam \Mux57~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N2
cycloneive_lcell_comb \Mux57~15 (
// Equation(s):
// \Mux57~15_combout  = (\Mux57~14_combout ) # ((\Reg[2][6]~q  & (!ifid_ifinstr_o_16 & ifid_ifinstr_o_17)))

	.dataa(\Reg[2][6]~q ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux57~14_combout ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux57~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~15 .lut_mask = 16'hF2F0;
defparam \Mux57~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N28
cycloneive_lcell_comb \Mux57~16 (
// Equation(s):
// \Mux57~16_combout  = (ifid_ifinstr_o_18 & ((\Mux57~13_combout ) # ((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (((!ifid_ifinstr_o_19 & \Mux57~15_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux57~13_combout ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux57~15_combout ),
	.cin(gnd),
	.combout(\Mux57~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~16 .lut_mask = 16'hADA8;
defparam \Mux57~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N8
cycloneive_lcell_comb \Reg[24][7]~feeder (
// Equation(s):
// \Reg[24][7]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat6),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[24][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[24][7]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[24][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N9
dffeas \Reg[24][7] (
	.clk(!CLK),
	.d(\Reg[24][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][7] .is_wysiwyg = "true";
defparam \Reg[24][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y33_N11
dffeas \Reg[16][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][7] .is_wysiwyg = "true";
defparam \Reg[16][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N28
cycloneive_lcell_comb \Mux56~4 (
// Equation(s):
// \Mux56~4_combout  = (ifid_ifinstr_o_19 & (((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Reg[20][7]~q ))) # (!ifid_ifinstr_o_18 & (\Reg[16][7]~q ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[16][7]~q ),
	.datac(\Reg[20][7]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux56~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~4 .lut_mask = 16'hFA44;
defparam \Mux56~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N22
cycloneive_lcell_comb \Mux56~5 (
// Equation(s):
// \Mux56~5_combout  = (ifid_ifinstr_o_19 & ((\Mux56~4_combout  & (\Reg[28][7]~q )) # (!\Mux56~4_combout  & ((\Reg[24][7]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux56~4_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[28][7]~q ),
	.datac(\Reg[24][7]~q ),
	.datad(\Mux56~4_combout ),
	.cin(gnd),
	.combout(\Mux56~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~5 .lut_mask = 16'hDDA0;
defparam \Mux56~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N12
cycloneive_lcell_comb \Mux56~2 (
// Equation(s):
// \Mux56~2_combout  = (ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19) # ((\Reg[22][7]~q )))) # (!ifid_ifinstr_o_18 & (!ifid_ifinstr_o_19 & (\Reg[18][7]~q )))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[18][7]~q ),
	.datad(\Reg[22][7]~q ),
	.cin(gnd),
	.combout(\Mux56~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~2 .lut_mask = 16'hBA98;
defparam \Mux56~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N31
dffeas \Reg[30][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][7] .is_wysiwyg = "true";
defparam \Reg[30][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N30
cycloneive_lcell_comb \Mux56~3 (
// Equation(s):
// \Mux56~3_combout  = (ifid_ifinstr_o_19 & ((\Mux56~2_combout  & (\Reg[30][7]~q )) # (!\Mux56~2_combout  & ((\Reg[26][7]~q ))))) # (!ifid_ifinstr_o_19 & (\Mux56~2_combout ))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Mux56~2_combout ),
	.datac(\Reg[30][7]~q ),
	.datad(\Reg[26][7]~q ),
	.cin(gnd),
	.combout(\Mux56~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~3 .lut_mask = 16'hE6C4;
defparam \Mux56~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N12
cycloneive_lcell_comb \Mux56~6 (
// Equation(s):
// \Mux56~6_combout  = (ifid_ifinstr_o_16 & (((ifid_ifinstr_o_17)))) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Mux56~3_combout ))) # (!ifid_ifinstr_o_17 & (\Mux56~5_combout ))))

	.dataa(\Mux56~5_combout ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux56~3_combout ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux56~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~6 .lut_mask = 16'hFC22;
defparam \Mux56~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N10
cycloneive_lcell_comb \Mux56~0 (
// Equation(s):
// \Mux56~0_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Reg[25][7]~q )) # (!ifid_ifinstr_o_19 & ((\Reg[17][7]~q )))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[25][7]~q ),
	.datac(\Reg[17][7]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux56~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~0 .lut_mask = 16'hEE50;
defparam \Mux56~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N12
cycloneive_lcell_comb \Reg[21][7]~feeder (
// Equation(s):
// \Reg[21][7]~feeder_combout  = \wdat~13_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat6),
	.cin(gnd),
	.combout(\Reg[21][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[21][7]~feeder .lut_mask = 16'hFF00;
defparam \Reg[21][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y38_N13
dffeas \Reg[21][7] (
	.clk(!CLK),
	.d(\Reg[21][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[21][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[21][7] .is_wysiwyg = "true";
defparam \Reg[21][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N2
cycloneive_lcell_comb \Mux56~1 (
// Equation(s):
// \Mux56~1_combout  = (\Mux56~0_combout  & ((\Reg[29][7]~q ) # ((!ifid_ifinstr_o_18)))) # (!\Mux56~0_combout  & (((ifid_ifinstr_o_18 & \Reg[21][7]~q ))))

	.dataa(\Mux56~0_combout ),
	.datab(\Reg[29][7]~q ),
	.datac(ifid_ifinstr_o_18),
	.datad(\Reg[21][7]~q ),
	.cin(gnd),
	.combout(\Mux56~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~1 .lut_mask = 16'hDA8A;
defparam \Mux56~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N22
cycloneive_lcell_comb \Mux56~7 (
// Equation(s):
// \Mux56~7_combout  = (ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18) # ((\Reg[27][7]~q )))) # (!ifid_ifinstr_o_19 & (!ifid_ifinstr_o_18 & (\Reg[19][7]~q )))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[19][7]~q ),
	.datad(\Reg[27][7]~q ),
	.cin(gnd),
	.combout(\Mux56~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~7 .lut_mask = 16'hBA98;
defparam \Mux56~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N18
cycloneive_lcell_comb \Mux56~8 (
// Equation(s):
// \Mux56~8_combout  = (ifid_ifinstr_o_18 & ((\Mux56~7_combout  & (\Reg[31][7]~q )) # (!\Mux56~7_combout  & ((\Reg[23][7]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux56~7_combout ))))

	.dataa(\Reg[31][7]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[23][7]~q ),
	.datad(\Mux56~7_combout ),
	.cin(gnd),
	.combout(\Mux56~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~8 .lut_mask = 16'hBBC0;
defparam \Mux56~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N17
dffeas \Reg[5][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][7] .is_wysiwyg = "true";
defparam \Reg[5][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N11
dffeas \Reg[4][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][7] .is_wysiwyg = "true";
defparam \Reg[4][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N16
cycloneive_lcell_comb \Mux56~10 (
// Equation(s):
// \Mux56~10_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[5][7]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[4][7]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[5][7]~q ),
	.datad(\Reg[4][7]~q ),
	.cin(gnd),
	.combout(\Mux56~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~10 .lut_mask = 16'hD9C8;
defparam \Mux56~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N8
cycloneive_lcell_comb \Mux56~11 (
// Equation(s):
// \Mux56~11_combout  = (\Mux56~10_combout  & ((\Reg[7][7]~q ) # ((!ifid_ifinstr_o_17)))) # (!\Mux56~10_combout  & (((\Reg[6][7]~q  & ifid_ifinstr_o_17))))

	.dataa(\Mux56~10_combout ),
	.datab(\Reg[7][7]~q ),
	.datac(\Reg[6][7]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux56~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~11 .lut_mask = 16'hD8AA;
defparam \Mux56~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N23
dffeas \Reg[12][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][7] .is_wysiwyg = "true";
defparam \Reg[12][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N22
cycloneive_lcell_comb \Mux56~17 (
// Equation(s):
// \Mux56~17_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[13][7]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[12][7]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[13][7]~q ),
	.datac(\Reg[12][7]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux56~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~17 .lut_mask = 16'hEE50;
defparam \Mux56~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N8
cycloneive_lcell_comb \Mux56~18 (
// Equation(s):
// \Mux56~18_combout  = (\Mux56~17_combout  & ((\Reg[15][7]~q ) # ((!ifid_ifinstr_o_17)))) # (!\Mux56~17_combout  & (((\Reg[14][7]~q  & ifid_ifinstr_o_17))))

	.dataa(\Mux56~17_combout ),
	.datab(\Reg[15][7]~q ),
	.datac(\Reg[14][7]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux56~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~18 .lut_mask = 16'hD8AA;
defparam \Mux56~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y31_N31
dffeas \Reg[8][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat6),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][7] .is_wysiwyg = "true";
defparam \Reg[8][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N30
cycloneive_lcell_comb \Mux56~12 (
// Equation(s):
// \Mux56~12_combout  = (ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16) # ((\Reg[10][7]~q )))) # (!ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & (\Reg[8][7]~q )))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[8][7]~q ),
	.datad(\Reg[10][7]~q ),
	.cin(gnd),
	.combout(\Mux56~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~12 .lut_mask = 16'hBA98;
defparam \Mux56~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N18
cycloneive_lcell_comb \Mux56~13 (
// Equation(s):
// \Mux56~13_combout  = (\Mux56~12_combout  & (((\Reg[11][7]~q ) # (!ifid_ifinstr_o_16)))) # (!\Mux56~12_combout  & (\Reg[9][7]~q  & ((ifid_ifinstr_o_16))))

	.dataa(\Reg[9][7]~q ),
	.datab(\Mux56~12_combout ),
	.datac(\Reg[11][7]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux56~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~13 .lut_mask = 16'hE2CC;
defparam \Mux56~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N24
cycloneive_lcell_comb \Mux56~14 (
// Equation(s):
// \Mux56~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][7]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][7]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[3][7]~q ),
	.datad(\Reg[1][7]~q ),
	.cin(gnd),
	.combout(\Mux56~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~14 .lut_mask = 16'hA280;
defparam \Mux56~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N24
cycloneive_lcell_comb \Mux56~15 (
// Equation(s):
// \Mux56~15_combout  = (\Mux56~14_combout ) # ((!ifid_ifinstr_o_16 & (ifid_ifinstr_o_17 & \Reg[2][7]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[2][7]~q ),
	.datad(\Mux56~14_combout ),
	.cin(gnd),
	.combout(\Mux56~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~15 .lut_mask = 16'hFF40;
defparam \Mux56~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N20
cycloneive_lcell_comb \Mux56~16 (
// Equation(s):
// \Mux56~16_combout  = (ifid_ifinstr_o_19 & ((\Mux56~13_combout ) # ((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & (((!ifid_ifinstr_o_18 & \Mux56~15_combout ))))

	.dataa(\Mux56~13_combout ),
	.datab(ifid_ifinstr_o_19),
	.datac(ifid_ifinstr_o_18),
	.datad(\Mux56~15_combout ),
	.cin(gnd),
	.combout(\Mux56~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~16 .lut_mask = 16'hCBC8;
defparam \Mux56~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N30
cycloneive_lcell_comb \Reg[19][8]~feeder (
// Equation(s):
// \Reg[19][8]~feeder_combout  = \wdat~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat5),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[19][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[19][8]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[19][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N31
dffeas \Reg[19][8] (
	.clk(!CLK),
	.d(\Reg[19][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[19][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[19][8] .is_wysiwyg = "true";
defparam \Reg[19][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N20
cycloneive_lcell_comb \Mux55~7 (
// Equation(s):
// \Mux55~7_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[23][8]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[19][8]~q )))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[23][8]~q ),
	.datad(\Reg[19][8]~q ),
	.cin(gnd),
	.combout(\Mux55~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~7 .lut_mask = 16'hD9C8;
defparam \Mux55~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N24
cycloneive_lcell_comb \Mux55~8 (
// Equation(s):
// \Mux55~8_combout  = (ifid_ifinstr_o_19 & ((\Mux55~7_combout  & (\Reg[31][8]~q )) # (!\Mux55~7_combout  & ((\Reg[27][8]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux55~7_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[31][8]~q ),
	.datac(\Mux55~7_combout ),
	.datad(\Reg[27][8]~q ),
	.cin(gnd),
	.combout(\Mux55~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~8 .lut_mask = 16'hDAD0;
defparam \Mux55~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N2
cycloneive_lcell_comb \Mux55~0 (
// Equation(s):
// \Mux55~0_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19) # (\Reg[21][8]~q )))) # (!ifid_ifinstr_o_18 & (\Reg[17][8]~q  & (!ifid_ifinstr_o_19)))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[17][8]~q ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Reg[21][8]~q ),
	.cin(gnd),
	.combout(\Mux55~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~0 .lut_mask = 16'hAEA4;
defparam \Mux55~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N14
cycloneive_lcell_comb \Mux55~1 (
// Equation(s):
// \Mux55~1_combout  = (ifid_ifinstr_o_19 & ((\Mux55~0_combout  & (\Reg[29][8]~q )) # (!\Mux55~0_combout  & ((\Reg[25][8]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux55~0_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[29][8]~q ),
	.datac(\Mux55~0_combout ),
	.datad(\Reg[25][8]~q ),
	.cin(gnd),
	.combout(\Mux55~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~1 .lut_mask = 16'hDAD0;
defparam \Mux55~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N3
dffeas \Reg[28][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat5),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][8] .is_wysiwyg = "true";
defparam \Reg[28][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N28
cycloneive_lcell_comb \Mux55~4 (
// Equation(s):
// \Mux55~4_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[24][8]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[16][8]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[16][8]~q ),
	.datac(\Reg[24][8]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux55~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~4 .lut_mask = 16'hFA44;
defparam \Mux55~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N2
cycloneive_lcell_comb \Mux55~5 (
// Equation(s):
// \Mux55~5_combout  = (ifid_ifinstr_o_18 & ((\Mux55~4_combout  & ((\Reg[28][8]~q ))) # (!\Mux55~4_combout  & (\Reg[20][8]~q )))) # (!ifid_ifinstr_o_18 & (((\Mux55~4_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[20][8]~q ),
	.datac(\Reg[28][8]~q ),
	.datad(\Mux55~4_combout ),
	.cin(gnd),
	.combout(\Mux55~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~5 .lut_mask = 16'hF588;
defparam \Mux55~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N6
cycloneive_lcell_comb \Mux55~2 (
// Equation(s):
// \Mux55~2_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Reg[26][8]~q )) # (!ifid_ifinstr_o_19 & ((\Reg[18][8]~q )))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[26][8]~q ),
	.datad(\Reg[18][8]~q ),
	.cin(gnd),
	.combout(\Mux55~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~2 .lut_mask = 16'hD9C8;
defparam \Mux55~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N14
cycloneive_lcell_comb \Mux55~3 (
// Equation(s):
// \Mux55~3_combout  = (ifid_ifinstr_o_18 & ((\Mux55~2_combout  & ((\Reg[30][8]~q ))) # (!\Mux55~2_combout  & (\Reg[22][8]~q )))) # (!ifid_ifinstr_o_18 & (((\Mux55~2_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[22][8]~q ),
	.datac(\Reg[30][8]~q ),
	.datad(\Mux55~2_combout ),
	.cin(gnd),
	.combout(\Mux55~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~3 .lut_mask = 16'hF588;
defparam \Mux55~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N6
cycloneive_lcell_comb \Mux55~6 (
// Equation(s):
// \Mux55~6_combout  = (ifid_ifinstr_o_16 & (((ifid_ifinstr_o_17)))) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Mux55~3_combout ))) # (!ifid_ifinstr_o_17 & (\Mux55~5_combout ))))

	.dataa(\Mux55~5_combout ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux55~3_combout ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux55~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~6 .lut_mask = 16'hFC22;
defparam \Mux55~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N22
cycloneive_lcell_comb \Mux55~17 (
// Equation(s):
// \Mux55~17_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17) # ((\Reg[13][8]~q )))) # (!ifid_ifinstr_o_16 & (!ifid_ifinstr_o_17 & (\Reg[12][8]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[12][8]~q ),
	.datad(\Reg[13][8]~q ),
	.cin(gnd),
	.combout(\Mux55~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~17 .lut_mask = 16'hBA98;
defparam \Mux55~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y37_N28
cycloneive_lcell_comb \Mux55~18 (
// Equation(s):
// \Mux55~18_combout  = (\Mux55~17_combout  & ((\Reg[15][8]~q ) # ((!ifid_ifinstr_o_17)))) # (!\Mux55~17_combout  & (((\Reg[14][8]~q  & ifid_ifinstr_o_17))))

	.dataa(\Reg[15][8]~q ),
	.datab(\Mux55~17_combout ),
	.datac(\Reg[14][8]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux55~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~18 .lut_mask = 16'hB8CC;
defparam \Mux55~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N4
cycloneive_lcell_comb \Mux55~10 (
// Equation(s):
// \Mux55~10_combout  = (ifid_ifinstr_o_16 & (((ifid_ifinstr_o_17)))) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[10][8]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[8][8]~q ))))

	.dataa(\Reg[8][8]~q ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[10][8]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux55~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~10 .lut_mask = 16'hFC22;
defparam \Mux55~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N16
cycloneive_lcell_comb \Reg[9][8]~feeder (
// Equation(s):
// \Reg[9][8]~feeder_combout  = \wdat~11_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat5),
	.cin(gnd),
	.combout(\Reg[9][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[9][8]~feeder .lut_mask = 16'hFF00;
defparam \Reg[9][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y35_N17
dffeas \Reg[9][8] (
	.clk(!CLK),
	.d(\Reg[9][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][8] .is_wysiwyg = "true";
defparam \Reg[9][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N28
cycloneive_lcell_comb \Mux55~11 (
// Equation(s):
// \Mux55~11_combout  = (ifid_ifinstr_o_16 & ((\Mux55~10_combout  & (\Reg[11][8]~q )) # (!\Mux55~10_combout  & ((\Reg[9][8]~q ))))) # (!ifid_ifinstr_o_16 & (\Mux55~10_combout ))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux55~10_combout ),
	.datac(\Reg[11][8]~q ),
	.datad(\Reg[9][8]~q ),
	.cin(gnd),
	.combout(\Mux55~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~11 .lut_mask = 16'hE6C4;
defparam \Mux55~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N4
cycloneive_lcell_comb \Mux55~14 (
// Equation(s):
// \Mux55~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[3][8]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[1][8]~q ))))

	.dataa(\Reg[1][8]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[3][8]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux55~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~14 .lut_mask = 16'hE200;
defparam \Mux55~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N0
cycloneive_lcell_comb \Mux55~15 (
// Equation(s):
// \Mux55~15_combout  = (\Mux55~14_combout ) # ((!ifid_ifinstr_o_16 & (ifid_ifinstr_o_17 & \Reg[2][8]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[2][8]~q ),
	.datad(\Mux55~14_combout ),
	.cin(gnd),
	.combout(\Mux55~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~15 .lut_mask = 16'hFF40;
defparam \Mux55~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N22
cycloneive_lcell_comb \Mux55~12 (
// Equation(s):
// \Mux55~12_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[5][8]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[4][8]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[5][8]~q ),
	.datac(\Reg[4][8]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux55~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~12 .lut_mask = 16'hEE50;
defparam \Mux55~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N6
cycloneive_lcell_comb \Mux55~13 (
// Equation(s):
// \Mux55~13_combout  = (ifid_ifinstr_o_17 & ((\Mux55~12_combout  & ((\Reg[7][8]~q ))) # (!\Mux55~12_combout  & (\Reg[6][8]~q )))) # (!ifid_ifinstr_o_17 & (((\Mux55~12_combout ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[6][8]~q ),
	.datac(\Reg[7][8]~q ),
	.datad(\Mux55~12_combout ),
	.cin(gnd),
	.combout(\Mux55~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~13 .lut_mask = 16'hF588;
defparam \Mux55~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N30
cycloneive_lcell_comb \Mux55~16 (
// Equation(s):
// \Mux55~16_combout  = (ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19) # ((\Mux55~13_combout )))) # (!ifid_ifinstr_o_18 & (!ifid_ifinstr_o_19 & (\Mux55~15_combout )))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Mux55~15_combout ),
	.datad(\Mux55~13_combout ),
	.cin(gnd),
	.combout(\Mux55~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~16 .lut_mask = 16'hBA98;
defparam \Mux55~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N8
cycloneive_lcell_comb \Mux36~7 (
// Equation(s):
// \Mux36~7_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Reg[27][27]~q )) # (!ifid_ifinstr_o_19 & ((\Reg[19][27]~q )))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[27][27]~q ),
	.datad(\Reg[19][27]~q ),
	.cin(gnd),
	.combout(\Mux36~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~7 .lut_mask = 16'hD9C8;
defparam \Mux36~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N22
cycloneive_lcell_comb \Mux36~8 (
// Equation(s):
// \Mux36~8_combout  = (ifid_ifinstr_o_18 & ((\Mux36~7_combout  & (\Reg[31][27]~q )) # (!\Mux36~7_combout  & ((\Reg[23][27]~q ))))) # (!ifid_ifinstr_o_18 & (\Mux36~7_combout ))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux36~7_combout ),
	.datac(\Reg[31][27]~q ),
	.datad(\Reg[23][27]~q ),
	.cin(gnd),
	.combout(\Mux36~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~8 .lut_mask = 16'hE6C4;
defparam \Mux36~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y38_N4
cycloneive_lcell_comb \Mux36~0 (
// Equation(s):
// \Mux36~0_combout  = (ifid_ifinstr_o_19 & (((\Reg[25][27]~q ) # (ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & (\Reg[17][27]~q  & ((!ifid_ifinstr_o_18))))

	.dataa(\Reg[17][27]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[25][27]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux36~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~0 .lut_mask = 16'hCCE2;
defparam \Mux36~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y38_N14
cycloneive_lcell_comb \Mux36~1 (
// Equation(s):
// \Mux36~1_combout  = (\Mux36~0_combout  & (((\Reg[29][27]~q )) # (!ifid_ifinstr_o_18))) # (!\Mux36~0_combout  & (ifid_ifinstr_o_18 & (\Reg[21][27]~q )))

	.dataa(\Mux36~0_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[21][27]~q ),
	.datad(\Reg[29][27]~q ),
	.cin(gnd),
	.combout(\Mux36~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~1 .lut_mask = 16'hEA62;
defparam \Mux36~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N15
dffeas \Reg[16][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat22),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][27] .is_wysiwyg = "true";
defparam \Reg[16][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N14
cycloneive_lcell_comb \Mux36~4 (
// Equation(s):
// \Mux36~4_combout  = (ifid_ifinstr_o_18 & ((\Reg[20][27]~q ) # ((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (((\Reg[16][27]~q  & !ifid_ifinstr_o_19))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[20][27]~q ),
	.datac(\Reg[16][27]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux36~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~4 .lut_mask = 16'hAAD8;
defparam \Mux36~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N18
cycloneive_lcell_comb \Mux36~5 (
// Equation(s):
// \Mux36~5_combout  = (ifid_ifinstr_o_19 & ((\Mux36~4_combout  & (\Reg[28][27]~q )) # (!\Mux36~4_combout  & ((\Reg[24][27]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux36~4_combout ))))

	.dataa(\Reg[28][27]~q ),
	.datab(\Reg[24][27]~q ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux36~4_combout ),
	.cin(gnd),
	.combout(\Mux36~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~5 .lut_mask = 16'hAFC0;
defparam \Mux36~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N2
cycloneive_lcell_comb \Mux36~2 (
// Equation(s):
// \Mux36~2_combout  = (ifid_ifinstr_o_18 & (((\Reg[22][27]~q ) # (ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (\Reg[18][27]~q  & ((!ifid_ifinstr_o_19))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[18][27]~q ),
	.datac(\Reg[22][27]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux36~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~2 .lut_mask = 16'hAAE4;
defparam \Mux36~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N30
cycloneive_lcell_comb \Reg[30][27]~feeder (
// Equation(s):
// \Reg[30][27]~feeder_combout  = \wdat~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat22),
	.cin(gnd),
	.combout(\Reg[30][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[30][27]~feeder .lut_mask = 16'hFF00;
defparam \Reg[30][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N31
dffeas \Reg[30][27] (
	.clk(!CLK),
	.d(\Reg[30][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][27] .is_wysiwyg = "true";
defparam \Reg[30][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N14
cycloneive_lcell_comb \Mux36~3 (
// Equation(s):
// \Mux36~3_combout  = (ifid_ifinstr_o_19 & ((\Mux36~2_combout  & (\Reg[30][27]~q )) # (!\Mux36~2_combout  & ((\Reg[26][27]~q ))))) # (!ifid_ifinstr_o_19 & (\Mux36~2_combout ))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Mux36~2_combout ),
	.datac(\Reg[30][27]~q ),
	.datad(\Reg[26][27]~q ),
	.cin(gnd),
	.combout(\Mux36~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~3 .lut_mask = 16'hE6C4;
defparam \Mux36~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N12
cycloneive_lcell_comb \Mux36~6 (
// Equation(s):
// \Mux36~6_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16) # (\Mux36~3_combout )))) # (!ifid_ifinstr_o_17 & (\Mux36~5_combout  & (!ifid_ifinstr_o_16)))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux36~5_combout ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux36~3_combout ),
	.cin(gnd),
	.combout(\Mux36~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~6 .lut_mask = 16'hAEA4;
defparam \Mux36~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N22
cycloneive_lcell_comb \Reg[13][27]~feeder (
// Equation(s):
// \Reg[13][27]~feeder_combout  = \wdat~47_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat22),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[13][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[13][27]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[13][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N23
dffeas \Reg[13][27] (
	.clk(!CLK),
	.d(\Reg[13][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[13][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[13][27] .is_wysiwyg = "true";
defparam \Reg[13][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N26
cycloneive_lcell_comb \Mux36~17 (
// Equation(s):
// \Mux36~17_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17) # ((\Reg[13][27]~q )))) # (!ifid_ifinstr_o_16 & (!ifid_ifinstr_o_17 & (\Reg[12][27]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[12][27]~q ),
	.datad(\Reg[13][27]~q ),
	.cin(gnd),
	.combout(\Mux36~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~17 .lut_mask = 16'hBA98;
defparam \Mux36~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N16
cycloneive_lcell_comb \Mux36~18 (
// Equation(s):
// \Mux36~18_combout  = (ifid_ifinstr_o_17 & ((\Mux36~17_combout  & ((\Reg[15][27]~q ))) # (!\Mux36~17_combout  & (\Reg[14][27]~q )))) # (!ifid_ifinstr_o_17 & (((\Mux36~17_combout ))))

	.dataa(\Reg[14][27]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux36~17_combout ),
	.datad(\Reg[15][27]~q ),
	.cin(gnd),
	.combout(\Mux36~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~18 .lut_mask = 16'hF838;
defparam \Mux36~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N24
cycloneive_lcell_comb \Mux36~10 (
// Equation(s):
// \Mux36~10_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[5][27]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[4][27]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[5][27]~q ),
	.datad(\Reg[4][27]~q ),
	.cin(gnd),
	.combout(\Mux36~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~10 .lut_mask = 16'hD9C8;
defparam \Mux36~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N8
cycloneive_lcell_comb \Mux36~11 (
// Equation(s):
// \Mux36~11_combout  = (\Mux36~10_combout  & ((\Reg[7][27]~q ) # ((!ifid_ifinstr_o_17)))) # (!\Mux36~10_combout  & (((\Reg[6][27]~q  & ifid_ifinstr_o_17))))

	.dataa(\Reg[7][27]~q ),
	.datab(\Mux36~10_combout ),
	.datac(\Reg[6][27]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux36~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~11 .lut_mask = 16'hB8CC;
defparam \Mux36~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N6
cycloneive_lcell_comb \Mux36~12 (
// Equation(s):
// \Mux36~12_combout  = (ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16) # ((\Reg[10][27]~q )))) # (!ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & (\Reg[8][27]~q )))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[8][27]~q ),
	.datad(\Reg[10][27]~q ),
	.cin(gnd),
	.combout(\Mux36~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~12 .lut_mask = 16'hBA98;
defparam \Mux36~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N18
cycloneive_lcell_comb \Mux36~13 (
// Equation(s):
// \Mux36~13_combout  = (\Mux36~12_combout  & (((\Reg[11][27]~q ) # (!ifid_ifinstr_o_16)))) # (!\Mux36~12_combout  & (\Reg[9][27]~q  & ((ifid_ifinstr_o_16))))

	.dataa(\Reg[9][27]~q ),
	.datab(\Mux36~12_combout ),
	.datac(\Reg[11][27]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux36~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~13 .lut_mask = 16'hE2CC;
defparam \Mux36~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N2
cycloneive_lcell_comb \Mux36~14 (
// Equation(s):
// \Mux36~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][27]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][27]~q )))))

	.dataa(\Reg[3][27]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[1][27]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux36~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~14 .lut_mask = 16'hB800;
defparam \Mux36~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N26
cycloneive_lcell_comb \Mux36~15 (
// Equation(s):
// \Mux36~15_combout  = (\Mux36~14_combout ) # ((!ifid_ifinstr_o_16 & (ifid_ifinstr_o_17 & \Reg[2][27]~q )))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[2][27]~q ),
	.datad(\Mux36~14_combout ),
	.cin(gnd),
	.combout(\Mux36~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~15 .lut_mask = 16'hFF40;
defparam \Mux36~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N28
cycloneive_lcell_comb \Mux36~16 (
// Equation(s):
// \Mux36~16_combout  = (ifid_ifinstr_o_19 & ((\Mux36~13_combout ) # ((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & (((!ifid_ifinstr_o_18 & \Mux36~15_combout ))))

	.dataa(\Mux36~13_combout ),
	.datab(ifid_ifinstr_o_19),
	.datac(ifid_ifinstr_o_18),
	.datad(\Mux36~15_combout ),
	.cin(gnd),
	.combout(\Mux36~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~16 .lut_mask = 16'hCBC8;
defparam \Mux36~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N22
cycloneive_lcell_comb \Reg[25][28]~feeder (
// Equation(s):
// \Reg[25][28]~feeder_combout  = \wdat~43_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat20),
	.cin(gnd),
	.combout(\Reg[25][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[25][28]~feeder .lut_mask = 16'hFF00;
defparam \Reg[25][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y37_N23
dffeas \Reg[25][28] (
	.clk(!CLK),
	.d(\Reg[25][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~2_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[25][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[25][28] .is_wysiwyg = "true";
defparam \Reg[25][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N24
cycloneive_lcell_comb \Mux35~0 (
// Equation(s):
// \Mux35~0_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19) # (\Reg[21][28]~q )))) # (!ifid_ifinstr_o_18 & (\Reg[17][28]~q  & (!ifid_ifinstr_o_19)))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[17][28]~q ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Reg[21][28]~q ),
	.cin(gnd),
	.combout(\Mux35~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~0 .lut_mask = 16'hAEA4;
defparam \Mux35~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N14
cycloneive_lcell_comb \Mux35~1 (
// Equation(s):
// \Mux35~1_combout  = (ifid_ifinstr_o_19 & ((\Mux35~0_combout  & (\Reg[29][28]~q )) # (!\Mux35~0_combout  & ((\Reg[25][28]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux35~0_combout ))))

	.dataa(\Reg[29][28]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[25][28]~q ),
	.datad(\Mux35~0_combout ),
	.cin(gnd),
	.combout(\Mux35~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~1 .lut_mask = 16'hBBC0;
defparam \Mux35~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N0
cycloneive_lcell_comb \Mux35~7 (
// Equation(s):
// \Mux35~7_combout  = (ifid_ifinstr_o_18 & (((\Reg[23][28]~q ) # (ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (\Reg[19][28]~q  & ((!ifid_ifinstr_o_19))))

	.dataa(\Reg[19][28]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[23][28]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux35~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~7 .lut_mask = 16'hCCE2;
defparam \Mux35~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N16
cycloneive_lcell_comb \Mux35~8 (
// Equation(s):
// \Mux35~8_combout  = (\Mux35~7_combout  & (((\Reg[31][28]~q ) # (!ifid_ifinstr_o_19)))) # (!\Mux35~7_combout  & (\Reg[27][28]~q  & ((ifid_ifinstr_o_19))))

	.dataa(\Mux35~7_combout ),
	.datab(\Reg[27][28]~q ),
	.datac(\Reg[31][28]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux35~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~8 .lut_mask = 16'hE4AA;
defparam \Mux35~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N16
cycloneive_lcell_comb \Mux35~2 (
// Equation(s):
// \Mux35~2_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Reg[26][28]~q )) # (!ifid_ifinstr_o_19 & ((\Reg[18][28]~q )))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[26][28]~q ),
	.datad(\Reg[18][28]~q ),
	.cin(gnd),
	.combout(\Mux35~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~2 .lut_mask = 16'hD9C8;
defparam \Mux35~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N4
cycloneive_lcell_comb \Mux35~3 (
// Equation(s):
// \Mux35~3_combout  = (ifid_ifinstr_o_18 & ((\Mux35~2_combout  & (\Reg[30][28]~q )) # (!\Mux35~2_combout  & ((\Reg[22][28]~q ))))) # (!ifid_ifinstr_o_18 & (\Mux35~2_combout ))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux35~2_combout ),
	.datac(\Reg[30][28]~q ),
	.datad(\Reg[22][28]~q ),
	.cin(gnd),
	.combout(\Mux35~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~3 .lut_mask = 16'hE6C4;
defparam \Mux35~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N14
cycloneive_lcell_comb \Mux35~5 (
// Equation(s):
// \Mux35~5_combout  = (\Mux35~4_combout  & (((\Reg[28][28]~q )) # (!ifid_ifinstr_o_18))) # (!\Mux35~4_combout  & (ifid_ifinstr_o_18 & ((\Reg[20][28]~q ))))

	.dataa(\Mux35~4_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[28][28]~q ),
	.datad(\Reg[20][28]~q ),
	.cin(gnd),
	.combout(\Mux35~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~5 .lut_mask = 16'hE6A2;
defparam \Mux35~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N2
cycloneive_lcell_comb \Mux35~6 (
// Equation(s):
// \Mux35~6_combout  = (ifid_ifinstr_o_17 & ((\Mux35~3_combout ) # ((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & (((!ifid_ifinstr_o_16 & \Mux35~5_combout ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux35~3_combout ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux35~5_combout ),
	.cin(gnd),
	.combout(\Mux35~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~6 .lut_mask = 16'hADA8;
defparam \Mux35~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N24
cycloneive_lcell_comb \Mux35~17 (
// Equation(s):
// \Mux35~17_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[13][28]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[12][28]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[12][28]~q ),
	.datad(\Reg[13][28]~q ),
	.cin(gnd),
	.combout(\Mux35~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~17 .lut_mask = 16'hDC98;
defparam \Mux35~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N6
cycloneive_lcell_comb \Mux35~18 (
// Equation(s):
// \Mux35~18_combout  = (\Mux35~17_combout  & (((\Reg[15][28]~q )) # (!ifid_ifinstr_o_17))) # (!\Mux35~17_combout  & (ifid_ifinstr_o_17 & ((\Reg[14][28]~q ))))

	.dataa(\Mux35~17_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[15][28]~q ),
	.datad(\Reg[14][28]~q ),
	.cin(gnd),
	.combout(\Mux35~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~18 .lut_mask = 16'hE6A2;
defparam \Mux35~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y31_N15
dffeas \Reg[8][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][28] .is_wysiwyg = "true";
defparam \Reg[8][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N17
dffeas \Reg[10][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat20),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][28] .is_wysiwyg = "true";
defparam \Reg[10][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N16
cycloneive_lcell_comb \Mux35~10 (
// Equation(s):
// \Mux35~10_combout  = (ifid_ifinstr_o_17 & (((\Reg[10][28]~q ) # (ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & (\Reg[8][28]~q  & ((!ifid_ifinstr_o_16))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[8][28]~q ),
	.datac(\Reg[10][28]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux35~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~10 .lut_mask = 16'hAAE4;
defparam \Mux35~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N24
cycloneive_lcell_comb \Mux35~11 (
// Equation(s):
// \Mux35~11_combout  = (\Mux35~10_combout  & ((\Reg[11][28]~q ) # ((!ifid_ifinstr_o_16)))) # (!\Mux35~10_combout  & (((\Reg[9][28]~q  & ifid_ifinstr_o_16))))

	.dataa(\Mux35~10_combout ),
	.datab(\Reg[11][28]~q ),
	.datac(\Reg[9][28]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux35~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~11 .lut_mask = 16'hD8AA;
defparam \Mux35~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N30
cycloneive_lcell_comb \Mux35~15 (
// Equation(s):
// \Mux35~15_combout  = (\Mux35~14_combout ) # ((ifid_ifinstr_o_17 & (\Reg[2][28]~q  & !ifid_ifinstr_o_16)))

	.dataa(\Mux35~14_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[2][28]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux35~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~15 .lut_mask = 16'hAAEA;
defparam \Mux35~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N12
cycloneive_lcell_comb \Mux35~13 (
// Equation(s):
// \Mux35~13_combout  = (\Mux35~12_combout  & (((\Reg[7][28]~q )) # (!ifid_ifinstr_o_17))) # (!\Mux35~12_combout  & (ifid_ifinstr_o_17 & ((\Reg[6][28]~q ))))

	.dataa(\Mux35~12_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[7][28]~q ),
	.datad(\Reg[6][28]~q ),
	.cin(gnd),
	.combout(\Mux35~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~13 .lut_mask = 16'hE6A2;
defparam \Mux35~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N26
cycloneive_lcell_comb \Mux35~16 (
// Equation(s):
// \Mux35~16_combout  = (ifid_ifinstr_o_19 & (((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Mux35~13_combout ))) # (!ifid_ifinstr_o_18 & (\Mux35~15_combout ))))

	.dataa(\Mux35~15_combout ),
	.datab(ifid_ifinstr_o_19),
	.datac(ifid_ifinstr_o_18),
	.datad(\Mux35~13_combout ),
	.cin(gnd),
	.combout(\Mux35~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~16 .lut_mask = 16'hF2C2;
defparam \Mux35~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N4
cycloneive_lcell_comb \Mux34~7 (
// Equation(s):
// \Mux34~7_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[27][29]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[19][29]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[19][29]~q ),
	.datac(\Reg[27][29]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux34~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~7 .lut_mask = 16'hFA44;
defparam \Mux34~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N10
cycloneive_lcell_comb \Mux34~8 (
// Equation(s):
// \Mux34~8_combout  = (ifid_ifinstr_o_18 & ((\Mux34~7_combout  & (\Reg[31][29]~q )) # (!\Mux34~7_combout  & ((\Reg[23][29]~q ))))) # (!ifid_ifinstr_o_18 & (\Mux34~7_combout ))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux34~7_combout ),
	.datac(\Reg[31][29]~q ),
	.datad(\Reg[23][29]~q ),
	.cin(gnd),
	.combout(\Mux34~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~8 .lut_mask = 16'hE6C4;
defparam \Mux34~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N0
cycloneive_lcell_comb \Mux34~0 (
// Equation(s):
// \Mux34~0_combout  = (ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18) # ((\Reg[25][29]~q )))) # (!ifid_ifinstr_o_19 & (!ifid_ifinstr_o_18 & (\Reg[17][29]~q )))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[17][29]~q ),
	.datad(\Reg[25][29]~q ),
	.cin(gnd),
	.combout(\Mux34~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~0 .lut_mask = 16'hBA98;
defparam \Mux34~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N16
cycloneive_lcell_comb \Mux34~1 (
// Equation(s):
// \Mux34~1_combout  = (\Mux34~0_combout  & (((\Reg[29][29]~q ) # (!ifid_ifinstr_o_18)))) # (!\Mux34~0_combout  & (\Reg[21][29]~q  & ((ifid_ifinstr_o_18))))

	.dataa(\Reg[21][29]~q ),
	.datab(\Mux34~0_combout ),
	.datac(\Reg[29][29]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux34~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~1 .lut_mask = 16'hE2CC;
defparam \Mux34~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N24
cycloneive_lcell_comb \Mux34~2 (
// Equation(s):
// \Mux34~2_combout  = (ifid_ifinstr_o_18 & (((\Reg[22][29]~q ) # (ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (\Reg[18][29]~q  & ((!ifid_ifinstr_o_19))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[18][29]~q ),
	.datac(\Reg[22][29]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux34~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~2 .lut_mask = 16'hAAE4;
defparam \Mux34~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N12
cycloneive_lcell_comb \Mux34~3 (
// Equation(s):
// \Mux34~3_combout  = (ifid_ifinstr_o_19 & ((\Mux34~2_combout  & (\Reg[30][29]~q )) # (!\Mux34~2_combout  & ((\Reg[26][29]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux34~2_combout ))))

	.dataa(\Reg[30][29]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[26][29]~q ),
	.datad(\Mux34~2_combout ),
	.cin(gnd),
	.combout(\Mux34~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~3 .lut_mask = 16'hBBC0;
defparam \Mux34~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N23
dffeas \Reg[16][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][29] .is_wysiwyg = "true";
defparam \Reg[16][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N22
cycloneive_lcell_comb \Mux34~4 (
// Equation(s):
// \Mux34~4_combout  = (ifid_ifinstr_o_19 & (((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[20][29]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[16][29]~q )))))

	.dataa(\Reg[20][29]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[16][29]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux34~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~4 .lut_mask = 16'hEE30;
defparam \Mux34~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N6
cycloneive_lcell_comb \Mux34~5 (
// Equation(s):
// \Mux34~5_combout  = (ifid_ifinstr_o_19 & ((\Mux34~4_combout  & (\Reg[28][29]~q )) # (!\Mux34~4_combout  & ((\Reg[24][29]~q ))))) # (!ifid_ifinstr_o_19 & (\Mux34~4_combout ))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Mux34~4_combout ),
	.datac(\Reg[28][29]~q ),
	.datad(\Reg[24][29]~q ),
	.cin(gnd),
	.combout(\Mux34~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~5 .lut_mask = 16'hE6C4;
defparam \Mux34~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N24
cycloneive_lcell_comb \Mux34~6 (
// Equation(s):
// \Mux34~6_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Mux34~3_combout )) # (!ifid_ifinstr_o_17 & ((\Mux34~5_combout )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux34~3_combout ),
	.datad(\Mux34~5_combout ),
	.cin(gnd),
	.combout(\Mux34~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~6 .lut_mask = 16'hD9C8;
defparam \Mux34~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N0
cycloneive_lcell_comb \Mux34~10 (
// Equation(s):
// \Mux34~10_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[5][29]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[4][29]~q ))))

	.dataa(\Reg[4][29]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[5][29]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux34~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~10 .lut_mask = 16'hFC22;
defparam \Mux34~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N26
cycloneive_lcell_comb \Mux34~11 (
// Equation(s):
// \Mux34~11_combout  = (\Mux34~10_combout  & ((\Reg[7][29]~q ) # ((!ifid_ifinstr_o_17)))) # (!\Mux34~10_combout  & (((\Reg[6][29]~q  & ifid_ifinstr_o_17))))

	.dataa(\Mux34~10_combout ),
	.datab(\Reg[7][29]~q ),
	.datac(\Reg[6][29]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux34~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~11 .lut_mask = 16'hD8AA;
defparam \Mux34~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N23
dffeas \Reg[1][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat18),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][29] .is_wysiwyg = "true";
defparam \Reg[1][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N22
cycloneive_lcell_comb \Mux34~14 (
// Equation(s):
// \Mux34~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][29]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][29]~q )))))

	.dataa(\Reg[3][29]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[1][29]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux34~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~14 .lut_mask = 16'hB800;
defparam \Mux34~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N14
cycloneive_lcell_comb \Mux34~15 (
// Equation(s):
// \Mux34~15_combout  = (\Mux34~14_combout ) # ((!ifid_ifinstr_o_16 & (\Reg[2][29]~q  & ifid_ifinstr_o_17)))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux34~14_combout ),
	.datac(\Reg[2][29]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux34~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~15 .lut_mask = 16'hDCCC;
defparam \Mux34~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N2
cycloneive_lcell_comb \Mux34~12 (
// Equation(s):
// \Mux34~12_combout  = (ifid_ifinstr_o_17 & ((\Reg[10][29]~q ) # ((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & (((\Reg[8][29]~q  & !ifid_ifinstr_o_16))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[10][29]~q ),
	.datac(\Reg[8][29]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux34~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~12 .lut_mask = 16'hAAD8;
defparam \Mux34~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N22
cycloneive_lcell_comb \Mux34~13 (
// Equation(s):
// \Mux34~13_combout  = (ifid_ifinstr_o_16 & ((\Mux34~12_combout  & ((\Reg[11][29]~q ))) # (!\Mux34~12_combout  & (\Reg[9][29]~q )))) # (!ifid_ifinstr_o_16 & (((\Mux34~12_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[9][29]~q ),
	.datac(\Reg[11][29]~q ),
	.datad(\Mux34~12_combout ),
	.cin(gnd),
	.combout(\Mux34~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~13 .lut_mask = 16'hF588;
defparam \Mux34~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N8
cycloneive_lcell_comb \Mux34~16 (
// Equation(s):
// \Mux34~16_combout  = (ifid_ifinstr_o_19 & (((ifid_ifinstr_o_18) # (\Mux34~13_combout )))) # (!ifid_ifinstr_o_19 & (\Mux34~15_combout  & (!ifid_ifinstr_o_18)))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Mux34~15_combout ),
	.datac(ifid_ifinstr_o_18),
	.datad(\Mux34~13_combout ),
	.cin(gnd),
	.combout(\Mux34~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~16 .lut_mask = 16'hAEA4;
defparam \Mux34~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N2
cycloneive_lcell_comb \Mux34~17 (
// Equation(s):
// \Mux34~17_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[13][29]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[12][29]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[13][29]~q ),
	.datac(\Reg[12][29]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux34~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~17 .lut_mask = 16'hEE50;
defparam \Mux34~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N22
cycloneive_lcell_comb \Mux34~18 (
// Equation(s):
// \Mux34~18_combout  = (\Mux34~17_combout  & (((\Reg[15][29]~q ) # (!ifid_ifinstr_o_17)))) # (!\Mux34~17_combout  & (\Reg[14][29]~q  & ((ifid_ifinstr_o_17))))

	.dataa(\Mux34~17_combout ),
	.datab(\Reg[14][29]~q ),
	.datac(\Reg[15][29]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux34~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~18 .lut_mask = 16'hE4AA;
defparam \Mux34~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N8
cycloneive_lcell_comb \Mux33~7 (
// Equation(s):
// \Mux33~7_combout  = (ifid_ifinstr_o_18 & (((\Reg[23][30]~q ) # (ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (\Reg[19][30]~q  & ((!ifid_ifinstr_o_19))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[19][30]~q ),
	.datac(\Reg[23][30]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux33~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~7 .lut_mask = 16'hAAE4;
defparam \Mux33~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N0
cycloneive_lcell_comb \Reg[27][30]~feeder (
// Equation(s):
// \Reg[27][30]~feeder_combout  = \wdat~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat19),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[27][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[27][30]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[27][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N1
dffeas \Reg[27][30] (
	.clk(!CLK),
	.d(\Reg[27][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[27][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[27][30] .is_wysiwyg = "true";
defparam \Reg[27][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N30
cycloneive_lcell_comb \Mux33~8 (
// Equation(s):
// \Mux33~8_combout  = (\Mux33~7_combout  & (((\Reg[31][30]~q ) # (!ifid_ifinstr_o_19)))) # (!\Mux33~7_combout  & (\Reg[27][30]~q  & ((ifid_ifinstr_o_19))))

	.dataa(\Mux33~7_combout ),
	.datab(\Reg[27][30]~q ),
	.datac(\Reg[31][30]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux33~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~8 .lut_mask = 16'hE4AA;
defparam \Mux33~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N4
cycloneive_lcell_comb \Mux33~5 (
// Equation(s):
// \Mux33~5_combout  = (\Mux33~4_combout  & (((\Reg[28][30]~q )) # (!ifid_ifinstr_o_18))) # (!\Mux33~4_combout  & (ifid_ifinstr_o_18 & (\Reg[20][30]~q )))

	.dataa(\Mux33~4_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[20][30]~q ),
	.datad(\Reg[28][30]~q ),
	.cin(gnd),
	.combout(\Mux33~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~5 .lut_mask = 16'hEA62;
defparam \Mux33~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N16
cycloneive_lcell_comb \Mux33~2 (
// Equation(s):
// \Mux33~2_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[26][30]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[18][30]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[18][30]~q ),
	.datad(\Reg[26][30]~q ),
	.cin(gnd),
	.combout(\Mux33~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~2 .lut_mask = 16'hDC98;
defparam \Mux33~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N30
cycloneive_lcell_comb \Mux33~3 (
// Equation(s):
// \Mux33~3_combout  = (ifid_ifinstr_o_18 & ((\Mux33~2_combout  & ((\Reg[30][30]~q ))) # (!\Mux33~2_combout  & (\Reg[22][30]~q )))) # (!ifid_ifinstr_o_18 & (((\Mux33~2_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[22][30]~q ),
	.datac(\Reg[30][30]~q ),
	.datad(\Mux33~2_combout ),
	.cin(gnd),
	.combout(\Mux33~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~3 .lut_mask = 16'hF588;
defparam \Mux33~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N30
cycloneive_lcell_comb \Mux33~6 (
// Equation(s):
// \Mux33~6_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Mux33~3_combout ))) # (!ifid_ifinstr_o_17 & (\Mux33~5_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux33~5_combout ),
	.datad(\Mux33~3_combout ),
	.cin(gnd),
	.combout(\Mux33~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~6 .lut_mask = 16'hDC98;
defparam \Mux33~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N4
cycloneive_lcell_comb \Mux33~0 (
// Equation(s):
// \Mux33~0_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[21][30]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[17][30]~q )))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[21][30]~q ),
	.datad(\Reg[17][30]~q ),
	.cin(gnd),
	.combout(\Mux33~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~0 .lut_mask = 16'hD9C8;
defparam \Mux33~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N14
cycloneive_lcell_comb \Mux33~1 (
// Equation(s):
// \Mux33~1_combout  = (\Mux33~0_combout  & ((\Reg[29][30]~q ) # ((!ifid_ifinstr_o_19)))) # (!\Mux33~0_combout  & (((\Reg[25][30]~q  & ifid_ifinstr_o_19))))

	.dataa(\Mux33~0_combout ),
	.datab(\Reg[29][30]~q ),
	.datac(\Reg[25][30]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux33~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~1 .lut_mask = 16'hD8AA;
defparam \Mux33~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N10
cycloneive_lcell_comb \Mux33~17 (
// Equation(s):
// \Mux33~17_combout  = (ifid_ifinstr_o_16 & (((\Reg[13][30]~q ) # (ifid_ifinstr_o_17)))) # (!ifid_ifinstr_o_16 & (\Reg[12][30]~q  & ((!ifid_ifinstr_o_17))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[12][30]~q ),
	.datac(\Reg[13][30]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux33~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~17 .lut_mask = 16'hAAE4;
defparam \Mux33~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N26
cycloneive_lcell_comb \Mux33~18 (
// Equation(s):
// \Mux33~18_combout  = (\Mux33~17_combout  & (((\Reg[15][30]~q ) # (!ifid_ifinstr_o_17)))) # (!\Mux33~17_combout  & (\Reg[14][30]~q  & ((ifid_ifinstr_o_17))))

	.dataa(\Mux33~17_combout ),
	.datab(\Reg[14][30]~q ),
	.datac(\Reg[15][30]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux33~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~18 .lut_mask = 16'hE4AA;
defparam \Mux33~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y36_N15
dffeas \Reg[8][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][30] .is_wysiwyg = "true";
defparam \Reg[8][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y36_N1
dffeas \Reg[10][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[10][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[10][30] .is_wysiwyg = "true";
defparam \Reg[10][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N0
cycloneive_lcell_comb \Mux33~10 (
// Equation(s):
// \Mux33~10_combout  = (ifid_ifinstr_o_16 & (((ifid_ifinstr_o_17)))) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[10][30]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[8][30]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[8][30]~q ),
	.datac(\Reg[10][30]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux33~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~10 .lut_mask = 16'hFA44;
defparam \Mux33~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N20
cycloneive_lcell_comb \Mux33~11 (
// Equation(s):
// \Mux33~11_combout  = (ifid_ifinstr_o_16 & ((\Mux33~10_combout  & ((\Reg[11][30]~q ))) # (!\Mux33~10_combout  & (\Reg[9][30]~q )))) # (!ifid_ifinstr_o_16 & (\Mux33~10_combout ))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Mux33~10_combout ),
	.datac(\Reg[9][30]~q ),
	.datad(\Reg[11][30]~q ),
	.cin(gnd),
	.combout(\Mux33~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~11 .lut_mask = 16'hEC64;
defparam \Mux33~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N13
dffeas \Reg[1][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat19),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][30] .is_wysiwyg = "true";
defparam \Reg[1][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N12
cycloneive_lcell_comb \Mux33~14 (
// Equation(s):
// \Mux33~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][30]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][30]~q )))))

	.dataa(\Reg[3][30]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[1][30]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux33~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~14 .lut_mask = 16'hB800;
defparam \Mux33~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N20
cycloneive_lcell_comb \Mux33~15 (
// Equation(s):
// \Mux33~15_combout  = (\Mux33~14_combout ) # ((\Reg[2][30]~q  & (ifid_ifinstr_o_17 & !ifid_ifinstr_o_16)))

	.dataa(\Reg[2][30]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux33~14_combout ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux33~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~15 .lut_mask = 16'hF0F8;
defparam \Mux33~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N16
cycloneive_lcell_comb \Mux33~13 (
// Equation(s):
// \Mux33~13_combout  = (\Mux33~12_combout  & (((\Reg[7][30]~q ) # (!ifid_ifinstr_o_17)))) # (!\Mux33~12_combout  & (\Reg[6][30]~q  & ((ifid_ifinstr_o_17))))

	.dataa(\Mux33~12_combout ),
	.datab(\Reg[6][30]~q ),
	.datac(\Reg[7][30]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux33~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~13 .lut_mask = 16'hE4AA;
defparam \Mux33~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N10
cycloneive_lcell_comb \Mux33~16 (
// Equation(s):
// \Mux33~16_combout  = (ifid_ifinstr_o_19 & (((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Mux33~13_combout ))) # (!ifid_ifinstr_o_18 & (\Mux33~15_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Mux33~15_combout ),
	.datac(ifid_ifinstr_o_18),
	.datad(\Mux33~13_combout ),
	.cin(gnd),
	.combout(\Mux33~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~16 .lut_mask = 16'hF4A4;
defparam \Mux33~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N22
cycloneive_lcell_comb \Mux54~7 (
// Equation(s):
// \Mux54~7_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[27][9]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[19][9]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[19][9]~q ),
	.datad(\Reg[27][9]~q ),
	.cin(gnd),
	.combout(\Mux54~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~7 .lut_mask = 16'hDC98;
defparam \Mux54~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N16
cycloneive_lcell_comb \Mux54~8 (
// Equation(s):
// \Mux54~8_combout  = (\Mux54~7_combout  & ((\Reg[31][9]~q ) # ((!ifid_ifinstr_o_18)))) # (!\Mux54~7_combout  & (((\Reg[23][9]~q  & ifid_ifinstr_o_18))))

	.dataa(\Mux54~7_combout ),
	.datab(\Reg[31][9]~q ),
	.datac(\Reg[23][9]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux54~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~8 .lut_mask = 16'hD8AA;
defparam \Mux54~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N28
cycloneive_lcell_comb \Mux54~0 (
// Equation(s):
// \Mux54~0_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[25][9]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[17][9]~q ))))

	.dataa(\Reg[17][9]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[25][9]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux54~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~0 .lut_mask = 16'hFC22;
defparam \Mux54~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N8
cycloneive_lcell_comb \Mux54~1 (
// Equation(s):
// \Mux54~1_combout  = (ifid_ifinstr_o_18 & ((\Mux54~0_combout  & (\Reg[29][9]~q )) # (!\Mux54~0_combout  & ((\Reg[21][9]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux54~0_combout ))))

	.dataa(\Reg[29][9]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[21][9]~q ),
	.datad(\Mux54~0_combout ),
	.cin(gnd),
	.combout(\Mux54~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~1 .lut_mask = 16'hBBC0;
defparam \Mux54~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N19
dffeas \Reg[16][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][9] .is_wysiwyg = "true";
defparam \Reg[16][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N18
cycloneive_lcell_comb \Mux54~4 (
// Equation(s):
// \Mux54~4_combout  = (ifid_ifinstr_o_19 & (((ifid_ifinstr_o_18)))) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[20][9]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[16][9]~q )))))

	.dataa(\Reg[20][9]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[16][9]~q ),
	.datad(ifid_ifinstr_o_18),
	.cin(gnd),
	.combout(\Mux54~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~4 .lut_mask = 16'hEE30;
defparam \Mux54~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N15
dffeas \Reg[28][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][9] .is_wysiwyg = "true";
defparam \Reg[28][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N14
cycloneive_lcell_comb \Mux54~5 (
// Equation(s):
// \Mux54~5_combout  = (\Mux54~4_combout  & (((\Reg[28][9]~q ) # (!ifid_ifinstr_o_19)))) # (!\Mux54~4_combout  & (\Reg[24][9]~q  & ((ifid_ifinstr_o_19))))

	.dataa(\Reg[24][9]~q ),
	.datab(\Mux54~4_combout ),
	.datac(\Reg[28][9]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux54~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~5 .lut_mask = 16'hE2CC;
defparam \Mux54~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N29
dffeas \Reg[22][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][9] .is_wysiwyg = "true";
defparam \Reg[22][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N28
cycloneive_lcell_comb \Mux54~2 (
// Equation(s):
// \Mux54~2_combout  = (ifid_ifinstr_o_18 & (((\Reg[22][9]~q ) # (ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (\Reg[18][9]~q  & ((!ifid_ifinstr_o_19))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[18][9]~q ),
	.datac(\Reg[22][9]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux54~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~2 .lut_mask = 16'hAAE4;
defparam \Mux54~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N8
cycloneive_lcell_comb \Mux54~3 (
// Equation(s):
// \Mux54~3_combout  = (ifid_ifinstr_o_19 & ((\Mux54~2_combout  & ((\Reg[30][9]~q ))) # (!\Mux54~2_combout  & (\Reg[26][9]~q )))) # (!ifid_ifinstr_o_19 & (((\Mux54~2_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[26][9]~q ),
	.datac(\Reg[30][9]~q ),
	.datad(\Mux54~2_combout ),
	.cin(gnd),
	.combout(\Mux54~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~3 .lut_mask = 16'hF588;
defparam \Mux54~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N28
cycloneive_lcell_comb \Mux54~6 (
// Equation(s):
// \Mux54~6_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Mux54~3_combout ))) # (!ifid_ifinstr_o_17 & (\Mux54~5_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux54~5_combout ),
	.datad(\Mux54~3_combout ),
	.cin(gnd),
	.combout(\Mux54~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~6 .lut_mask = 16'hDC98;
defparam \Mux54~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N28
cycloneive_lcell_comb \Mux54~10 (
// Equation(s):
// \Mux54~10_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[5][9]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[4][9]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[5][9]~q ),
	.datad(\Reg[4][9]~q ),
	.cin(gnd),
	.combout(\Mux54~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~10 .lut_mask = 16'hD9C8;
defparam \Mux54~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N4
cycloneive_lcell_comb \Mux54~11 (
// Equation(s):
// \Mux54~11_combout  = (ifid_ifinstr_o_17 & ((\Mux54~10_combout  & (\Reg[7][9]~q )) # (!\Mux54~10_combout  & ((\Reg[6][9]~q ))))) # (!ifid_ifinstr_o_17 & (((\Mux54~10_combout ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[7][9]~q ),
	.datac(\Reg[6][9]~q ),
	.datad(\Mux54~10_combout ),
	.cin(gnd),
	.combout(\Mux54~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~11 .lut_mask = 16'hDDA0;
defparam \Mux54~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N20
cycloneive_lcell_comb \Mux54~17 (
// Equation(s):
// \Mux54~17_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[13][9]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[12][9]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[12][9]~q ),
	.datac(\Reg[13][9]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux54~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~17 .lut_mask = 16'hFA44;
defparam \Mux54~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N2
cycloneive_lcell_comb \Mux54~18 (
// Equation(s):
// \Mux54~18_combout  = (ifid_ifinstr_o_17 & ((\Mux54~17_combout  & (\Reg[15][9]~q )) # (!\Mux54~17_combout  & ((\Reg[14][9]~q ))))) # (!ifid_ifinstr_o_17 & (((\Mux54~17_combout ))))

	.dataa(\Reg[15][9]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[14][9]~q ),
	.datad(\Mux54~17_combout ),
	.cin(gnd),
	.combout(\Mux54~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~18 .lut_mask = 16'hBBC0;
defparam \Mux54~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y36_N1
dffeas \Reg[1][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat16),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[1][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[1][9] .is_wysiwyg = "true";
defparam \Reg[1][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N0
cycloneive_lcell_comb \Mux54~14 (
// Equation(s):
// \Mux54~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][9]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][9]~q )))))

	.dataa(\Reg[3][9]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[1][9]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux54~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~14 .lut_mask = 16'hB800;
defparam \Mux54~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N2
cycloneive_lcell_comb \Mux54~15 (
// Equation(s):
// \Mux54~15_combout  = (\Mux54~14_combout ) # ((!ifid_ifinstr_o_16 & (\Reg[2][9]~q  & ifid_ifinstr_o_17)))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[2][9]~q ),
	.datac(\Mux54~14_combout ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux54~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~15 .lut_mask = 16'hF4F0;
defparam \Mux54~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N10
cycloneive_lcell_comb \Mux54~12 (
// Equation(s):
// \Mux54~12_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[10][9]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[8][9]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[8][9]~q ),
	.datad(\Reg[10][9]~q ),
	.cin(gnd),
	.combout(\Mux54~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~12 .lut_mask = 16'hDC98;
defparam \Mux54~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N6
cycloneive_lcell_comb \Mux54~13 (
// Equation(s):
// \Mux54~13_combout  = (ifid_ifinstr_o_16 & ((\Mux54~12_combout  & ((\Reg[11][9]~q ))) # (!\Mux54~12_combout  & (\Reg[9][9]~q )))) # (!ifid_ifinstr_o_16 & (((\Mux54~12_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[9][9]~q ),
	.datac(\Reg[11][9]~q ),
	.datad(\Mux54~12_combout ),
	.cin(gnd),
	.combout(\Mux54~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~13 .lut_mask = 16'hF588;
defparam \Mux54~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N0
cycloneive_lcell_comb \Mux54~16 (
// Equation(s):
// \Mux54~16_combout  = (ifid_ifinstr_o_19 & (((ifid_ifinstr_o_18) # (\Mux54~13_combout )))) # (!ifid_ifinstr_o_19 & (\Mux54~15_combout  & (!ifid_ifinstr_o_18)))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Mux54~15_combout ),
	.datac(ifid_ifinstr_o_18),
	.datad(\Mux54~13_combout ),
	.cin(gnd),
	.combout(\Mux54~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~16 .lut_mask = 16'hAEA4;
defparam \Mux54~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N28
cycloneive_lcell_comb \Mux49~7 (
// Equation(s):
// \Mux49~7_combout  = (ifid_ifinstr_o_18 & (((\Reg[23][14]~q ) # (ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (\Reg[19][14]~q  & ((!ifid_ifinstr_o_19))))

	.dataa(\Reg[19][14]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[23][14]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux49~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~7 .lut_mask = 16'hCCE2;
defparam \Mux49~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N30
cycloneive_lcell_comb \Mux49~8 (
// Equation(s):
// \Mux49~8_combout  = (ifid_ifinstr_o_19 & ((\Mux49~7_combout  & ((\Reg[31][14]~q ))) # (!\Mux49~7_combout  & (\Reg[27][14]~q )))) # (!ifid_ifinstr_o_19 & (((\Mux49~7_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[27][14]~q ),
	.datac(\Reg[31][14]~q ),
	.datad(\Mux49~7_combout ),
	.cin(gnd),
	.combout(\Mux49~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~8 .lut_mask = 16'hF588;
defparam \Mux49~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N2
cycloneive_lcell_comb \Mux49~0 (
// Equation(s):
// \Mux49~0_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Reg[21][14]~q ))) # (!ifid_ifinstr_o_18 & (\Reg[17][14]~q ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[17][14]~q ),
	.datad(\Reg[21][14]~q ),
	.cin(gnd),
	.combout(\Mux49~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~0 .lut_mask = 16'hDC98;
defparam \Mux49~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N12
cycloneive_lcell_comb \Mux49~1 (
// Equation(s):
// \Mux49~1_combout  = (\Mux49~0_combout  & (((\Reg[29][14]~q ) # (!ifid_ifinstr_o_19)))) # (!\Mux49~0_combout  & (\Reg[25][14]~q  & ((ifid_ifinstr_o_19))))

	.dataa(\Reg[25][14]~q ),
	.datab(\Mux49~0_combout ),
	.datac(\Reg[29][14]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux49~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~1 .lut_mask = 16'hE2CC;
defparam \Mux49~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N15
dffeas \Reg[16][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][14] .is_wysiwyg = "true";
defparam \Reg[16][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N14
cycloneive_lcell_comb \Mux49~4 (
// Equation(s):
// \Mux49~4_combout  = (ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18) # ((\Reg[24][14]~q )))) # (!ifid_ifinstr_o_19 & (!ifid_ifinstr_o_18 & (\Reg[16][14]~q )))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[16][14]~q ),
	.datad(\Reg[24][14]~q ),
	.cin(gnd),
	.combout(\Mux49~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~4 .lut_mask = 16'hBA98;
defparam \Mux49~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y34_N17
dffeas \Reg[20][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat11),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~11_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[20][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[20][14] .is_wysiwyg = "true";
defparam \Reg[20][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N10
cycloneive_lcell_comb \Mux49~5 (
// Equation(s):
// \Mux49~5_combout  = (\Mux49~4_combout  & ((\Reg[28][14]~q ) # ((!ifid_ifinstr_o_18)))) # (!\Mux49~4_combout  & (((ifid_ifinstr_o_18 & \Reg[20][14]~q ))))

	.dataa(\Reg[28][14]~q ),
	.datab(\Mux49~4_combout ),
	.datac(ifid_ifinstr_o_18),
	.datad(\Reg[20][14]~q ),
	.cin(gnd),
	.combout(\Mux49~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~5 .lut_mask = 16'hBC8C;
defparam \Mux49~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N0
cycloneive_lcell_comb \Mux49~2 (
// Equation(s):
// \Mux49~2_combout  = (ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18) # ((\Reg[26][14]~q )))) # (!ifid_ifinstr_o_19 & (!ifid_ifinstr_o_18 & ((\Reg[18][14]~q ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[26][14]~q ),
	.datad(\Reg[18][14]~q ),
	.cin(gnd),
	.combout(\Mux49~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~2 .lut_mask = 16'hB9A8;
defparam \Mux49~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N26
cycloneive_lcell_comb \Mux49~3 (
// Equation(s):
// \Mux49~3_combout  = (ifid_ifinstr_o_18 & ((\Mux49~2_combout  & (\Reg[30][14]~q )) # (!\Mux49~2_combout  & ((\Reg[22][14]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux49~2_combout ))))

	.dataa(\Reg[30][14]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Mux49~2_combout ),
	.datad(\Reg[22][14]~q ),
	.cin(gnd),
	.combout(\Mux49~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~3 .lut_mask = 16'hBCB0;
defparam \Mux49~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N6
cycloneive_lcell_comb \Mux49~6 (
// Equation(s):
// \Mux49~6_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16) # (\Mux49~3_combout )))) # (!ifid_ifinstr_o_17 & (\Mux49~5_combout  & (!ifid_ifinstr_o_16)))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux49~5_combout ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux49~3_combout ),
	.cin(gnd),
	.combout(\Mux49~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~6 .lut_mask = 16'hAEA4;
defparam \Mux49~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N10
cycloneive_lcell_comb \Mux49~14 (
// Equation(s):
// \Mux49~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[3][14]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[1][14]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[1][14]~q ),
	.datad(\Reg[3][14]~q ),
	.cin(gnd),
	.combout(\Mux49~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~14 .lut_mask = 16'hA820;
defparam \Mux49~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N10
cycloneive_lcell_comb \Mux49~15 (
// Equation(s):
// \Mux49~15_combout  = (\Mux49~14_combout ) # ((ifid_ifinstr_o_17 & (\Reg[2][14]~q  & !ifid_ifinstr_o_16)))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[2][14]~q ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux49~14_combout ),
	.cin(gnd),
	.combout(\Mux49~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~15 .lut_mask = 16'hFF08;
defparam \Mux49~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N30
cycloneive_lcell_comb \Mux49~13 (
// Equation(s):
// \Mux49~13_combout  = (\Mux49~12_combout  & (((\Reg[7][14]~q )) # (!ifid_ifinstr_o_17))) # (!\Mux49~12_combout  & (ifid_ifinstr_o_17 & ((\Reg[6][14]~q ))))

	.dataa(\Mux49~12_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[7][14]~q ),
	.datad(\Reg[6][14]~q ),
	.cin(gnd),
	.combout(\Mux49~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~13 .lut_mask = 16'hE6A2;
defparam \Mux49~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N12
cycloneive_lcell_comb \Mux49~16 (
// Equation(s):
// \Mux49~16_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19) # (\Mux49~13_combout )))) # (!ifid_ifinstr_o_18 & (\Mux49~15_combout  & (!ifid_ifinstr_o_19)))

	.dataa(\Mux49~15_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux49~13_combout ),
	.cin(gnd),
	.combout(\Mux49~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~16 .lut_mask = 16'hCEC2;
defparam \Mux49~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N24
cycloneive_lcell_comb \Mux49~10 (
// Equation(s):
// \Mux49~10_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[10][14]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[8][14]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[10][14]~q ),
	.datad(\Reg[8][14]~q ),
	.cin(gnd),
	.combout(\Mux49~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~10 .lut_mask = 16'hD9C8;
defparam \Mux49~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N20
cycloneive_lcell_comb \Mux49~11 (
// Equation(s):
// \Mux49~11_combout  = (ifid_ifinstr_o_16 & ((\Mux49~10_combout  & (\Reg[11][14]~q )) # (!\Mux49~10_combout  & ((\Reg[9][14]~q ))))) # (!ifid_ifinstr_o_16 & (((\Mux49~10_combout ))))

	.dataa(\Reg[11][14]~q ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[9][14]~q ),
	.datad(\Mux49~10_combout ),
	.cin(gnd),
	.combout(\Mux49~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~11 .lut_mask = 16'hBBC0;
defparam \Mux49~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N16
cycloneive_lcell_comb \Mux49~17 (
// Equation(s):
// \Mux49~17_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[13][14]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[12][14]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[13][14]~q ),
	.datad(\Reg[12][14]~q ),
	.cin(gnd),
	.combout(\Mux49~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~17 .lut_mask = 16'hD9C8;
defparam \Mux49~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N18
cycloneive_lcell_comb \Mux49~18 (
// Equation(s):
// \Mux49~18_combout  = (\Mux49~17_combout  & ((\Reg[15][14]~q ) # ((!ifid_ifinstr_o_17)))) # (!\Mux49~17_combout  & (((\Reg[14][14]~q  & ifid_ifinstr_o_17))))

	.dataa(\Reg[15][14]~q ),
	.datab(\Reg[14][14]~q ),
	.datac(\Mux49~17_combout ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux49~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~18 .lut_mask = 16'hACF0;
defparam \Mux49~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N28
cycloneive_lcell_comb \Mux48~7 (
// Equation(s):
// \Mux48~7_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Reg[27][15]~q )) # (!ifid_ifinstr_o_19 & ((\Reg[19][15]~q )))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[27][15]~q ),
	.datad(\Reg[19][15]~q ),
	.cin(gnd),
	.combout(\Mux48~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~7 .lut_mask = 16'hD9C8;
defparam \Mux48~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N18
cycloneive_lcell_comb \Mux48~8 (
// Equation(s):
// \Mux48~8_combout  = (ifid_ifinstr_o_18 & ((\Mux48~7_combout  & (\Reg[31][15]~q )) # (!\Mux48~7_combout  & ((\Reg[23][15]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux48~7_combout ))))

	.dataa(\Reg[31][15]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[23][15]~q ),
	.datad(\Mux48~7_combout ),
	.cin(gnd),
	.combout(\Mux48~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~8 .lut_mask = 16'hBBC0;
defparam \Mux48~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N18
cycloneive_lcell_comb \Mux48~0 (
// Equation(s):
// \Mux48~0_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[25][15]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[17][15]~q ))))

	.dataa(\Reg[17][15]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(ifid_ifinstr_o_19),
	.datad(\Reg[25][15]~q ),
	.cin(gnd),
	.combout(\Mux48~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~0 .lut_mask = 16'hF2C2;
defparam \Mux48~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y37_N24
cycloneive_lcell_comb \Mux48~1 (
// Equation(s):
// \Mux48~1_combout  = (ifid_ifinstr_o_18 & ((\Mux48~0_combout  & (\Reg[29][15]~q )) # (!\Mux48~0_combout  & ((\Reg[21][15]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux48~0_combout ))))

	.dataa(\Reg[29][15]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[21][15]~q ),
	.datad(\Mux48~0_combout ),
	.cin(gnd),
	.combout(\Mux48~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~1 .lut_mask = 16'hBBC0;
defparam \Mux48~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y33_N22
cycloneive_lcell_comb \Mux48~4 (
// Equation(s):
// \Mux48~4_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[20][15]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[16][15]~q )))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[20][15]~q ),
	.datad(\Reg[16][15]~q ),
	.cin(gnd),
	.combout(\Mux48~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~4 .lut_mask = 16'hD9C8;
defparam \Mux48~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N20
cycloneive_lcell_comb \Mux48~5 (
// Equation(s):
// \Mux48~5_combout  = (ifid_ifinstr_o_19 & ((\Mux48~4_combout  & (\Reg[28][15]~q )) # (!\Mux48~4_combout  & ((\Reg[24][15]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux48~4_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[28][15]~q ),
	.datac(\Reg[24][15]~q ),
	.datad(\Mux48~4_combout ),
	.cin(gnd),
	.combout(\Mux48~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~5 .lut_mask = 16'hDDA0;
defparam \Mux48~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N7
dffeas \Reg[18][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][15] .is_wysiwyg = "true";
defparam \Reg[18][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N6
cycloneive_lcell_comb \Mux48~2 (
// Equation(s):
// \Mux48~2_combout  = (ifid_ifinstr_o_18 & ((\Reg[22][15]~q ) # ((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (((\Reg[18][15]~q  & !ifid_ifinstr_o_19))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[22][15]~q ),
	.datac(\Reg[18][15]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux48~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~2 .lut_mask = 16'hAAD8;
defparam \Mux48~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N24
cycloneive_lcell_comb \Mux48~3 (
// Equation(s):
// \Mux48~3_combout  = (ifid_ifinstr_o_19 & ((\Mux48~2_combout  & (\Reg[30][15]~q )) # (!\Mux48~2_combout  & ((\Reg[26][15]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux48~2_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[30][15]~q ),
	.datac(\Reg[26][15]~q ),
	.datad(\Mux48~2_combout ),
	.cin(gnd),
	.combout(\Mux48~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~3 .lut_mask = 16'hDDA0;
defparam \Mux48~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N18
cycloneive_lcell_comb \Mux48~6 (
// Equation(s):
// \Mux48~6_combout  = (ifid_ifinstr_o_16 & (((ifid_ifinstr_o_17)))) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Mux48~3_combout ))) # (!ifid_ifinstr_o_17 & (\Mux48~5_combout ))))

	.dataa(\Mux48~5_combout ),
	.datab(\Mux48~3_combout ),
	.datac(ifid_ifinstr_o_16),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux48~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~6 .lut_mask = 16'hFC0A;
defparam \Mux48~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y35_N30
cycloneive_lcell_comb \Mux48~13 (
// Equation(s):
// \Mux48~13_combout  = (\Mux48~12_combout  & ((\Reg[11][15]~q ) # ((!ifid_ifinstr_o_16)))) # (!\Mux48~12_combout  & (((\Reg[9][15]~q  & ifid_ifinstr_o_16))))

	.dataa(\Mux48~12_combout ),
	.datab(\Reg[11][15]~q ),
	.datac(\Reg[9][15]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux48~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~13 .lut_mask = 16'hD8AA;
defparam \Mux48~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N18
cycloneive_lcell_comb \Mux48~14 (
// Equation(s):
// \Mux48~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[3][15]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[1][15]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[1][15]~q ),
	.datad(\Reg[3][15]~q ),
	.cin(gnd),
	.combout(\Mux48~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~14 .lut_mask = 16'hA820;
defparam \Mux48~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N24
cycloneive_lcell_comb \Mux48~15 (
// Equation(s):
// \Mux48~15_combout  = (\Mux48~14_combout ) # ((ifid_ifinstr_o_17 & (\Reg[2][15]~q  & !ifid_ifinstr_o_16)))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux48~14_combout ),
	.datac(\Reg[2][15]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux48~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~15 .lut_mask = 16'hCCEC;
defparam \Mux48~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N10
cycloneive_lcell_comb \Mux48~16 (
// Equation(s):
// \Mux48~16_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Mux48~13_combout )) # (!ifid_ifinstr_o_19 & ((\Mux48~15_combout )))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux48~13_combout ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux48~15_combout ),
	.cin(gnd),
	.combout(\Mux48~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~16 .lut_mask = 16'hE5E0;
defparam \Mux48~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N8
cycloneive_lcell_comb \Mux48~17 (
// Equation(s):
// \Mux48~17_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[13][15]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[12][15]~q )))))

	.dataa(\Reg[13][15]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[12][15]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux48~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~17 .lut_mask = 16'hEE30;
defparam \Mux48~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N18
cycloneive_lcell_comb \Mux48~18 (
// Equation(s):
// \Mux48~18_combout  = (ifid_ifinstr_o_17 & ((\Mux48~17_combout  & ((\Reg[15][15]~q ))) # (!\Mux48~17_combout  & (\Reg[14][15]~q )))) # (!ifid_ifinstr_o_17 & (((\Mux48~17_combout ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[14][15]~q ),
	.datac(\Reg[15][15]~q ),
	.datad(\Mux48~17_combout ),
	.cin(gnd),
	.combout(\Mux48~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~18 .lut_mask = 16'hF588;
defparam \Mux48~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y39_N13
dffeas \Reg[5][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][15] .is_wysiwyg = "true";
defparam \Reg[5][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y39_N19
dffeas \Reg[4][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat10),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][15] .is_wysiwyg = "true";
defparam \Reg[4][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N12
cycloneive_lcell_comb \Mux48~10 (
// Equation(s):
// \Mux48~10_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[5][15]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[4][15]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[5][15]~q ),
	.datad(\Reg[4][15]~q ),
	.cin(gnd),
	.combout(\Mux48~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~10 .lut_mask = 16'hD9C8;
defparam \Mux48~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N4
cycloneive_lcell_comb \Mux48~11 (
// Equation(s):
// \Mux48~11_combout  = (\Mux48~10_combout  & ((\Reg[7][15]~q ) # ((!ifid_ifinstr_o_17)))) # (!\Mux48~10_combout  & (((\Reg[6][15]~q  & ifid_ifinstr_o_17))))

	.dataa(\Mux48~10_combout ),
	.datab(\Reg[7][15]~q ),
	.datac(\Reg[6][15]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux48~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~11 .lut_mask = 16'hD8AA;
defparam \Mux48~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N10
cycloneive_lcell_comb \Mux53~7 (
// Equation(s):
// \Mux53~7_combout  = (ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19) # ((\Reg[23][10]~q )))) # (!ifid_ifinstr_o_18 & (!ifid_ifinstr_o_19 & (\Reg[19][10]~q )))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[19][10]~q ),
	.datad(\Reg[23][10]~q ),
	.cin(gnd),
	.combout(\Mux53~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~7 .lut_mask = 16'hBA98;
defparam \Mux53~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N8
cycloneive_lcell_comb \Mux53~8 (
// Equation(s):
// \Mux53~8_combout  = (\Mux53~7_combout  & (((\Reg[31][10]~q )) # (!ifid_ifinstr_o_19))) # (!\Mux53~7_combout  & (ifid_ifinstr_o_19 & ((\Reg[27][10]~q ))))

	.dataa(\Mux53~7_combout ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[31][10]~q ),
	.datad(\Reg[27][10]~q ),
	.cin(gnd),
	.combout(\Mux53~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~8 .lut_mask = 16'hE6A2;
defparam \Mux53~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N2
cycloneive_lcell_comb \Mux53~4 (
// Equation(s):
// \Mux53~4_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[24][10]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[16][10]~q ))))

	.dataa(\Reg[16][10]~q ),
	.datab(\Reg[24][10]~q ),
	.datac(ifid_ifinstr_o_18),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux53~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~4 .lut_mask = 16'hFC0A;
defparam \Mux53~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N30
cycloneive_lcell_comb \Mux53~5 (
// Equation(s):
// \Mux53~5_combout  = (ifid_ifinstr_o_18 & ((\Mux53~4_combout  & (\Reg[28][10]~q )) # (!\Mux53~4_combout  & ((\Reg[20][10]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux53~4_combout ))))

	.dataa(\Reg[28][10]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[20][10]~q ),
	.datad(\Mux53~4_combout ),
	.cin(gnd),
	.combout(\Mux53~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~5 .lut_mask = 16'hBBC0;
defparam \Mux53~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y36_N19
dffeas \Reg[30][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~9_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[30][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[30][10] .is_wysiwyg = "true";
defparam \Reg[30][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N18
cycloneive_lcell_comb \Mux53~3 (
// Equation(s):
// \Mux53~3_combout  = (\Mux53~2_combout  & (((\Reg[30][10]~q )) # (!ifid_ifinstr_o_18))) # (!\Mux53~2_combout  & (ifid_ifinstr_o_18 & ((\Reg[22][10]~q ))))

	.dataa(\Mux53~2_combout ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[30][10]~q ),
	.datad(\Reg[22][10]~q ),
	.cin(gnd),
	.combout(\Mux53~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~3 .lut_mask = 16'hE6A2;
defparam \Mux53~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N28
cycloneive_lcell_comb \Mux53~6 (
// Equation(s):
// \Mux53~6_combout  = (ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16) # ((\Mux53~3_combout )))) # (!ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & (\Mux53~5_combout )))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux53~5_combout ),
	.datad(\Mux53~3_combout ),
	.cin(gnd),
	.combout(\Mux53~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~6 .lut_mask = 16'hBA98;
defparam \Mux53~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N24
cycloneive_lcell_comb \Mux53~0 (
// Equation(s):
// \Mux53~0_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Reg[21][10]~q ))) # (!ifid_ifinstr_o_18 & (\Reg[17][10]~q ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[17][10]~q ),
	.datad(\Reg[21][10]~q ),
	.cin(gnd),
	.combout(\Mux53~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~0 .lut_mask = 16'hDC98;
defparam \Mux53~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N10
cycloneive_lcell_comb \Mux53~1 (
// Equation(s):
// \Mux53~1_combout  = (ifid_ifinstr_o_19 & ((\Mux53~0_combout  & (\Reg[29][10]~q )) # (!\Mux53~0_combout  & ((\Reg[25][10]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux53~0_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[29][10]~q ),
	.datac(\Mux53~0_combout ),
	.datad(\Reg[25][10]~q ),
	.cin(gnd),
	.combout(\Mux53~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~1 .lut_mask = 16'hDAD0;
defparam \Mux53~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N31
dffeas \Reg[12][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat15),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][10] .is_wysiwyg = "true";
defparam \Reg[12][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N30
cycloneive_lcell_comb \Mux53~17 (
// Equation(s):
// \Mux53~17_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[13][10]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[12][10]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[12][10]~q ),
	.datad(\Reg[13][10]~q ),
	.cin(gnd),
	.combout(\Mux53~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~17 .lut_mask = 16'hDC98;
defparam \Mux53~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N12
cycloneive_lcell_comb \Mux53~18 (
// Equation(s):
// \Mux53~18_combout  = (\Mux53~17_combout  & (((\Reg[15][10]~q ) # (!ifid_ifinstr_o_17)))) # (!\Mux53~17_combout  & (\Reg[14][10]~q  & ((ifid_ifinstr_o_17))))

	.dataa(\Reg[14][10]~q ),
	.datab(\Mux53~17_combout ),
	.datac(\Reg[15][10]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux53~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~18 .lut_mask = 16'hE2CC;
defparam \Mux53~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N30
cycloneive_lcell_comb \Mux53~12 (
// Equation(s):
// \Mux53~12_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & (\Reg[5][10]~q )) # (!ifid_ifinstr_o_16 & ((\Reg[4][10]~q )))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[5][10]~q ),
	.datac(\Reg[4][10]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux53~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~12 .lut_mask = 16'hEE50;
defparam \Mux53~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N10
cycloneive_lcell_comb \Mux53~13 (
// Equation(s):
// \Mux53~13_combout  = (\Mux53~12_combout  & (((\Reg[7][10]~q ) # (!ifid_ifinstr_o_17)))) # (!\Mux53~12_combout  & (\Reg[6][10]~q  & ((ifid_ifinstr_o_17))))

	.dataa(\Reg[6][10]~q ),
	.datab(\Mux53~12_combout ),
	.datac(\Reg[7][10]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux53~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~13 .lut_mask = 16'hE2CC;
defparam \Mux53~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N20
cycloneive_lcell_comb \Mux53~14 (
// Equation(s):
// \Mux53~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][10]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][10]~q )))))

	.dataa(\Reg[3][10]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[1][10]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux53~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~14 .lut_mask = 16'hB800;
defparam \Mux53~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N10
cycloneive_lcell_comb \Mux53~15 (
// Equation(s):
// \Mux53~15_combout  = (\Mux53~14_combout ) # ((ifid_ifinstr_o_17 & (\Reg[2][10]~q  & !ifid_ifinstr_o_16)))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux53~14_combout ),
	.datac(\Reg[2][10]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux53~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~15 .lut_mask = 16'hCCEC;
defparam \Mux53~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N8
cycloneive_lcell_comb \Mux53~16 (
// Equation(s):
// \Mux53~16_combout  = (ifid_ifinstr_o_18 & ((\Mux53~13_combout ) # ((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (((!ifid_ifinstr_o_19 & \Mux53~15_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux53~13_combout ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux53~15_combout ),
	.cin(gnd),
	.combout(\Mux53~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~16 .lut_mask = 16'hADA8;
defparam \Mux53~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N16
cycloneive_lcell_comb \Mux53~10 (
// Equation(s):
// \Mux53~10_combout  = (ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16) # ((\Reg[10][10]~q )))) # (!ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & ((\Reg[8][10]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[10][10]~q ),
	.datad(\Reg[8][10]~q ),
	.cin(gnd),
	.combout(\Mux53~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~10 .lut_mask = 16'hB9A8;
defparam \Mux53~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N24
cycloneive_lcell_comb \Reg[9][10]~feeder (
// Equation(s):
// \Reg[9][10]~feeder_combout  = \wdat~33_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat15),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[9][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[9][10]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[9][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y32_N25
dffeas \Reg[9][10] (
	.clk(!CLK),
	.d(\Reg[9][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[9][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[9][10] .is_wysiwyg = "true";
defparam \Reg[9][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N14
cycloneive_lcell_comb \Mux53~11 (
// Equation(s):
// \Mux53~11_combout  = (ifid_ifinstr_o_16 & ((\Mux53~10_combout  & (\Reg[11][10]~q )) # (!\Mux53~10_combout  & ((\Reg[9][10]~q ))))) # (!ifid_ifinstr_o_16 & (((\Mux53~10_combout ))))

	.dataa(\Reg[11][10]~q ),
	.datab(ifid_ifinstr_o_16),
	.datac(\Mux53~10_combout ),
	.datad(\Reg[9][10]~q ),
	.cin(gnd),
	.combout(\Mux53~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~11 .lut_mask = 16'hBCB0;
defparam \Mux53~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N12
cycloneive_lcell_comb \Mux52~7 (
// Equation(s):
// \Mux52~7_combout  = (ifid_ifinstr_o_18 & (((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[27][11]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[19][11]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[19][11]~q ),
	.datac(\Reg[27][11]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux52~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~7 .lut_mask = 16'hFA44;
defparam \Mux52~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N14
cycloneive_lcell_comb \Mux52~8 (
// Equation(s):
// \Mux52~8_combout  = (ifid_ifinstr_o_18 & ((\Mux52~7_combout  & (\Reg[31][11]~q )) # (!\Mux52~7_combout  & ((\Reg[23][11]~q ))))) # (!ifid_ifinstr_o_18 & (\Mux52~7_combout ))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Mux52~7_combout ),
	.datac(\Reg[31][11]~q ),
	.datad(\Reg[23][11]~q ),
	.cin(gnd),
	.combout(\Mux52~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~8 .lut_mask = 16'hE6C4;
defparam \Mux52~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N8
cycloneive_lcell_comb \Mux52~3 (
// Equation(s):
// \Mux52~3_combout  = (\Mux52~2_combout  & (((\Reg[30][11]~q )) # (!ifid_ifinstr_o_19))) # (!\Mux52~2_combout  & (ifid_ifinstr_o_19 & (\Reg[26][11]~q )))

	.dataa(\Mux52~2_combout ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[26][11]~q ),
	.datad(\Reg[30][11]~q ),
	.cin(gnd),
	.combout(\Mux52~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~3 .lut_mask = 16'hEA62;
defparam \Mux52~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N29
dffeas \Reg[16][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~12_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[16][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[16][11] .is_wysiwyg = "true";
defparam \Reg[16][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N28
cycloneive_lcell_comb \Mux52~4 (
// Equation(s):
// \Mux52~4_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & ((\Reg[20][11]~q ))) # (!ifid_ifinstr_o_18 & (\Reg[16][11]~q ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[16][11]~q ),
	.datad(\Reg[20][11]~q ),
	.cin(gnd),
	.combout(\Mux52~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~4 .lut_mask = 16'hDC98;
defparam \Mux52~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N17
dffeas \Reg[24][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][11] .is_wysiwyg = "true";
defparam \Reg[24][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N22
cycloneive_lcell_comb \Mux52~5 (
// Equation(s):
// \Mux52~5_combout  = (ifid_ifinstr_o_19 & ((\Mux52~4_combout  & (\Reg[28][11]~q )) # (!\Mux52~4_combout  & ((\Reg[24][11]~q ))))) # (!ifid_ifinstr_o_19 & (\Mux52~4_combout ))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Mux52~4_combout ),
	.datac(\Reg[28][11]~q ),
	.datad(\Reg[24][11]~q ),
	.cin(gnd),
	.combout(\Mux52~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~5 .lut_mask = 16'hE6C4;
defparam \Mux52~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N14
cycloneive_lcell_comb \Mux52~6 (
// Equation(s):
// \Mux52~6_combout  = (ifid_ifinstr_o_17 & ((\Mux52~3_combout ) # ((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & (((!ifid_ifinstr_o_16 & \Mux52~5_combout ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux52~3_combout ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux52~5_combout ),
	.cin(gnd),
	.combout(\Mux52~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~6 .lut_mask = 16'hADA8;
defparam \Mux52~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N20
cycloneive_lcell_comb \Mux52~0 (
// Equation(s):
// \Mux52~0_combout  = (ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18) # ((\Reg[25][11]~q )))) # (!ifid_ifinstr_o_19 & (!ifid_ifinstr_o_18 & (\Reg[17][11]~q )))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[17][11]~q ),
	.datad(\Reg[25][11]~q ),
	.cin(gnd),
	.combout(\Mux52~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~0 .lut_mask = 16'hBA98;
defparam \Mux52~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N30
cycloneive_lcell_comb \Mux52~1 (
// Equation(s):
// \Mux52~1_combout  = (ifid_ifinstr_o_18 & ((\Mux52~0_combout  & ((\Reg[29][11]~q ))) # (!\Mux52~0_combout  & (\Reg[21][11]~q )))) # (!ifid_ifinstr_o_18 & (((\Mux52~0_combout ))))

	.dataa(\Reg[21][11]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[29][11]~q ),
	.datad(\Mux52~0_combout ),
	.cin(gnd),
	.combout(\Mux52~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~1 .lut_mask = 16'hF388;
defparam \Mux52~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N14
cycloneive_lcell_comb \Mux52~14 (
// Equation(s):
// \Mux52~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[3][11]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[1][11]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[3][11]~q ),
	.datac(\Reg[1][11]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux52~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~14 .lut_mask = 16'h88A0;
defparam \Mux52~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N22
cycloneive_lcell_comb \Mux52~15 (
// Equation(s):
// \Mux52~15_combout  = (\Mux52~14_combout ) # ((ifid_ifinstr_o_17 & (!ifid_ifinstr_o_16 & \Reg[2][11]~q )))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[2][11]~q ),
	.datad(\Mux52~14_combout ),
	.cin(gnd),
	.combout(\Mux52~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~15 .lut_mask = 16'hFF20;
defparam \Mux52~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y36_N27
dffeas \Reg[8][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[8][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[8][11] .is_wysiwyg = "true";
defparam \Reg[8][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N26
cycloneive_lcell_comb \Mux52~12 (
// Equation(s):
// \Mux52~12_combout  = (ifid_ifinstr_o_16 & (((ifid_ifinstr_o_17)))) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & (\Reg[10][11]~q )) # (!ifid_ifinstr_o_17 & ((\Reg[8][11]~q )))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[10][11]~q ),
	.datac(\Reg[8][11]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux52~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~12 .lut_mask = 16'hEE50;
defparam \Mux52~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N20
cycloneive_lcell_comb \Mux52~13 (
// Equation(s):
// \Mux52~13_combout  = (\Mux52~12_combout  & (((\Reg[11][11]~q ) # (!ifid_ifinstr_o_16)))) # (!\Mux52~12_combout  & (\Reg[9][11]~q  & ((ifid_ifinstr_o_16))))

	.dataa(\Reg[9][11]~q ),
	.datab(\Mux52~12_combout ),
	.datac(\Reg[11][11]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux52~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~13 .lut_mask = 16'hE2CC;
defparam \Mux52~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N2
cycloneive_lcell_comb \Mux52~16 (
// Equation(s):
// \Mux52~16_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Mux52~13_combout ))) # (!ifid_ifinstr_o_19 & (\Mux52~15_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Mux52~15_combout ),
	.datad(\Mux52~13_combout ),
	.cin(gnd),
	.combout(\Mux52~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~16 .lut_mask = 16'hDC98;
defparam \Mux52~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N16
cycloneive_lcell_comb \Mux52~10 (
// Equation(s):
// \Mux52~10_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[5][11]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[4][11]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[4][11]~q ),
	.datac(\Reg[5][11]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux52~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~10 .lut_mask = 16'hFA44;
defparam \Mux52~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N28
cycloneive_lcell_comb \Mux52~11 (
// Equation(s):
// \Mux52~11_combout  = (ifid_ifinstr_o_17 & ((\Mux52~10_combout  & (\Reg[7][11]~q )) # (!\Mux52~10_combout  & ((\Reg[6][11]~q ))))) # (!ifid_ifinstr_o_17 & (((\Mux52~10_combout ))))

	.dataa(\Reg[7][11]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[6][11]~q ),
	.datad(\Mux52~10_combout ),
	.cin(gnd),
	.combout(\Mux52~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~11 .lut_mask = 16'hBBC0;
defparam \Mux52~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N27
dffeas \Reg[12][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat14),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[12][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[12][11] .is_wysiwyg = "true";
defparam \Reg[12][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N26
cycloneive_lcell_comb \Mux52~17 (
// Equation(s):
// \Mux52~17_combout  = (ifid_ifinstr_o_17 & (ifid_ifinstr_o_16)) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[13][11]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[12][11]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[12][11]~q ),
	.datad(\Reg[13][11]~q ),
	.cin(gnd),
	.combout(\Mux52~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~17 .lut_mask = 16'hDC98;
defparam \Mux52~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N12
cycloneive_lcell_comb \Mux52~18 (
// Equation(s):
// \Mux52~18_combout  = (ifid_ifinstr_o_17 & ((\Mux52~17_combout  & ((\Reg[15][11]~q ))) # (!\Mux52~17_combout  & (\Reg[14][11]~q )))) # (!ifid_ifinstr_o_17 & (((\Mux52~17_combout ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[14][11]~q ),
	.datac(\Mux52~17_combout ),
	.datad(\Reg[15][11]~q ),
	.cin(gnd),
	.combout(\Mux52~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~18 .lut_mask = 16'hF858;
defparam \Mux52~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N22
cycloneive_lcell_comb \Mux51~0 (
// Equation(s):
// \Mux51~0_combout  = (ifid_ifinstr_o_19 & (ifid_ifinstr_o_18)) # (!ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18 & (\Reg[21][12]~q )) # (!ifid_ifinstr_o_18 & ((\Reg[17][12]~q )))))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[21][12]~q ),
	.datad(\Reg[17][12]~q ),
	.cin(gnd),
	.combout(\Mux51~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~0 .lut_mask = 16'hD9C8;
defparam \Mux51~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N4
cycloneive_lcell_comb \Mux51~1 (
// Equation(s):
// \Mux51~1_combout  = (ifid_ifinstr_o_19 & ((\Mux51~0_combout  & ((\Reg[29][12]~q ))) # (!\Mux51~0_combout  & (\Reg[25][12]~q )))) # (!ifid_ifinstr_o_19 & (((\Mux51~0_combout ))))

	.dataa(\Reg[25][12]~q ),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[29][12]~q ),
	.datad(\Mux51~0_combout ),
	.cin(gnd),
	.combout(\Mux51~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~1 .lut_mask = 16'hF388;
defparam \Mux51~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N16
cycloneive_lcell_comb \Mux51~7 (
// Equation(s):
// \Mux51~7_combout  = (ifid_ifinstr_o_18 & (((\Reg[23][12]~q ) # (ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (\Reg[19][12]~q  & ((!ifid_ifinstr_o_19))))

	.dataa(\Reg[19][12]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[23][12]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux51~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~7 .lut_mask = 16'hCCE2;
defparam \Mux51~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N26
cycloneive_lcell_comb \Mux51~8 (
// Equation(s):
// \Mux51~8_combout  = (ifid_ifinstr_o_19 & ((\Mux51~7_combout  & ((\Reg[31][12]~q ))) # (!\Mux51~7_combout  & (\Reg[27][12]~q )))) # (!ifid_ifinstr_o_19 & (((\Mux51~7_combout ))))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Reg[27][12]~q ),
	.datac(\Reg[31][12]~q ),
	.datad(\Mux51~7_combout ),
	.cin(gnd),
	.combout(\Mux51~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~8 .lut_mask = 16'hF588;
defparam \Mux51~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N23
dffeas \Reg[18][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat13),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[18][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[18][12] .is_wysiwyg = "true";
defparam \Reg[18][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N22
cycloneive_lcell_comb \Mux51~2 (
// Equation(s):
// \Mux51~2_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[26][12]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[18][12]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[18][12]~q ),
	.datad(\Reg[26][12]~q ),
	.cin(gnd),
	.combout(\Mux51~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~2 .lut_mask = 16'hDC98;
defparam \Mux51~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N22
cycloneive_lcell_comb \Mux51~3 (
// Equation(s):
// \Mux51~3_combout  = (ifid_ifinstr_o_18 & ((\Mux51~2_combout  & (\Reg[30][12]~q )) # (!\Mux51~2_combout  & ((\Reg[22][12]~q ))))) # (!ifid_ifinstr_o_18 & (((\Mux51~2_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[30][12]~q ),
	.datac(\Mux51~2_combout ),
	.datad(\Reg[22][12]~q ),
	.cin(gnd),
	.combout(\Mux51~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~3 .lut_mask = 16'hDAD0;
defparam \Mux51~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N12
cycloneive_lcell_comb \Reg[24][12]~feeder (
// Equation(s):
// \Reg[24][12]~feeder_combout  = \wdat~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat13),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[24][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[24][12]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[24][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N13
dffeas \Reg[24][12] (
	.clk(!CLK),
	.d(\Reg[24][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[24][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[24][12] .is_wysiwyg = "true";
defparam \Reg[24][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N22
cycloneive_lcell_comb \Mux51~4 (
// Equation(s):
// \Mux51~4_combout  = (ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18) # ((\Reg[24][12]~q )))) # (!ifid_ifinstr_o_19 & (!ifid_ifinstr_o_18 & (\Reg[16][12]~q )))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[16][12]~q ),
	.datad(\Reg[24][12]~q ),
	.cin(gnd),
	.combout(\Mux51~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~4 .lut_mask = 16'hBA98;
defparam \Mux51~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N26
cycloneive_lcell_comb \Mux51~5 (
// Equation(s):
// \Mux51~5_combout  = (ifid_ifinstr_o_18 & ((\Mux51~4_combout  & ((\Reg[28][12]~q ))) # (!\Mux51~4_combout  & (\Reg[20][12]~q )))) # (!ifid_ifinstr_o_18 & (((\Mux51~4_combout ))))

	.dataa(\Reg[20][12]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[28][12]~q ),
	.datad(\Mux51~4_combout ),
	.cin(gnd),
	.combout(\Mux51~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~5 .lut_mask = 16'hF388;
defparam \Mux51~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y36_N8
cycloneive_lcell_comb \Mux51~6 (
// Equation(s):
// \Mux51~6_combout  = (ifid_ifinstr_o_17 & ((\Mux51~3_combout ) # ((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & (((\Mux51~5_combout  & !ifid_ifinstr_o_16))))

	.dataa(\Mux51~3_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Mux51~5_combout ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux51~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~6 .lut_mask = 16'hCCB8;
defparam \Mux51~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N0
cycloneive_lcell_comb \Mux51~17 (
// Equation(s):
// \Mux51~17_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17) # ((\Reg[13][12]~q )))) # (!ifid_ifinstr_o_16 & (!ifid_ifinstr_o_17 & ((\Reg[12][12]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[13][12]~q ),
	.datad(\Reg[12][12]~q ),
	.cin(gnd),
	.combout(\Mux51~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~17 .lut_mask = 16'hB9A8;
defparam \Mux51~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N0
cycloneive_lcell_comb \Mux51~18 (
// Equation(s):
// \Mux51~18_combout  = (ifid_ifinstr_o_17 & ((\Mux51~17_combout  & (\Reg[15][12]~q )) # (!\Mux51~17_combout  & ((\Reg[14][12]~q ))))) # (!ifid_ifinstr_o_17 & (((\Mux51~17_combout ))))

	.dataa(\Reg[15][12]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[14][12]~q ),
	.datad(\Mux51~17_combout ),
	.cin(gnd),
	.combout(\Mux51~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~18 .lut_mask = 16'hBBC0;
defparam \Mux51~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N28
cycloneive_lcell_comb \Mux51~10 (
// Equation(s):
// \Mux51~10_combout  = (ifid_ifinstr_o_17 & (((\Reg[10][12]~q ) # (ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & (\Reg[8][12]~q  & ((!ifid_ifinstr_o_16))))

	.dataa(\Reg[8][12]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[10][12]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux51~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~10 .lut_mask = 16'hCCE2;
defparam \Mux51~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N28
cycloneive_lcell_comb \Mux51~11 (
// Equation(s):
// \Mux51~11_combout  = (\Mux51~10_combout  & ((\Reg[11][12]~q ) # ((!ifid_ifinstr_o_16)))) # (!\Mux51~10_combout  & (((\Reg[9][12]~q  & ifid_ifinstr_o_16))))

	.dataa(\Reg[11][12]~q ),
	.datab(\Mux51~10_combout ),
	.datac(\Reg[9][12]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux51~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~11 .lut_mask = 16'hB8CC;
defparam \Mux51~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y39_N2
cycloneive_lcell_comb \Mux51~13 (
// Equation(s):
// \Mux51~13_combout  = (\Mux51~12_combout  & (((\Reg[7][12]~q )) # (!ifid_ifinstr_o_17))) # (!\Mux51~12_combout  & (ifid_ifinstr_o_17 & ((\Reg[6][12]~q ))))

	.dataa(\Mux51~12_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[7][12]~q ),
	.datad(\Reg[6][12]~q ),
	.cin(gnd),
	.combout(\Mux51~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~13 .lut_mask = 16'hE6A2;
defparam \Mux51~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N18
cycloneive_lcell_comb \Mux51~15 (
// Equation(s):
// \Mux51~15_combout  = (\Mux51~14_combout ) # ((ifid_ifinstr_o_17 & (\Reg[2][12]~q  & !ifid_ifinstr_o_16)))

	.dataa(\Mux51~14_combout ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[2][12]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux51~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~15 .lut_mask = 16'hAAEA;
defparam \Mux51~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N8
cycloneive_lcell_comb \Mux51~16 (
// Equation(s):
// \Mux51~16_combout  = (ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19) # ((\Mux51~13_combout )))) # (!ifid_ifinstr_o_18 & (!ifid_ifinstr_o_19 & ((\Mux51~15_combout ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Mux51~13_combout ),
	.datad(\Mux51~15_combout ),
	.cin(gnd),
	.combout(\Mux51~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~16 .lut_mask = 16'hB9A8;
defparam \Mux51~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y37_N14
cycloneive_lcell_comb \Mux50~0 (
// Equation(s):
// \Mux50~0_combout  = (ifid_ifinstr_o_19 & ((ifid_ifinstr_o_18) # ((\Reg[25][13]~q )))) # (!ifid_ifinstr_o_19 & (!ifid_ifinstr_o_18 & (\Reg[17][13]~q )))

	.dataa(ifid_ifinstr_o_19),
	.datab(ifid_ifinstr_o_18),
	.datac(\Reg[17][13]~q ),
	.datad(\Reg[25][13]~q ),
	.cin(gnd),
	.combout(\Mux50~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~0 .lut_mask = 16'hBA98;
defparam \Mux50~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N6
cycloneive_lcell_comb \Mux50~1 (
// Equation(s):
// \Mux50~1_combout  = (\Mux50~0_combout  & ((\Reg[29][13]~q ) # ((!ifid_ifinstr_o_18)))) # (!\Mux50~0_combout  & (((ifid_ifinstr_o_18 & \Reg[21][13]~q ))))

	.dataa(\Reg[29][13]~q ),
	.datab(\Mux50~0_combout ),
	.datac(ifid_ifinstr_o_18),
	.datad(\Reg[21][13]~q ),
	.cin(gnd),
	.combout(\Mux50~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~1 .lut_mask = 16'hBC8C;
defparam \Mux50~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N18
cycloneive_lcell_comb \Mux50~7 (
// Equation(s):
// \Mux50~7_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & ((\Reg[27][13]~q ))) # (!ifid_ifinstr_o_19 & (\Reg[19][13]~q ))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Reg[19][13]~q ),
	.datad(\Reg[27][13]~q ),
	.cin(gnd),
	.combout(\Mux50~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~7 .lut_mask = 16'hDC98;
defparam \Mux50~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N18
cycloneive_lcell_comb \Mux50~8 (
// Equation(s):
// \Mux50~8_combout  = (ifid_ifinstr_o_18 & ((\Mux50~7_combout  & ((\Reg[31][13]~q ))) # (!\Mux50~7_combout  & (\Reg[23][13]~q )))) # (!ifid_ifinstr_o_18 & (((\Mux50~7_combout ))))

	.dataa(\Reg[23][13]~q ),
	.datab(\Reg[31][13]~q ),
	.datac(ifid_ifinstr_o_18),
	.datad(\Mux50~7_combout ),
	.cin(gnd),
	.combout(\Mux50~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~8 .lut_mask = 16'hCFA0;
defparam \Mux50~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N0
cycloneive_lcell_comb \Mux50~4 (
// Equation(s):
// \Mux50~4_combout  = (ifid_ifinstr_o_18 & ((\Reg[20][13]~q ) # ((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (((!ifid_ifinstr_o_19 & \Reg[16][13]~q ))))

	.dataa(\Reg[20][13]~q ),
	.datab(ifid_ifinstr_o_18),
	.datac(ifid_ifinstr_o_19),
	.datad(\Reg[16][13]~q ),
	.cin(gnd),
	.combout(\Mux50~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~4 .lut_mask = 16'hCBC8;
defparam \Mux50~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N26
cycloneive_lcell_comb \Reg[28][13]~feeder (
// Equation(s):
// \Reg[28][13]~feeder_combout  = \wdat~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(wdat12),
	.datad(gnd),
	.cin(gnd),
	.combout(\Reg[28][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[28][13]~feeder .lut_mask = 16'hF0F0;
defparam \Reg[28][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N27
dffeas \Reg[28][13] (
	.clk(!CLK),
	.d(\Reg[28][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[28][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[28][13] .is_wysiwyg = "true";
defparam \Reg[28][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N6
cycloneive_lcell_comb \Mux50~5 (
// Equation(s):
// \Mux50~5_combout  = (ifid_ifinstr_o_19 & ((\Mux50~4_combout  & ((\Reg[28][13]~q ))) # (!\Mux50~4_combout  & (\Reg[24][13]~q )))) # (!ifid_ifinstr_o_19 & (\Mux50~4_combout ))

	.dataa(ifid_ifinstr_o_19),
	.datab(\Mux50~4_combout ),
	.datac(\Reg[24][13]~q ),
	.datad(\Reg[28][13]~q ),
	.cin(gnd),
	.combout(\Mux50~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~5 .lut_mask = 16'hEC64;
defparam \Mux50~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N10
cycloneive_lcell_comb \Reg[22][13]~feeder (
// Equation(s):
// \Reg[22][13]~feeder_combout  = \wdat~27_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(wdat12),
	.cin(gnd),
	.combout(\Reg[22][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \Reg[22][13]~feeder .lut_mask = 16'hFF00;
defparam \Reg[22][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y36_N11
dffeas \Reg[22][13] (
	.clk(!CLK),
	.d(\Reg[22][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~7_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[22][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[22][13] .is_wysiwyg = "true";
defparam \Reg[22][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N10
cycloneive_lcell_comb \Mux50~2 (
// Equation(s):
// \Mux50~2_combout  = (ifid_ifinstr_o_18 & ((\Reg[22][13]~q ) # ((ifid_ifinstr_o_19)))) # (!ifid_ifinstr_o_18 & (((\Reg[18][13]~q  & !ifid_ifinstr_o_19))))

	.dataa(ifid_ifinstr_o_18),
	.datab(\Reg[22][13]~q ),
	.datac(\Reg[18][13]~q ),
	.datad(ifid_ifinstr_o_19),
	.cin(gnd),
	.combout(\Mux50~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~2 .lut_mask = 16'hAAD8;
defparam \Mux50~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N0
cycloneive_lcell_comb \Mux50~3 (
// Equation(s):
// \Mux50~3_combout  = (ifid_ifinstr_o_19 & ((\Mux50~2_combout  & (\Reg[30][13]~q )) # (!\Mux50~2_combout  & ((\Reg[26][13]~q ))))) # (!ifid_ifinstr_o_19 & (((\Mux50~2_combout ))))

	.dataa(\Reg[30][13]~q ),
	.datab(\Reg[26][13]~q ),
	.datac(ifid_ifinstr_o_19),
	.datad(\Mux50~2_combout ),
	.cin(gnd),
	.combout(\Mux50~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~3 .lut_mask = 16'hAFC0;
defparam \Mux50~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N2
cycloneive_lcell_comb \Mux50~6 (
// Equation(s):
// \Mux50~6_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16) # (\Mux50~3_combout )))) # (!ifid_ifinstr_o_17 & (\Mux50~5_combout  & (!ifid_ifinstr_o_16)))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux50~5_combout ),
	.datac(ifid_ifinstr_o_16),
	.datad(\Mux50~3_combout ),
	.cin(gnd),
	.combout(\Mux50~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~6 .lut_mask = 16'hAEA4;
defparam \Mux50~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y36_N6
cycloneive_lcell_comb \Mux50~12 (
// Equation(s):
// \Mux50~12_combout  = (ifid_ifinstr_o_16 & (ifid_ifinstr_o_17)) # (!ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[10][13]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[8][13]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[8][13]~q ),
	.datad(\Reg[10][13]~q ),
	.cin(gnd),
	.combout(\Mux50~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~12 .lut_mask = 16'hDC98;
defparam \Mux50~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N30
cycloneive_lcell_comb \Mux50~13 (
// Equation(s):
// \Mux50~13_combout  = (ifid_ifinstr_o_16 & ((\Mux50~12_combout  & ((\Reg[11][13]~q ))) # (!\Mux50~12_combout  & (\Reg[9][13]~q )))) # (!ifid_ifinstr_o_16 & (((\Mux50~12_combout ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(\Reg[9][13]~q ),
	.datac(\Reg[11][13]~q ),
	.datad(\Mux50~12_combout ),
	.cin(gnd),
	.combout(\Mux50~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~13 .lut_mask = 16'hF588;
defparam \Mux50~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N2
cycloneive_lcell_comb \Mux50~14 (
// Equation(s):
// \Mux50~14_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17 & ((\Reg[3][13]~q ))) # (!ifid_ifinstr_o_17 & (\Reg[1][13]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(ifid_ifinstr_o_16),
	.datac(\Reg[1][13]~q ),
	.datad(\Reg[3][13]~q ),
	.cin(gnd),
	.combout(\Mux50~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~14 .lut_mask = 16'hC840;
defparam \Mux50~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N28
cycloneive_lcell_comb \Mux50~15 (
// Equation(s):
// \Mux50~15_combout  = (\Mux50~14_combout ) # ((ifid_ifinstr_o_17 & (\Reg[2][13]~q  & !ifid_ifinstr_o_16)))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Mux50~14_combout ),
	.datac(\Reg[2][13]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux50~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~15 .lut_mask = 16'hCCEC;
defparam \Mux50~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y36_N14
cycloneive_lcell_comb \Mux50~16 (
// Equation(s):
// \Mux50~16_combout  = (ifid_ifinstr_o_18 & (ifid_ifinstr_o_19)) # (!ifid_ifinstr_o_18 & ((ifid_ifinstr_o_19 & (\Mux50~13_combout )) # (!ifid_ifinstr_o_19 & ((\Mux50~15_combout )))))

	.dataa(ifid_ifinstr_o_18),
	.datab(ifid_ifinstr_o_19),
	.datac(\Mux50~13_combout ),
	.datad(\Mux50~15_combout ),
	.cin(gnd),
	.combout(\Mux50~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~16 .lut_mask = 16'hD9C8;
defparam \Mux50~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N8
cycloneive_lcell_comb \Mux50~17 (
// Equation(s):
// \Mux50~17_combout  = (ifid_ifinstr_o_16 & ((ifid_ifinstr_o_17) # ((\Reg[13][13]~q )))) # (!ifid_ifinstr_o_16 & (!ifid_ifinstr_o_17 & ((\Reg[12][13]~q ))))

	.dataa(ifid_ifinstr_o_16),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[13][13]~q ),
	.datad(\Reg[12][13]~q ),
	.cin(gnd),
	.combout(\Mux50~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~17 .lut_mask = 16'hB9A8;
defparam \Mux50~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N14
cycloneive_lcell_comb \Mux50~18 (
// Equation(s):
// \Mux50~18_combout  = (ifid_ifinstr_o_17 & ((\Mux50~17_combout  & (\Reg[15][13]~q )) # (!\Mux50~17_combout  & ((\Reg[14][13]~q ))))) # (!ifid_ifinstr_o_17 & (((\Mux50~17_combout ))))

	.dataa(\Reg[15][13]~q ),
	.datab(ifid_ifinstr_o_17),
	.datac(\Reg[14][13]~q ),
	.datad(\Mux50~17_combout ),
	.cin(gnd),
	.combout(\Mux50~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~18 .lut_mask = 16'hBBC0;
defparam \Mux50~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y39_N23
dffeas \Reg[4][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~22_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[4][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[4][13] .is_wysiwyg = "true";
defparam \Reg[4][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y39_N25
dffeas \Reg[5][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(wdat12),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\Reg[5][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \Reg[5][13] .is_wysiwyg = "true";
defparam \Reg[5][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y39_N24
cycloneive_lcell_comb \Mux50~10 (
// Equation(s):
// \Mux50~10_combout  = (ifid_ifinstr_o_17 & (((ifid_ifinstr_o_16)))) # (!ifid_ifinstr_o_17 & ((ifid_ifinstr_o_16 & ((\Reg[5][13]~q ))) # (!ifid_ifinstr_o_16 & (\Reg[4][13]~q ))))

	.dataa(ifid_ifinstr_o_17),
	.datab(\Reg[4][13]~q ),
	.datac(\Reg[5][13]~q ),
	.datad(ifid_ifinstr_o_16),
	.cin(gnd),
	.combout(\Mux50~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~10 .lut_mask = 16'hFA44;
defparam \Mux50~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N20
cycloneive_lcell_comb \Mux50~11 (
// Equation(s):
// \Mux50~11_combout  = (\Mux50~10_combout  & ((\Reg[7][13]~q ) # ((!ifid_ifinstr_o_17)))) # (!\Mux50~10_combout  & (((\Reg[6][13]~q  & ifid_ifinstr_o_17))))

	.dataa(\Reg[7][13]~q ),
	.datab(\Mux50~10_combout ),
	.datac(\Reg[6][13]~q ),
	.datad(ifid_ifinstr_o_17),
	.cin(gnd),
	.combout(\Mux50~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~11 .lut_mask = 16'hB8CC;
defparam \Mux50~11 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module memory_control (
	exmem_ifdWEN_o,
	exmem_ifdREN_o,
	always1,
	always11,
	always12,
	ramstate,
	always13,
	devpor,
	devclrn,
	devoe);
input 	exmem_ifdWEN_o;
input 	exmem_ifdREN_o;
input 	always1;
input 	always11;
output 	always12;
input 	ramstate;
output 	always13;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X55_Y28_N14
cycloneive_lcell_comb \always1~0 (
// Equation(s):
// always12 = (!exmem_ifdREN_o & !exmem_ifdWEN_o)

	.dataa(gnd),
	.datab(exmem_ifdREN_o),
	.datac(exmem_ifdWEN_o),
	.datad(gnd),
	.cin(gnd),
	.combout(always12),
	.cout());
// synopsys translate_off
defparam \always1~0 .lut_mask = 16'h0303;
defparam \always1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N4
cycloneive_lcell_comb \always1~1 (
// Equation(s):
// always13 = (!ramstate & (always12 & ((always1) # (always11))))

	.dataa(always1),
	.datab(ramstate),
	.datac(always12),
	.datad(always11),
	.cin(gnd),
	.combout(always13),
	.cout());
// synopsys translate_off
defparam \always1~1 .lut_mask = 16'h3020;
defparam \always1~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module ram (
	is_in_use_reg,
	ramiframload_0,
	ramaddr,
	ramaddr1,
	ramaddr2,
	ramaddr3,
	ramaddr4,
	ramaddr5,
	ramaddr6,
	ramaddr7,
	ramaddr8,
	ramaddr9,
	ramaddr10,
	ramaddr11,
	ramaddr12,
	ramaddr13,
	ramaddr14,
	ramaddr15,
	\ramif.ramaddr ,
	ramaddr16,
	ramaddr17,
	ramaddr18,
	ramaddr19,
	ramaddr20,
	ramaddr21,
	ramaddr22,
	ramaddr23,
	ramaddr24,
	ramaddr25,
	ramaddr26,
	ramiframload_01,
	ramiframload_1,
	ramiframload_11,
	always1,
	always11,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_111,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	ramWEN,
	ramstore,
	ramREN,
	ramstate,
	ramstore1,
	ramstore2,
	ramstore3,
	ramstore4,
	ramstore5,
	ramstore6,
	ramstore7,
	ramstore8,
	ramstore9,
	ramstore10,
	ramstore11,
	ramstore12,
	ramstore13,
	ramstore14,
	ramstore15,
	ramstore16,
	ramstore17,
	ramstore18,
	ramstore19,
	ramstore20,
	ramstore21,
	ramstore22,
	ramstore23,
	ramstore24,
	ramstore25,
	ramstore26,
	ramstore27,
	ramstore28,
	ramstore29,
	ramstore30,
	ramstore31,
	ramaddr27,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	nRST,
	syiftbCTRL,
	syifWEN,
	syifREN,
	altera_internal_jtag1,
	nRST1,
	CLK,
	devpor,
	devclrn,
	devoe);
output 	is_in_use_reg;
output 	ramiframload_0;
input 	ramaddr;
input 	ramaddr1;
input 	ramaddr2;
input 	ramaddr3;
input 	ramaddr4;
input 	ramaddr5;
input 	ramaddr6;
input 	ramaddr7;
input 	ramaddr8;
input 	ramaddr9;
input 	ramaddr10;
input 	ramaddr11;
input 	ramaddr12;
input 	ramaddr13;
input 	ramaddr14;
input 	ramaddr15;
input 	[31:0] \ramif.ramaddr ;
input 	ramaddr16;
input 	ramaddr17;
input 	ramaddr18;
input 	ramaddr19;
input 	ramaddr20;
input 	ramaddr21;
input 	ramaddr22;
input 	ramaddr23;
input 	ramaddr24;
input 	ramaddr25;
input 	ramaddr26;
output 	ramiframload_01;
output 	ramiframload_1;
output 	ramiframload_11;
output 	always1;
output 	always11;
output 	ramiframload_2;
output 	ramiframload_3;
output 	ramiframload_4;
output 	ramiframload_5;
output 	ramiframload_6;
output 	ramiframload_7;
output 	ramiframload_8;
output 	ramiframload_9;
output 	ramiframload_10;
output 	ramiframload_111;
output 	ramiframload_12;
output 	ramiframload_13;
output 	ramiframload_14;
output 	ramiframload_15;
output 	ramiframload_16;
output 	ramiframload_17;
output 	ramiframload_18;
output 	ramiframload_19;
output 	ramiframload_20;
output 	ramiframload_21;
output 	ramiframload_22;
output 	ramiframload_23;
output 	ramiframload_24;
output 	ramiframload_25;
output 	ramiframload_26;
output 	ramiframload_27;
output 	ramiframload_28;
output 	ramiframload_29;
output 	ramiframload_30;
output 	ramiframload_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	ramWEN;
input 	ramstore;
input 	ramREN;
output 	ramstate;
input 	ramstore1;
input 	ramstore2;
input 	ramstore3;
input 	ramstore4;
input 	ramstore5;
input 	ramstore6;
input 	ramstore7;
input 	ramstore8;
input 	ramstore9;
input 	ramstore10;
input 	ramstore11;
input 	ramstore12;
input 	ramstore13;
input 	ramstore14;
input 	ramstore15;
input 	ramstore16;
input 	ramstore17;
input 	ramstore18;
input 	ramstore19;
input 	ramstore20;
input 	ramstore21;
input 	ramstore22;
input 	ramstore23;
input 	ramstore24;
input 	ramstore25;
input 	ramstore26;
input 	ramstore27;
input 	ramstore28;
input 	ramstore29;
input 	ramstore30;
input 	ramstore31;
input 	ramaddr27;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	nRST;
input 	syiftbCTRL;
input 	syifWEN;
input 	syifREN;
input 	altera_internal_jtag1;
input 	nRST1;
input 	CLK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ;
wire \Equal2~3_combout ;
wire \Equal2~8_combout ;
wire \Equal2~10_combout ;
wire \Equal2~17_combout ;
wire \addr[5]~feeder_combout ;
wire \addr[21]~feeder_combout ;
wire \always0~0_combout ;
wire \always0~1_combout ;
wire \Equal2~5_combout ;
wire \Equal2~7_combout ;
wire \Equal2~6_combout ;
wire \Equal2~9_combout ;
wire \Equal2~15_combout ;
wire \Equal2~16_combout ;
wire \Equal2~18_combout ;
wire \Equal2~19_combout ;
wire \Equal2~13_combout ;
wire \Equal2~12_combout ;
wire \Equal2~11_combout ;
wire \Equal2~14_combout ;
wire \Equal2~1_combout ;
wire \Equal2~0_combout ;
wire \Equal2~2_combout ;
wire \Equal2~4_combout ;
wire \Equal2~20_combout ;
wire \ramif.ramload[0]~1_combout ;
wire \ramif.ramload[1]~4_combout ;
wire [1:0] en;
wire [31:0] addr;
wire [0:0] \altsyncram_component|auto_generated|altsyncram1|address_reg_a ;


altsyncram_1 altsyncram_component(
	.ram_block3a32(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.ram_block3a0(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.ram_block3a33(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.ram_block3a1(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.ram_block3a34(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.ram_block3a2(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.ram_block3a35(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.ram_block3a3(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.ram_block3a36(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.ram_block3a4(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.ram_block3a37(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.ram_block3a5(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.ram_block3a38(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.ram_block3a6(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.ram_block3a39(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.ram_block3a7(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.ram_block3a40(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.ram_block3a8(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.ram_block3a41(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.ram_block3a9(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.ram_block3a42(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.ram_block3a10(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.ram_block3a43(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.ram_block3a11(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.ram_block3a44(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.ram_block3a12(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.ram_block3a45(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.ram_block3a13(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.ram_block3a46(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.ram_block3a14(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.ram_block3a47(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.ram_block3a15(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.ram_block3a48(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.ram_block3a16(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.ram_block3a49(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.ram_block3a17(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.ram_block3a50(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.ram_block3a18(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.ram_block3a51(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.ram_block3a19(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.ram_block3a52(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.ram_block3a20(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.ram_block3a53(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.ram_block3a21(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.ram_block3a54(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.ram_block3a22(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.ram_block3a55(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.ram_block3a23(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.ram_block3a56(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.ram_block3a24(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.ram_block3a57(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.ram_block3a25(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.ram_block3a58(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.ram_block3a26(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.ram_block3a59(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.ram_block3a27(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.ram_block3a60(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.ram_block3a28(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.ram_block3a61(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.ram_block3a29(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.ram_block3a62(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.ram_block3a30(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.ram_block3a63(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.ram_block3a31(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.address_a({gnd,ramaddr15,ramaddr12,ramaddr13,ramaddr10,ramaddr11,ramaddr8,ramaddr9,ramaddr6,ramaddr7,ramaddr4,ramaddr5,ramaddr2,ramaddr3}),
	.ramaddr(ramaddr14),
	.always1(always11),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.ramWEN(ramWEN),
	.data_a({ramstore31,ramstore30,ramstore29,ramstore28,ramstore27,ramstore26,ramstore25,ramstore24,ramstore23,ramstore22,ramstore21,ramstore20,ramstore19,ramstore18,ramstore17,ramstore16,ramstore15,ramstore14,ramstore13,ramstore12,ramstore11,ramstore10,ramstore9,ramstore8,ramstore7,ramstore6,
ramstore5,ramstore4,ramstore3,ramstore2,ramstore1,ramstore}),
	.ramaddr1(ramaddr27),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(CLK),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: FF_X54_Y33_N27
dffeas \addr[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[1]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[1] .is_wysiwyg = "true";
defparam \addr[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y28_N23
dffeas \addr[5] (
	.clk(CLK),
	.d(\addr[5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[5]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[5] .is_wysiwyg = "true";
defparam \addr[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y29_N9
dffeas \addr[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr7),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[6]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[6] .is_wysiwyg = "true";
defparam \addr[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y29_N31
dffeas \addr[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr6),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[7]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[7] .is_wysiwyg = "true";
defparam \addr[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N8
cycloneive_lcell_comb \Equal2~3 (
// Equation(s):
// \Equal2~3_combout  = (addr[7] & (\ramaddr~13_combout  & (\ramaddr~15_combout  $ (!addr[6])))) # (!addr[7] & (!\ramaddr~13_combout  & (\ramaddr~15_combout  $ (!addr[6]))))

	.dataa(addr[7]),
	.datab(ramaddr7),
	.datac(addr[6]),
	.datad(ramaddr6),
	.cin(gnd),
	.combout(\Equal2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~3 .lut_mask = 16'h8241;
defparam \Equal2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N9
dffeas \addr[9] (
	.clk(CLK),
	.d(ramaddr8),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[9]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[9] .is_wysiwyg = "true";
defparam \addr[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N31
dffeas \addr[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr10),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[11]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[11] .is_wysiwyg = "true";
defparam \addr[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N27
dffeas \addr[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr15),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[14]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[14] .is_wysiwyg = "true";
defparam \addr[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N1
dffeas \addr[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr27),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[15]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[15] .is_wysiwyg = "true";
defparam \addr[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N26
cycloneive_lcell_comb \Equal2~8 (
// Equation(s):
// \Equal2~8_combout  = (\ramaddr~29_combout  & (!addr[15] & (\ramaddr~31_combout  $ (!addr[14])))) # (!\ramaddr~29_combout  & (addr[15] & (\ramaddr~31_combout  $ (!addr[14]))))

	.dataa(ramaddr14),
	.datab(ramaddr15),
	.datac(addr[14]),
	.datad(addr[15]),
	.cin(gnd),
	.combout(\Equal2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~8 .lut_mask = 16'h4182;
defparam \Equal2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y31_N1
dffeas \addr[16] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr16),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[16]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[16] .is_wysiwyg = "true";
defparam \addr[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N31
dffeas \addr[17] (
	.clk(CLK),
	.d(\ramif.ramaddr [17]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[17]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[17] .is_wysiwyg = "true";
defparam \addr[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N0
cycloneive_lcell_comb \Equal2~10 (
// Equation(s):
// \Equal2~10_combout  = (\ramaddr~33_combout  & (addr[17] & (addr[16] $ (!\ramaddr~35_combout )))) # (!\ramaddr~33_combout  & (!addr[17] & (addr[16] $ (!\ramaddr~35_combout ))))

	.dataa(\ramif.ramaddr [17]),
	.datab(addr[17]),
	.datac(addr[16]),
	.datad(ramaddr16),
	.cin(gnd),
	.combout(\Equal2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~10 .lut_mask = 16'h9009;
defparam \Equal2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y32_N31
dffeas \addr[21] (
	.clk(CLK),
	.d(\addr[21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[21]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[21] .is_wysiwyg = "true";
defparam \addr[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y32_N3
dffeas \addr[27] (
	.clk(CLK),
	.d(\ramif.ramaddr [27]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[27]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[27] .is_wysiwyg = "true";
defparam \addr[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N15
dffeas \addr[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr24),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[28]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[28] .is_wysiwyg = "true";
defparam \addr[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N21
dffeas \addr[29] (
	.clk(CLK),
	.d(\ramif.ramaddr [29]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[29]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[29] .is_wysiwyg = "true";
defparam \addr[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N14
cycloneive_lcell_comb \Equal2~17 (
// Equation(s):
// \Equal2~17_combout  = (addr[29] & (\ramaddr~57_combout  & (\ramaddr~59_combout  $ (!addr[28])))) # (!addr[29] & (!\ramaddr~57_combout  & (\ramaddr~59_combout  $ (!addr[28]))))

	.dataa(addr[29]),
	.datab(ramaddr24),
	.datac(addr[28]),
	.datad(\ramif.ramaddr [29]),
	.cin(gnd),
	.combout(\Equal2~17_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~17 .lut_mask = 16'h8241;
defparam \Equal2~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y32_N13
dffeas \addr[31] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr25),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[31]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[31] .is_wysiwyg = "true";
defparam \addr[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N19
dffeas \en[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramWEN),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[0]),
	.prn(vcc));
// synopsys translate_off
defparam \en[0] .is_wysiwyg = "true";
defparam \en[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N22
cycloneive_lcell_comb \addr[5]~feeder (
// Equation(s):
// \addr[5]~feeder_combout  = \ramaddr~9_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr4),
	.cin(gnd),
	.combout(\addr[5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[5]~feeder .lut_mask = 16'hFF00;
defparam \addr[5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N30
cycloneive_lcell_comb \addr[21]~feeder (
// Equation(s):
// \addr[21]~feeder_combout  = \ramaddr~41_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(ramaddr19),
	.datad(gnd),
	.cin(gnd),
	.combout(\addr[21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[21]~feeder .lut_mask = 16'hF0F0;
defparam \addr[21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N28
cycloneive_lcell_comb \ramif.ramload[0]~0 (
// Equation(s):
// ramiframload_0 = (address_reg_a_0 & (ram_block3a321)) # (!address_reg_a_0 & ((ram_block3a01)))

	.dataa(gnd),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.cin(gnd),
	.combout(ramiframload_0),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[0]~0 .lut_mask = 16'hF3C0;
defparam \ramif.ramload[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N28
cycloneive_lcell_comb \ramif.ramload[0]~2 (
// Equation(s):
// ramiframload_01 = (ramiframload_0) # ((\nRST~input_o  & ((\ramif.ramload[0]~1_combout ) # (!\Equal2~20_combout ))))

	.dataa(\Equal2~20_combout ),
	.datab(ramiframload_0),
	.datac(nRST),
	.datad(\ramif.ramload[0]~1_combout ),
	.cin(gnd),
	.combout(ramiframload_01),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[0]~2 .lut_mask = 16'hFCDC;
defparam \ramif.ramload[0]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N22
cycloneive_lcell_comb \ramif.ramload[1]~3 (
// Equation(s):
// ramiframload_1 = (address_reg_a_0 & ((ram_block3a331))) # (!address_reg_a_0 & (ram_block3a110))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(gnd),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.cin(gnd),
	.combout(ramiframload_1),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[1]~3 .lut_mask = 16'hEE22;
defparam \ramif.ramload[1]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N12
cycloneive_lcell_comb \ramif.ramload[1]~5 (
// Equation(s):
// ramiframload_11 = (ramiframload_1 & (((\Equal2~20_combout  & \ramif.ramload[1]~4_combout )) # (!\nRST~input_o )))

	.dataa(\Equal2~20_combout ),
	.datab(ramiframload_1),
	.datac(nRST),
	.datad(\ramif.ramload[1]~4_combout ),
	.cin(gnd),
	.combout(ramiframload_11),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[1]~5 .lut_mask = 16'h8C0C;
defparam \ramif.ramload[1]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N18
cycloneive_lcell_comb \always1~0 (
// Equation(s):
// always1 = (!\syif.WEN~input_o  & (\syif.tbCTRL~input_o  & !\syif.REN~input_o ))

	.dataa(gnd),
	.datab(syifWEN),
	.datac(syiftbCTRL),
	.datad(syifREN),
	.cin(gnd),
	.combout(always1),
	.cout());
// synopsys translate_off
defparam \always1~0 .lut_mask = 16'h0030;
defparam \always1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N20
cycloneive_lcell_comb \always1~1 (
// Equation(s):
// always11 = ((!always1 & \Equal2~20_combout )) # (!\nRST~input_o )

	.dataa(always1),
	.datab(nRST),
	.datac(gnd),
	.datad(\Equal2~20_combout ),
	.cin(gnd),
	.combout(always11),
	.cout());
// synopsys translate_off
defparam \always1~1 .lut_mask = 16'h7733;
defparam \always1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N0
cycloneive_lcell_comb \ramif.ramload[2]~6 (
// Equation(s):
// ramiframload_2 = (always11 & ((address_reg_a_0 & (ram_block3a341)) # (!address_reg_a_0 & ((ram_block3a210)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.cin(gnd),
	.combout(ramiframload_2),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[2]~6 .lut_mask = 16'hC480;
defparam \ramif.ramload[2]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N18
cycloneive_lcell_comb \ramif.ramload[3]~7 (
// Equation(s):
// ramiframload_3 = (always11 & ((address_reg_a_0 & (ram_block3a351)) # (!address_reg_a_0 & ((ram_block3a310)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always11),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.cin(gnd),
	.combout(ramiframload_3),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[3]~7 .lut_mask = 16'hB080;
defparam \ramif.ramload[3]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N22
cycloneive_lcell_comb \ramif.ramload[4]~8 (
// Equation(s):
// ramiframload_4 = ((address_reg_a_0 & ((ram_block3a361))) # (!address_reg_a_0 & (ram_block3a410))) # (!always11)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.cin(gnd),
	.combout(ramiframload_4),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[4]~8 .lut_mask = 16'hFB73;
defparam \ramif.ramload[4]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N0
cycloneive_lcell_comb \ramif.ramload[5]~9 (
// Equation(s):
// ramiframload_5 = (always11 & ((address_reg_a_0 & (ram_block3a371)) # (!address_reg_a_0 & ((ram_block3a510)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.cin(gnd),
	.combout(ramiframload_5),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[5]~9 .lut_mask = 16'hC480;
defparam \ramif.ramload[5]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N12
cycloneive_lcell_comb \ramif.ramload[6]~10 (
// Equation(s):
// ramiframload_6 = ((address_reg_a_0 & ((ram_block3a381))) # (!address_reg_a_0 & (ram_block3a64))) # (!always11)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.cin(gnd),
	.combout(ramiframload_6),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[6]~10 .lut_mask = 16'hFB73;
defparam \ramif.ramload[6]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N30
cycloneive_lcell_comb \ramif.ramload[7]~11 (
// Equation(s):
// ramiframload_7 = ((address_reg_a_0 & ((ram_block3a391))) # (!address_reg_a_0 & (ram_block3a71))) # (!always11)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.cin(gnd),
	.combout(ramiframload_7),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[7]~11 .lut_mask = 16'hFB73;
defparam \ramif.ramload[7]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N12
cycloneive_lcell_comb \ramif.ramload[8]~12 (
// Equation(s):
// ramiframload_8 = (always11 & ((address_reg_a_0 & (ram_block3a401)) # (!address_reg_a_0 & ((ram_block3a81)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.cin(gnd),
	.combout(ramiframload_8),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[8]~12 .lut_mask = 16'hC480;
defparam \ramif.ramload[8]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N4
cycloneive_lcell_comb \ramif.ramload[9]~13 (
// Equation(s):
// ramiframload_9 = ((address_reg_a_0 & ((ram_block3a412))) # (!address_reg_a_0 & (ram_block3a91))) # (!always11)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.cin(gnd),
	.combout(ramiframload_9),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[9]~13 .lut_mask = 16'hFB73;
defparam \ramif.ramload[9]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N16
cycloneive_lcell_comb \ramif.ramload[10]~14 (
// Equation(s):
// ramiframload_10 = (always11 & ((address_reg_a_0 & ((ram_block3a421))) # (!address_reg_a_0 & (ram_block3a101))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.datad(always11),
	.cin(gnd),
	.combout(ramiframload_10),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[10]~14 .lut_mask = 16'hE400;
defparam \ramif.ramload[10]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N4
cycloneive_lcell_comb \ramif.ramload[11]~15 (
// Equation(s):
// ramiframload_111 = ((address_reg_a_0 & ((ram_block3a431))) # (!address_reg_a_0 & (ram_block3a112))) # (!always11)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.cin(gnd),
	.combout(ramiframload_111),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[11]~15 .lut_mask = 16'hFB3B;
defparam \ramif.ramload[11]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N16
cycloneive_lcell_comb \ramif.ramload[12]~16 (
// Equation(s):
// ramiframload_12 = ((address_reg_a_0 & (ram_block3a441)) # (!address_reg_a_0 & ((ram_block3a121)))) # (!always11)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.cin(gnd),
	.combout(ramiframload_12),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[12]~16 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[12]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N8
cycloneive_lcell_comb \ramif.ramload[13]~17 (
// Equation(s):
// ramiframload_13 = ((address_reg_a_0 & ((ram_block3a451))) # (!address_reg_a_0 & (ram_block3a131))) # (!always11)

	.dataa(always11),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.cin(gnd),
	.combout(ramiframload_13),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[13]~17 .lut_mask = 16'hFD75;
defparam \ramif.ramload[13]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N14
cycloneive_lcell_comb \ramif.ramload[14]~18 (
// Equation(s):
// ramiframload_14 = (always11 & ((address_reg_a_0 & (ram_block3a461)) # (!address_reg_a_0 & ((ram_block3a141)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.cin(gnd),
	.combout(ramiframload_14),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[14]~18 .lut_mask = 16'hC480;
defparam \ramif.ramload[14]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N22
cycloneive_lcell_comb \ramif.ramload[15]~19 (
// Equation(s):
// ramiframload_15 = ((address_reg_a_0 & ((ram_block3a471))) # (!address_reg_a_0 & (ram_block3a151))) # (!always11)

	.dataa(always11),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.cin(gnd),
	.combout(ramiframload_15),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[15]~19 .lut_mask = 16'hFD75;
defparam \ramif.ramload[15]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N14
cycloneive_lcell_comb \ramif.ramload[16]~20 (
// Equation(s):
// ramiframload_16 = ((address_reg_a_0 & (ram_block3a481)) # (!address_reg_a_0 & ((ram_block3a161)))) # (!always11)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.cin(gnd),
	.combout(ramiframload_16),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[16]~20 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[16]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N18
cycloneive_lcell_comb \ramif.ramload[17]~21 (
// Equation(s):
// ramiframload_17 = (always11 & ((address_reg_a_0 & ((ram_block3a491))) # (!address_reg_a_0 & (ram_block3a171))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.cin(gnd),
	.combout(ramiframload_17),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[17]~21 .lut_mask = 16'hC840;
defparam \ramif.ramload[17]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N24
cycloneive_lcell_comb \ramif.ramload[18]~22 (
// Equation(s):
// ramiframload_18 = (always11 & ((address_reg_a_0 & (ram_block3a501)) # (!address_reg_a_0 & ((ram_block3a181)))))

	.dataa(always11),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.cin(gnd),
	.combout(ramiframload_18),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[18]~22 .lut_mask = 16'hA280;
defparam \ramif.ramload[18]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N8
cycloneive_lcell_comb \ramif.ramload[19]~23 (
// Equation(s):
// ramiframload_19 = (always11 & ((address_reg_a_0 & (ram_block3a512)) # (!address_reg_a_0 & ((ram_block3a191)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.cin(gnd),
	.combout(ramiframload_19),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[19]~23 .lut_mask = 16'hC480;
defparam \ramif.ramload[19]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N8
cycloneive_lcell_comb \ramif.ramload[20]~24 (
// Equation(s):
// ramiframload_20 = ((address_reg_a_0 & ((ram_block3a521))) # (!address_reg_a_0 & (ram_block3a201))) # (!always11)

	.dataa(always11),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.cin(gnd),
	.combout(ramiframload_20),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[20]~24 .lut_mask = 16'hFD75;
defparam \ramif.ramload[20]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N24
cycloneive_lcell_comb \ramif.ramload[21]~25 (
// Equation(s):
// ramiframload_21 = (always11 & ((address_reg_a_0 & (ram_block3a531)) # (!address_reg_a_0 & ((ram_block3a212)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.cin(gnd),
	.combout(ramiframload_21),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[21]~25 .lut_mask = 16'hC480;
defparam \ramif.ramload[21]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N20
cycloneive_lcell_comb \ramif.ramload[22]~26 (
// Equation(s):
// ramiframload_22 = ((address_reg_a_0 & (ram_block3a541)) # (!address_reg_a_0 & ((ram_block3a221)))) # (!always11)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.datad(always11),
	.cin(gnd),
	.combout(ramiframload_22),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[22]~26 .lut_mask = 16'hB8FF;
defparam \ramif.ramload[22]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N24
cycloneive_lcell_comb \ramif.ramload[23]~27 (
// Equation(s):
// ramiframload_23 = ((address_reg_a_0 & (ram_block3a551)) # (!address_reg_a_0 & ((ram_block3a231)))) # (!always11)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.cin(gnd),
	.combout(ramiframload_23),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[23]~27 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[23]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N24
cycloneive_lcell_comb \ramif.ramload[24]~28 (
// Equation(s):
// ramiframload_24 = (always11 & ((address_reg_a_0 & ((ram_block3a561))) # (!address_reg_a_0 & (ram_block3a241))))

	.dataa(always11),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.cin(gnd),
	.combout(ramiframload_24),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[24]~28 .lut_mask = 16'hA820;
defparam \ramif.ramload[24]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N0
cycloneive_lcell_comb \ramif.ramload[25]~29 (
// Equation(s):
// ramiframload_25 = ((address_reg_a_0 & (ram_block3a571)) # (!address_reg_a_0 & ((ram_block3a251)))) # (!always11)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.cin(gnd),
	.combout(ramiframload_25),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[25]~29 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[25]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N10
cycloneive_lcell_comb \ramif.ramload[26]~30 (
// Equation(s):
// ramiframload_26 = (always11 & ((address_reg_a_0 & (ram_block3a581)) # (!address_reg_a_0 & ((ram_block3a261)))))

	.dataa(always11),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.cin(gnd),
	.combout(ramiframload_26),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[26]~30 .lut_mask = 16'hA280;
defparam \ramif.ramload[26]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N14
cycloneive_lcell_comb \ramif.ramload[27]~31 (
// Equation(s):
// ramiframload_27 = ((address_reg_a_0 & (ram_block3a591)) # (!address_reg_a_0 & ((ram_block3a271)))) # (!always11)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.cin(gnd),
	.combout(ramiframload_27),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[27]~31 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[27]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N4
cycloneive_lcell_comb \ramif.ramload[28]~32 (
// Equation(s):
// ramiframload_28 = ((address_reg_a_0 & ((ram_block3a601))) # (!address_reg_a_0 & (ram_block3a281))) # (!always11)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.cin(gnd),
	.combout(ramiframload_28),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[28]~32 .lut_mask = 16'hFB73;
defparam \ramif.ramload[28]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N8
cycloneive_lcell_comb \ramif.ramload[29]~33 (
// Equation(s):
// ramiframload_29 = ((address_reg_a_0 & (ram_block3a611)) # (!address_reg_a_0 & ((ram_block3a291)))) # (!always11)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always11),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.cin(gnd),
	.combout(ramiframload_29),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[29]~33 .lut_mask = 16'hF7B3;
defparam \ramif.ramload[29]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N20
cycloneive_lcell_comb \ramif.ramload[30]~34 (
// Equation(s):
// ramiframload_30 = (always11 & ((address_reg_a_0 & (ram_block3a621)) # (!address_reg_a_0 & ((ram_block3a301)))))

	.dataa(always11),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.cin(gnd),
	.combout(ramiframload_30),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[30]~34 .lut_mask = 16'hA280;
defparam \ramif.ramload[30]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N8
cycloneive_lcell_comb \ramif.ramload[31]~35 (
// Equation(s):
// ramiframload_31 = ((address_reg_a_0 & (ram_block3a631)) # (!address_reg_a_0 & ((ram_block3a312)))) # (!always11)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.datac(always11),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.cin(gnd),
	.combout(ramiframload_31),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[31]~35 .lut_mask = 16'hDF8F;
defparam \ramif.ramload[31]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N16
cycloneive_lcell_comb \ramstate~0 (
// Equation(s):
// ramstate = (\nRST~input_o  & ((\ramREN~0_combout  & ((\ramWEN~0_combout ) # (!\Equal2~20_combout ))) # (!\ramREN~0_combout  & (\ramWEN~0_combout  & !\Equal2~20_combout ))))

	.dataa(ramREN),
	.datab(ramWEN),
	.datac(nRST),
	.datad(\Equal2~20_combout ),
	.cin(gnd),
	.combout(ramstate),
	.cout());
// synopsys translate_off
defparam \ramstate~0 .lut_mask = 16'h80E0;
defparam \ramstate~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y28_N29
dffeas \en[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramREN),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[1]),
	.prn(vcc));
// synopsys translate_off
defparam \en[1] .is_wysiwyg = "true";
defparam \en[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N24
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// \always0~0_combout  = (en[0] & ((en[1] $ (\ramREN~0_combout )) # (!\ramWEN~0_combout ))) # (!en[0] & ((\ramWEN~0_combout ) # (en[1] $ (\ramREN~0_combout ))))

	.dataa(en[0]),
	.datab(en[1]),
	.datac(ramREN),
	.datad(ramWEN),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'h7DBE;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N0
cycloneive_lcell_comb \always0~1 (
// Equation(s):
// \always0~1_combout  = (always1) # ((\always0~0_combout ) # (!\Equal2~20_combout ))

	.dataa(always1),
	.datab(\always0~0_combout ),
	.datac(gnd),
	.datad(\Equal2~20_combout ),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
// synopsys translate_off
defparam \always0~1 .lut_mask = 16'hEEFF;
defparam \always0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N23
dffeas \addr[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr9),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[8]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[8] .is_wysiwyg = "true";
defparam \addr[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N22
cycloneive_lcell_comb \Equal2~5 (
// Equation(s):
// \Equal2~5_combout  = (addr[9] & (\ramaddr~17_combout  & (addr[8] $ (!\ramaddr~19_combout )))) # (!addr[9] & (!\ramaddr~17_combout  & (addr[8] $ (!\ramaddr~19_combout ))))

	.dataa(addr[9]),
	.datab(ramaddr8),
	.datac(addr[8]),
	.datad(ramaddr9),
	.cin(gnd),
	.combout(\Equal2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~5 .lut_mask = 16'h9009;
defparam \Equal2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y31_N11
dffeas \addr[13] (
	.clk(CLK),
	.d(ramaddr12),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[13]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[13] .is_wysiwyg = "true";
defparam \addr[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N25
dffeas \addr[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr13),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[12]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[12] .is_wysiwyg = "true";
defparam \addr[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N24
cycloneive_lcell_comb \Equal2~7 (
// Equation(s):
// \Equal2~7_combout  = (\ramaddr~25_combout  & (addr[13] & (addr[12] $ (!\ramaddr~27_combout )))) # (!\ramaddr~25_combout  & (!addr[13] & (addr[12] $ (!\ramaddr~27_combout ))))

	.dataa(ramaddr12),
	.datab(addr[13]),
	.datac(addr[12]),
	.datad(ramaddr13),
	.cin(gnd),
	.combout(\Equal2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~7 .lut_mask = 16'h9009;
defparam \Equal2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N13
dffeas \addr[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr11),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[10]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[10] .is_wysiwyg = "true";
defparam \addr[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N12
cycloneive_lcell_comb \Equal2~6 (
// Equation(s):
// \Equal2~6_combout  = (addr[11] & (\ramaddr~21_combout  & (addr[10] $ (!\ramaddr~23_combout )))) # (!addr[11] & (!\ramaddr~21_combout  & (addr[10] $ (!\ramaddr~23_combout ))))

	.dataa(addr[11]),
	.datab(ramaddr10),
	.datac(addr[10]),
	.datad(ramaddr11),
	.cin(gnd),
	.combout(\Equal2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~6 .lut_mask = 16'h9009;
defparam \Equal2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N22
cycloneive_lcell_comb \Equal2~9 (
// Equation(s):
// \Equal2~9_combout  = (\Equal2~8_combout  & (\Equal2~5_combout  & (\Equal2~7_combout  & \Equal2~6_combout )))

	.dataa(\Equal2~8_combout ),
	.datab(\Equal2~5_combout ),
	.datac(\Equal2~7_combout ),
	.datad(\Equal2~6_combout ),
	.cin(gnd),
	.combout(\Equal2~9_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~9 .lut_mask = 16'h8000;
defparam \Equal2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y32_N7
dffeas \addr[25] (
	.clk(CLK),
	.d(\ramif.ramaddr [25]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[25]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[25] .is_wysiwyg = "true";
defparam \addr[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y32_N25
dffeas \addr[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr22),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[24]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[24] .is_wysiwyg = "true";
defparam \addr[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N24
cycloneive_lcell_comb \Equal2~15 (
// Equation(s):
// \Equal2~15_combout  = (\ramaddr~49_combout  & (addr[25] & (addr[24] $ (!\ramaddr~51_combout )))) # (!\ramaddr~49_combout  & (!addr[25] & (addr[24] $ (!\ramaddr~51_combout ))))

	.dataa(\ramif.ramaddr [25]),
	.datab(addr[25]),
	.datac(addr[24]),
	.datad(ramaddr22),
	.cin(gnd),
	.combout(\Equal2~15_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~15 .lut_mask = 16'h9009;
defparam \Equal2~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y32_N5
dffeas \addr[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr23),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[26]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[26] .is_wysiwyg = "true";
defparam \addr[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N4
cycloneive_lcell_comb \Equal2~16 (
// Equation(s):
// \Equal2~16_combout  = (addr[27] & (\ramaddr~53_combout  & (\ramaddr~55_combout  $ (!addr[26])))) # (!addr[27] & (!\ramaddr~53_combout  & (\ramaddr~55_combout  $ (!addr[26]))))

	.dataa(addr[27]),
	.datab(ramaddr23),
	.datac(addr[26]),
	.datad(\ramif.ramaddr [27]),
	.cin(gnd),
	.combout(\Equal2~16_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~16 .lut_mask = 16'h8241;
defparam \Equal2~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y32_N11
dffeas \addr[30] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr26),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[30]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[30] .is_wysiwyg = "true";
defparam \addr[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N10
cycloneive_lcell_comb \Equal2~18 (
// Equation(s):
// \Equal2~18_combout  = (addr[31] & (\ramaddr~61_combout  & (\ramaddr~63_combout  $ (!addr[30])))) # (!addr[31] & (!\ramaddr~61_combout  & (\ramaddr~63_combout  $ (!addr[30]))))

	.dataa(addr[31]),
	.datab(ramaddr26),
	.datac(addr[30]),
	.datad(ramaddr25),
	.cin(gnd),
	.combout(\Equal2~18_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~18 .lut_mask = 16'h8241;
defparam \Equal2~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N16
cycloneive_lcell_comb \Equal2~19 (
// Equation(s):
// \Equal2~19_combout  = (\Equal2~17_combout  & (\Equal2~15_combout  & (\Equal2~16_combout  & \Equal2~18_combout )))

	.dataa(\Equal2~17_combout ),
	.datab(\Equal2~15_combout ),
	.datac(\Equal2~16_combout ),
	.datad(\Equal2~18_combout ),
	.cin(gnd),
	.combout(\Equal2~19_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~19 .lut_mask = 16'h8000;
defparam \Equal2~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y32_N11
dffeas \addr[23] (
	.clk(CLK),
	.d(\ramif.ramaddr [23]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[23]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[23] .is_wysiwyg = "true";
defparam \addr[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N29
dffeas \addr[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr21),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[22]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[22] .is_wysiwyg = "true";
defparam \addr[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N28
cycloneive_lcell_comb \Equal2~13 (
// Equation(s):
// \Equal2~13_combout  = (\ramaddr~45_combout  & (addr[23] & (addr[22] $ (!\ramaddr~47_combout )))) # (!\ramaddr~45_combout  & (!addr[23] & (addr[22] $ (!\ramaddr~47_combout ))))

	.dataa(\ramif.ramaddr [23]),
	.datab(addr[23]),
	.datac(addr[22]),
	.datad(ramaddr21),
	.cin(gnd),
	.combout(\Equal2~13_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~13 .lut_mask = 16'h9009;
defparam \Equal2~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y32_N9
dffeas \addr[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr20),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[20]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[20] .is_wysiwyg = "true";
defparam \addr[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N8
cycloneive_lcell_comb \Equal2~12 (
// Equation(s):
// \Equal2~12_combout  = (addr[21] & (\ramaddr~41_combout  & (\ramaddr~43_combout  $ (!addr[20])))) # (!addr[21] & (!\ramaddr~41_combout  & (\ramaddr~43_combout  $ (!addr[20]))))

	.dataa(addr[21]),
	.datab(ramaddr20),
	.datac(addr[20]),
	.datad(ramaddr19),
	.cin(gnd),
	.combout(\Equal2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~12 .lut_mask = 16'h8241;
defparam \Equal2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y32_N5
dffeas \addr[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr17),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[19]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[19] .is_wysiwyg = "true";
defparam \addr[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y32_N25
dffeas \addr[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr18),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[18]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[18] .is_wysiwyg = "true";
defparam \addr[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N24
cycloneive_lcell_comb \Equal2~11 (
// Equation(s):
// \Equal2~11_combout  = (\ramaddr~37_combout  & (addr[19] & (addr[18] $ (!\ramaddr~39_combout )))) # (!\ramaddr~37_combout  & (!addr[19] & (addr[18] $ (!\ramaddr~39_combout ))))

	.dataa(ramaddr17),
	.datab(addr[19]),
	.datac(addr[18]),
	.datad(ramaddr18),
	.cin(gnd),
	.combout(\Equal2~11_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~11 .lut_mask = 16'h9009;
defparam \Equal2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N4
cycloneive_lcell_comb \Equal2~14 (
// Equation(s):
// \Equal2~14_combout  = (\Equal2~10_combout  & (\Equal2~13_combout  & (\Equal2~12_combout  & \Equal2~11_combout )))

	.dataa(\Equal2~10_combout ),
	.datab(\Equal2~13_combout ),
	.datac(\Equal2~12_combout ),
	.datad(\Equal2~11_combout ),
	.cin(gnd),
	.combout(\Equal2~14_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~14 .lut_mask = 16'h8000;
defparam \Equal2~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y32_N15
dffeas \addr[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr2),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[3]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[3] .is_wysiwyg = "true";
defparam \addr[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N21
dffeas \addr[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr3),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[2]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[2] .is_wysiwyg = "true";
defparam \addr[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N20
cycloneive_lcell_comb \Equal2~1 (
// Equation(s):
// \Equal2~1_combout  = (\ramaddr~7_combout  & (addr[2] & (addr[3] $ (!\ramaddr~5_combout )))) # (!\ramaddr~7_combout  & (!addr[2] & (addr[3] $ (!\ramaddr~5_combout ))))

	.dataa(ramaddr3),
	.datab(addr[3]),
	.datac(addr[2]),
	.datad(ramaddr2),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~1 .lut_mask = 16'h8421;
defparam \Equal2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N9
dffeas \addr[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr1),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[0]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[0] .is_wysiwyg = "true";
defparam \addr[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N8
cycloneive_lcell_comb \Equal2~0 (
// Equation(s):
// \Equal2~0_combout  = (addr[1] & (\ramaddr~1_combout  & (addr[0] $ (!\ramaddr~3_combout )))) # (!addr[1] & (!\ramaddr~1_combout  & (addr[0] $ (!\ramaddr~3_combout ))))

	.dataa(addr[1]),
	.datab(ramaddr),
	.datac(addr[0]),
	.datad(ramaddr1),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~0 .lut_mask = 16'h9009;
defparam \Equal2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y28_N25
dffeas \addr[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr5),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[4]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[4] .is_wysiwyg = "true";
defparam \addr[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N24
cycloneive_lcell_comb \Equal2~2 (
// Equation(s):
// \Equal2~2_combout  = (addr[5] & (\ramaddr~9_combout  & (\ramaddr~11_combout  $ (!addr[4])))) # (!addr[5] & (!\ramaddr~9_combout  & (\ramaddr~11_combout  $ (!addr[4]))))

	.dataa(addr[5]),
	.datab(ramaddr5),
	.datac(addr[4]),
	.datad(ramaddr4),
	.cin(gnd),
	.combout(\Equal2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~2 .lut_mask = 16'h8241;
defparam \Equal2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N28
cycloneive_lcell_comb \Equal2~4 (
// Equation(s):
// \Equal2~4_combout  = (\Equal2~3_combout  & (\Equal2~1_combout  & (\Equal2~0_combout  & \Equal2~2_combout )))

	.dataa(\Equal2~3_combout ),
	.datab(\Equal2~1_combout ),
	.datac(\Equal2~0_combout ),
	.datad(\Equal2~2_combout ),
	.cin(gnd),
	.combout(\Equal2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~4 .lut_mask = 16'h8000;
defparam \Equal2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N6
cycloneive_lcell_comb \Equal2~20 (
// Equation(s):
// \Equal2~20_combout  = (\Equal2~9_combout  & (\Equal2~19_combout  & (\Equal2~14_combout  & \Equal2~4_combout )))

	.dataa(\Equal2~9_combout ),
	.datab(\Equal2~19_combout ),
	.datac(\Equal2~14_combout ),
	.datad(\Equal2~4_combout ),
	.cin(gnd),
	.combout(\Equal2~20_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~20 .lut_mask = 16'h8000;
defparam \Equal2~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N10
cycloneive_lcell_comb \ramif.ramload[0]~1 (
// Equation(s):
// \ramif.ramload[0]~1_combout  = (!\syif.WEN~input_o  & (\syif.tbCTRL~input_o  & !\syif.REN~input_o ))

	.dataa(gnd),
	.datab(syifWEN),
	.datac(syiftbCTRL),
	.datad(syifREN),
	.cin(gnd),
	.combout(\ramif.ramload[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[0]~1 .lut_mask = 16'h0030;
defparam \ramif.ramload[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N6
cycloneive_lcell_comb \ramif.ramload[1]~4 (
// Equation(s):
// \ramif.ramload[1]~4_combout  = (\syif.WEN~input_o ) # ((\syif.REN~input_o ) # (!\syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(syifWEN),
	.datac(syiftbCTRL),
	.datad(syifREN),
	.cin(gnd),
	.combout(\ramif.ramload[1]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[1]~4 .lut_mask = 16'hFFCF;
defparam \ramif.ramload[1]~4 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module altsyncram_1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	ramWEN,
	data_a,
	ramaddr1,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	ramWEN;
input 	[31:0] data_a;
input 	ramaddr1;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



altsyncram_99f1 auto_generated(
	.ram_block3a32(ram_block3a32),
	.ram_block3a0(ram_block3a0),
	.ram_block3a33(ram_block3a33),
	.ram_block3a1(ram_block3a1),
	.ram_block3a34(ram_block3a34),
	.ram_block3a2(ram_block3a2),
	.ram_block3a35(ram_block3a35),
	.ram_block3a3(ram_block3a3),
	.ram_block3a36(ram_block3a36),
	.ram_block3a4(ram_block3a4),
	.ram_block3a37(ram_block3a37),
	.ram_block3a5(ram_block3a5),
	.ram_block3a38(ram_block3a38),
	.ram_block3a6(ram_block3a6),
	.ram_block3a39(ram_block3a39),
	.ram_block3a7(ram_block3a7),
	.ram_block3a40(ram_block3a40),
	.ram_block3a8(ram_block3a8),
	.ram_block3a41(ram_block3a41),
	.ram_block3a9(ram_block3a9),
	.ram_block3a42(ram_block3a42),
	.ram_block3a10(ram_block3a10),
	.ram_block3a43(ram_block3a43),
	.ram_block3a11(ram_block3a11),
	.ram_block3a44(ram_block3a44),
	.ram_block3a12(ram_block3a12),
	.ram_block3a45(ram_block3a45),
	.ram_block3a13(ram_block3a13),
	.ram_block3a46(ram_block3a46),
	.ram_block3a14(ram_block3a14),
	.ram_block3a47(ram_block3a47),
	.ram_block3a15(ram_block3a15),
	.ram_block3a48(ram_block3a48),
	.ram_block3a16(ram_block3a16),
	.ram_block3a49(ram_block3a49),
	.ram_block3a17(ram_block3a17),
	.ram_block3a50(ram_block3a50),
	.ram_block3a18(ram_block3a18),
	.ram_block3a51(ram_block3a51),
	.ram_block3a19(ram_block3a19),
	.ram_block3a52(ram_block3a52),
	.ram_block3a20(ram_block3a20),
	.ram_block3a53(ram_block3a53),
	.ram_block3a21(ram_block3a21),
	.ram_block3a54(ram_block3a54),
	.ram_block3a22(ram_block3a22),
	.ram_block3a55(ram_block3a55),
	.ram_block3a23(ram_block3a23),
	.ram_block3a56(ram_block3a56),
	.ram_block3a24(ram_block3a24),
	.ram_block3a57(ram_block3a57),
	.ram_block3a25(ram_block3a25),
	.ram_block3a58(ram_block3a58),
	.ram_block3a26(ram_block3a26),
	.ram_block3a59(ram_block3a59),
	.ram_block3a27(ram_block3a27),
	.ram_block3a60(ram_block3a60),
	.ram_block3a28(ram_block3a28),
	.ram_block3a61(ram_block3a61),
	.ram_block3a29(ram_block3a29),
	.ram_block3a62(ram_block3a62),
	.ram_block3a30(ram_block3a30),
	.ram_block3a63(ram_block3a63),
	.ram_block3a31(ram_block3a31),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(address_reg_a_0),
	.address_a({gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.ramWEN(ramWEN),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.ramaddr1(ramaddr1),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_99f1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	ramWEN,
	data_a,
	ramaddr1,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	ramWEN;
input 	[31:0] data_a;
input 	ramaddr1;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram1|ram_block3a32~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a0~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a33~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a1~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a34~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a2~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a35~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a3~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a36~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a4~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a37~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a5~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a38~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a6~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a39~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a7~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a40~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a8~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a41~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a9~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a42~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a10~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a43~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a11~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a44~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a12~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a45~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a13~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a46~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a14~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a47~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a15~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a48~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a16~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a49~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a17~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a50~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a18~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a51~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a19~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a52~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a20~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a53~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a21~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a54~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a22~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a55~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a23~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a56~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a24~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a57~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a25~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a58~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a26~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a59~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a27~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a60~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a28~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a61~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a29~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a62~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a30~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a63~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a31~PORTBDATAOUT0 ;
wire \mgl_prim2|sdr~0_combout ;
wire [0:0] \altsyncram1|address_reg_b ;
wire [31:0] \mgl_prim2|ram_rom_data_reg ;
wire [13:0] \mgl_prim2|ram_rom_addr_reg ;


sld_mod_ram_rom mgl_prim2(
	.ram_block3a32(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a0(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a33(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a1(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a34(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a2(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a35(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a3(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a36(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a4(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a37(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a5(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a38(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a6(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a39(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a7(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a40(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a8(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a41(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a9(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a42(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a10(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a43(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a11(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a44(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a12(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a45(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a13(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a46(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a14(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a47(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a15(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a48(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a16(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a49(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a17(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a50(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a18(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a51(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a19(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a52(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a20(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a53(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a21(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a54(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a22(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a55(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a23(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a56(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a24(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a57(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a25(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a58(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a26(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a59(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a27(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a60(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a28(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a61(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a29(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a62(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a30(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a63(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a31(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.is_in_use_reg1(is_in_use_reg),
	.ram_rom_data_reg_0(\mgl_prim2|ram_rom_data_reg [0]),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.ram_rom_addr_reg_0(\mgl_prim2|ram_rom_addr_reg [0]),
	.ram_rom_addr_reg_1(\mgl_prim2|ram_rom_addr_reg [1]),
	.ram_rom_addr_reg_2(\mgl_prim2|ram_rom_addr_reg [2]),
	.ram_rom_addr_reg_3(\mgl_prim2|ram_rom_addr_reg [3]),
	.ram_rom_addr_reg_4(\mgl_prim2|ram_rom_addr_reg [4]),
	.ram_rom_addr_reg_5(\mgl_prim2|ram_rom_addr_reg [5]),
	.ram_rom_addr_reg_6(\mgl_prim2|ram_rom_addr_reg [6]),
	.ram_rom_addr_reg_7(\mgl_prim2|ram_rom_addr_reg [7]),
	.ram_rom_addr_reg_8(\mgl_prim2|ram_rom_addr_reg [8]),
	.ram_rom_addr_reg_9(\mgl_prim2|ram_rom_addr_reg [9]),
	.ram_rom_addr_reg_10(\mgl_prim2|ram_rom_addr_reg [10]),
	.ram_rom_addr_reg_11(\mgl_prim2|ram_rom_addr_reg [11]),
	.ram_rom_addr_reg_12(\mgl_prim2|ram_rom_addr_reg [12]),
	.ram_rom_data_reg_1(\mgl_prim2|ram_rom_data_reg [1]),
	.ram_rom_data_reg_2(\mgl_prim2|ram_rom_data_reg [2]),
	.ram_rom_data_reg_3(\mgl_prim2|ram_rom_data_reg [3]),
	.ram_rom_data_reg_4(\mgl_prim2|ram_rom_data_reg [4]),
	.ram_rom_data_reg_5(\mgl_prim2|ram_rom_data_reg [5]),
	.ram_rom_data_reg_6(\mgl_prim2|ram_rom_data_reg [6]),
	.ram_rom_data_reg_7(\mgl_prim2|ram_rom_data_reg [7]),
	.ram_rom_data_reg_8(\mgl_prim2|ram_rom_data_reg [8]),
	.ram_rom_data_reg_9(\mgl_prim2|ram_rom_data_reg [9]),
	.ram_rom_data_reg_10(\mgl_prim2|ram_rom_data_reg [10]),
	.ram_rom_data_reg_11(\mgl_prim2|ram_rom_data_reg [11]),
	.ram_rom_data_reg_12(\mgl_prim2|ram_rom_data_reg [12]),
	.ram_rom_data_reg_13(\mgl_prim2|ram_rom_data_reg [13]),
	.ram_rom_data_reg_14(\mgl_prim2|ram_rom_data_reg [14]),
	.ram_rom_data_reg_15(\mgl_prim2|ram_rom_data_reg [15]),
	.ram_rom_data_reg_16(\mgl_prim2|ram_rom_data_reg [16]),
	.ram_rom_data_reg_17(\mgl_prim2|ram_rom_data_reg [17]),
	.ram_rom_data_reg_18(\mgl_prim2|ram_rom_data_reg [18]),
	.ram_rom_data_reg_19(\mgl_prim2|ram_rom_data_reg [19]),
	.ram_rom_data_reg_20(\mgl_prim2|ram_rom_data_reg [20]),
	.ram_rom_data_reg_21(\mgl_prim2|ram_rom_data_reg [21]),
	.ram_rom_data_reg_22(\mgl_prim2|ram_rom_data_reg [22]),
	.ram_rom_data_reg_23(\mgl_prim2|ram_rom_data_reg [23]),
	.ram_rom_data_reg_24(\mgl_prim2|ram_rom_data_reg [24]),
	.ram_rom_data_reg_25(\mgl_prim2|ram_rom_data_reg [25]),
	.ram_rom_data_reg_26(\mgl_prim2|ram_rom_data_reg [26]),
	.ram_rom_data_reg_27(\mgl_prim2|ram_rom_data_reg [27]),
	.ram_rom_data_reg_28(\mgl_prim2|ram_rom_data_reg [28]),
	.ram_rom_data_reg_29(\mgl_prim2|ram_rom_data_reg [29]),
	.ram_rom_data_reg_30(\mgl_prim2|ram_rom_data_reg [30]),
	.ram_rom_data_reg_31(\mgl_prim2|ram_rom_data_reg [31]),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.ir_in({gnd,irf_reg_3_1,gnd,gnd,irf_reg_0_1}),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.raw_tck(altera_internal_jtag1),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

altsyncram_fta2 altsyncram1(
	.ram_block3a321(ram_block3a32),
	.ram_block3a322(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a01(ram_block3a0),
	.ram_block3a02(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a331(ram_block3a33),
	.ram_block3a332(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a110(ram_block3a1),
	.ram_block3a111(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a341(ram_block3a34),
	.ram_block3a342(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a210(ram_block3a2),
	.ram_block3a211(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a351(ram_block3a35),
	.ram_block3a352(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a310(ram_block3a3),
	.ram_block3a311(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a361(ram_block3a36),
	.ram_block3a362(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a410(ram_block3a4),
	.ram_block3a411(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a371(ram_block3a37),
	.ram_block3a372(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a510(ram_block3a5),
	.ram_block3a511(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a381(ram_block3a38),
	.ram_block3a382(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a64(ram_block3a6),
	.ram_block3a65(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a391(ram_block3a39),
	.ram_block3a392(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a71(ram_block3a7),
	.ram_block3a72(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a401(ram_block3a40),
	.ram_block3a402(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a81(ram_block3a8),
	.ram_block3a82(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a412(ram_block3a41),
	.ram_block3a413(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a91(ram_block3a9),
	.ram_block3a92(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a421(ram_block3a42),
	.ram_block3a422(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a101(ram_block3a10),
	.ram_block3a102(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a431(ram_block3a43),
	.ram_block3a432(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a112(ram_block3a11),
	.ram_block3a113(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a441(ram_block3a44),
	.ram_block3a442(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a121(ram_block3a12),
	.ram_block3a122(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a451(ram_block3a45),
	.ram_block3a452(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a131(ram_block3a13),
	.ram_block3a132(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a461(ram_block3a46),
	.ram_block3a462(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a141(ram_block3a14),
	.ram_block3a142(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a471(ram_block3a47),
	.ram_block3a472(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a151(ram_block3a15),
	.ram_block3a152(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a481(ram_block3a48),
	.ram_block3a482(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a161(ram_block3a16),
	.ram_block3a162(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a491(ram_block3a49),
	.ram_block3a492(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a171(ram_block3a17),
	.ram_block3a172(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a501(ram_block3a50),
	.ram_block3a502(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a181(ram_block3a18),
	.ram_block3a182(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a512(ram_block3a51),
	.ram_block3a513(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a191(ram_block3a19),
	.ram_block3a192(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a521(ram_block3a52),
	.ram_block3a522(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a201(ram_block3a20),
	.ram_block3a202(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a531(ram_block3a53),
	.ram_block3a532(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a212(ram_block3a21),
	.ram_block3a213(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a541(ram_block3a54),
	.ram_block3a542(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a221(ram_block3a22),
	.ram_block3a222(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a551(ram_block3a55),
	.ram_block3a552(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a231(ram_block3a23),
	.ram_block3a232(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a561(ram_block3a56),
	.ram_block3a562(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a241(ram_block3a24),
	.ram_block3a242(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a571(ram_block3a57),
	.ram_block3a572(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a251(ram_block3a25),
	.ram_block3a252(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a581(ram_block3a58),
	.ram_block3a582(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a261(ram_block3a26),
	.ram_block3a262(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a591(ram_block3a59),
	.ram_block3a592(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a271(ram_block3a27),
	.ram_block3a272(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a601(ram_block3a60),
	.ram_block3a602(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a281(ram_block3a28),
	.ram_block3a282(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a611(ram_block3a61),
	.ram_block3a612(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a291(ram_block3a29),
	.ram_block3a292(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a621(ram_block3a62),
	.ram_block3a622(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a301(ram_block3a30),
	.ram_block3a302(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a631(ram_block3a63),
	.ram_block3a632(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a312(ram_block3a31),
	.ram_block3a313(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.data_b({\mgl_prim2|ram_rom_data_reg [31],\mgl_prim2|ram_rom_data_reg [30],\mgl_prim2|ram_rom_data_reg [29],\mgl_prim2|ram_rom_data_reg [28],\mgl_prim2|ram_rom_data_reg [27],\mgl_prim2|ram_rom_data_reg [26],\mgl_prim2|ram_rom_data_reg [25],\mgl_prim2|ram_rom_data_reg [24],\mgl_prim2|ram_rom_data_reg [23],
\mgl_prim2|ram_rom_data_reg [22],\mgl_prim2|ram_rom_data_reg [21],\mgl_prim2|ram_rom_data_reg [20],\mgl_prim2|ram_rom_data_reg [19],\mgl_prim2|ram_rom_data_reg [18],\mgl_prim2|ram_rom_data_reg [17],\mgl_prim2|ram_rom_data_reg [16],\mgl_prim2|ram_rom_data_reg [15],\mgl_prim2|ram_rom_data_reg [14],
\mgl_prim2|ram_rom_data_reg [13],\mgl_prim2|ram_rom_data_reg [12],\mgl_prim2|ram_rom_data_reg [11],\mgl_prim2|ram_rom_data_reg [10],\mgl_prim2|ram_rom_data_reg [9],\mgl_prim2|ram_rom_data_reg [8],\mgl_prim2|ram_rom_data_reg [7],\mgl_prim2|ram_rom_data_reg [6],\mgl_prim2|ram_rom_data_reg [5],
\mgl_prim2|ram_rom_data_reg [4],\mgl_prim2|ram_rom_data_reg [3],\mgl_prim2|ram_rom_data_reg [2],\mgl_prim2|ram_rom_data_reg [1],\mgl_prim2|ram_rom_data_reg [0]}),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.address_b({gnd,\mgl_prim2|ram_rom_addr_reg [12],\mgl_prim2|ram_rom_addr_reg [11],\mgl_prim2|ram_rom_addr_reg [10],\mgl_prim2|ram_rom_addr_reg [9],\mgl_prim2|ram_rom_addr_reg [8],\mgl_prim2|ram_rom_addr_reg [7],\mgl_prim2|ram_rom_addr_reg [6],\mgl_prim2|ram_rom_addr_reg [5],\mgl_prim2|ram_rom_addr_reg [4],
\mgl_prim2|ram_rom_addr_reg [3],\mgl_prim2|ram_rom_addr_reg [2],\mgl_prim2|ram_rom_addr_reg [1],\mgl_prim2|ram_rom_addr_reg [0]}),
	.address_reg_a_0(address_reg_a_0),
	.address_a({gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.always1(always1),
	.ramWEN(ramWEN),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.ramaddr1(ramaddr1),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.clock1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_fta2 (
	ram_block3a321,
	ram_block3a322,
	ram_block3a01,
	ram_block3a02,
	ram_block3a331,
	ram_block3a332,
	ram_block3a110,
	ram_block3a111,
	ram_block3a341,
	ram_block3a342,
	ram_block3a210,
	ram_block3a211,
	ram_block3a351,
	ram_block3a352,
	ram_block3a310,
	ram_block3a311,
	ram_block3a361,
	ram_block3a362,
	ram_block3a410,
	ram_block3a411,
	ram_block3a371,
	ram_block3a372,
	ram_block3a510,
	ram_block3a511,
	ram_block3a381,
	ram_block3a382,
	ram_block3a64,
	ram_block3a65,
	ram_block3a391,
	ram_block3a392,
	ram_block3a71,
	ram_block3a72,
	ram_block3a401,
	ram_block3a402,
	ram_block3a81,
	ram_block3a82,
	ram_block3a412,
	ram_block3a413,
	ram_block3a91,
	ram_block3a92,
	ram_block3a421,
	ram_block3a422,
	ram_block3a101,
	ram_block3a102,
	ram_block3a431,
	ram_block3a432,
	ram_block3a112,
	ram_block3a113,
	ram_block3a441,
	ram_block3a442,
	ram_block3a121,
	ram_block3a122,
	ram_block3a451,
	ram_block3a452,
	ram_block3a131,
	ram_block3a132,
	ram_block3a461,
	ram_block3a462,
	ram_block3a141,
	ram_block3a142,
	ram_block3a471,
	ram_block3a472,
	ram_block3a151,
	ram_block3a152,
	ram_block3a481,
	ram_block3a482,
	ram_block3a161,
	ram_block3a162,
	ram_block3a491,
	ram_block3a492,
	ram_block3a171,
	ram_block3a172,
	ram_block3a501,
	ram_block3a502,
	ram_block3a181,
	ram_block3a182,
	ram_block3a512,
	ram_block3a513,
	ram_block3a191,
	ram_block3a192,
	ram_block3a521,
	ram_block3a522,
	ram_block3a201,
	ram_block3a202,
	ram_block3a531,
	ram_block3a532,
	ram_block3a212,
	ram_block3a213,
	ram_block3a541,
	ram_block3a542,
	ram_block3a221,
	ram_block3a222,
	ram_block3a551,
	ram_block3a552,
	ram_block3a231,
	ram_block3a232,
	ram_block3a561,
	ram_block3a562,
	ram_block3a241,
	ram_block3a242,
	ram_block3a571,
	ram_block3a572,
	ram_block3a251,
	ram_block3a252,
	ram_block3a581,
	ram_block3a582,
	ram_block3a261,
	ram_block3a262,
	ram_block3a591,
	ram_block3a592,
	ram_block3a271,
	ram_block3a272,
	ram_block3a601,
	ram_block3a602,
	ram_block3a281,
	ram_block3a282,
	ram_block3a611,
	ram_block3a612,
	ram_block3a291,
	ram_block3a292,
	ram_block3a621,
	ram_block3a622,
	ram_block3a301,
	ram_block3a302,
	ram_block3a631,
	ram_block3a632,
	ram_block3a312,
	ram_block3a313,
	data_b,
	ram_rom_addr_reg_13,
	address_b,
	address_reg_a_0,
	address_a,
	ramaddr,
	always1,
	ramWEN,
	sdr,
	data_a,
	address_reg_b_0,
	ramaddr1,
	irf_reg_2_1,
	state_5,
	clock1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a321;
output 	ram_block3a322;
output 	ram_block3a01;
output 	ram_block3a02;
output 	ram_block3a331;
output 	ram_block3a332;
output 	ram_block3a110;
output 	ram_block3a111;
output 	ram_block3a341;
output 	ram_block3a342;
output 	ram_block3a210;
output 	ram_block3a211;
output 	ram_block3a351;
output 	ram_block3a352;
output 	ram_block3a310;
output 	ram_block3a311;
output 	ram_block3a361;
output 	ram_block3a362;
output 	ram_block3a410;
output 	ram_block3a411;
output 	ram_block3a371;
output 	ram_block3a372;
output 	ram_block3a510;
output 	ram_block3a511;
output 	ram_block3a381;
output 	ram_block3a382;
output 	ram_block3a64;
output 	ram_block3a65;
output 	ram_block3a391;
output 	ram_block3a392;
output 	ram_block3a71;
output 	ram_block3a72;
output 	ram_block3a401;
output 	ram_block3a402;
output 	ram_block3a81;
output 	ram_block3a82;
output 	ram_block3a412;
output 	ram_block3a413;
output 	ram_block3a91;
output 	ram_block3a92;
output 	ram_block3a421;
output 	ram_block3a422;
output 	ram_block3a101;
output 	ram_block3a102;
output 	ram_block3a431;
output 	ram_block3a432;
output 	ram_block3a112;
output 	ram_block3a113;
output 	ram_block3a441;
output 	ram_block3a442;
output 	ram_block3a121;
output 	ram_block3a122;
output 	ram_block3a451;
output 	ram_block3a452;
output 	ram_block3a131;
output 	ram_block3a132;
output 	ram_block3a461;
output 	ram_block3a462;
output 	ram_block3a141;
output 	ram_block3a142;
output 	ram_block3a471;
output 	ram_block3a472;
output 	ram_block3a151;
output 	ram_block3a152;
output 	ram_block3a481;
output 	ram_block3a482;
output 	ram_block3a161;
output 	ram_block3a162;
output 	ram_block3a491;
output 	ram_block3a492;
output 	ram_block3a171;
output 	ram_block3a172;
output 	ram_block3a501;
output 	ram_block3a502;
output 	ram_block3a181;
output 	ram_block3a182;
output 	ram_block3a512;
output 	ram_block3a513;
output 	ram_block3a191;
output 	ram_block3a192;
output 	ram_block3a521;
output 	ram_block3a522;
output 	ram_block3a201;
output 	ram_block3a202;
output 	ram_block3a531;
output 	ram_block3a532;
output 	ram_block3a212;
output 	ram_block3a213;
output 	ram_block3a541;
output 	ram_block3a542;
output 	ram_block3a221;
output 	ram_block3a222;
output 	ram_block3a551;
output 	ram_block3a552;
output 	ram_block3a231;
output 	ram_block3a232;
output 	ram_block3a561;
output 	ram_block3a562;
output 	ram_block3a241;
output 	ram_block3a242;
output 	ram_block3a571;
output 	ram_block3a572;
output 	ram_block3a251;
output 	ram_block3a252;
output 	ram_block3a581;
output 	ram_block3a582;
output 	ram_block3a261;
output 	ram_block3a262;
output 	ram_block3a591;
output 	ram_block3a592;
output 	ram_block3a271;
output 	ram_block3a272;
output 	ram_block3a601;
output 	ram_block3a602;
output 	ram_block3a281;
output 	ram_block3a282;
output 	ram_block3a611;
output 	ram_block3a612;
output 	ram_block3a291;
output 	ram_block3a292;
output 	ram_block3a621;
output 	ram_block3a622;
output 	ram_block3a301;
output 	ram_block3a302;
output 	ram_block3a631;
output 	ram_block3a632;
output 	ram_block3a312;
output 	ram_block3a313;
input 	[31:0] data_b;
input 	ram_rom_addr_reg_13;
input 	[13:0] address_b;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	always1;
input 	ramWEN;
input 	sdr;
input 	[31:0] data_a;
output 	address_reg_b_0;
input 	ramaddr1;
input 	irf_reg_2_1;
input 	state_5;
input 	clock1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \decode4|eq_node[1]~0_combout ;
wire \decode5|eq_node[1]~0_combout ;
wire \decode4|eq_node[0]~1_combout ;
wire \decode5|eq_node[0]~1_combout ;
wire \address_reg_b[0]~feeder_combout ;

wire [0:0] ram_block3a32_PORTADATAOUT_bus;
wire [0:0] ram_block3a32_PORTBDATAOUT_bus;
wire [0:0] ram_block3a0_PORTADATAOUT_bus;
wire [0:0] ram_block3a0_PORTBDATAOUT_bus;
wire [0:0] ram_block3a33_PORTADATAOUT_bus;
wire [0:0] ram_block3a33_PORTBDATAOUT_bus;
wire [0:0] ram_block3a1_PORTADATAOUT_bus;
wire [0:0] ram_block3a1_PORTBDATAOUT_bus;
wire [0:0] ram_block3a34_PORTADATAOUT_bus;
wire [0:0] ram_block3a34_PORTBDATAOUT_bus;
wire [0:0] ram_block3a2_PORTADATAOUT_bus;
wire [0:0] ram_block3a2_PORTBDATAOUT_bus;
wire [0:0] ram_block3a35_PORTADATAOUT_bus;
wire [0:0] ram_block3a35_PORTBDATAOUT_bus;
wire [0:0] ram_block3a3_PORTADATAOUT_bus;
wire [0:0] ram_block3a3_PORTBDATAOUT_bus;
wire [0:0] ram_block3a36_PORTADATAOUT_bus;
wire [0:0] ram_block3a36_PORTBDATAOUT_bus;
wire [0:0] ram_block3a4_PORTADATAOUT_bus;
wire [0:0] ram_block3a4_PORTBDATAOUT_bus;
wire [0:0] ram_block3a37_PORTADATAOUT_bus;
wire [0:0] ram_block3a37_PORTBDATAOUT_bus;
wire [0:0] ram_block3a5_PORTADATAOUT_bus;
wire [0:0] ram_block3a5_PORTBDATAOUT_bus;
wire [0:0] ram_block3a38_PORTADATAOUT_bus;
wire [0:0] ram_block3a38_PORTBDATAOUT_bus;
wire [0:0] ram_block3a6_PORTADATAOUT_bus;
wire [0:0] ram_block3a6_PORTBDATAOUT_bus;
wire [0:0] ram_block3a39_PORTADATAOUT_bus;
wire [0:0] ram_block3a39_PORTBDATAOUT_bus;
wire [0:0] ram_block3a7_PORTADATAOUT_bus;
wire [0:0] ram_block3a7_PORTBDATAOUT_bus;
wire [0:0] ram_block3a40_PORTADATAOUT_bus;
wire [0:0] ram_block3a40_PORTBDATAOUT_bus;
wire [0:0] ram_block3a8_PORTADATAOUT_bus;
wire [0:0] ram_block3a8_PORTBDATAOUT_bus;
wire [0:0] ram_block3a41_PORTADATAOUT_bus;
wire [0:0] ram_block3a41_PORTBDATAOUT_bus;
wire [0:0] ram_block3a9_PORTADATAOUT_bus;
wire [0:0] ram_block3a9_PORTBDATAOUT_bus;
wire [0:0] ram_block3a42_PORTADATAOUT_bus;
wire [0:0] ram_block3a42_PORTBDATAOUT_bus;
wire [0:0] ram_block3a10_PORTADATAOUT_bus;
wire [0:0] ram_block3a10_PORTBDATAOUT_bus;
wire [0:0] ram_block3a43_PORTADATAOUT_bus;
wire [0:0] ram_block3a43_PORTBDATAOUT_bus;
wire [0:0] ram_block3a11_PORTADATAOUT_bus;
wire [0:0] ram_block3a11_PORTBDATAOUT_bus;
wire [0:0] ram_block3a44_PORTADATAOUT_bus;
wire [0:0] ram_block3a44_PORTBDATAOUT_bus;
wire [0:0] ram_block3a12_PORTADATAOUT_bus;
wire [0:0] ram_block3a12_PORTBDATAOUT_bus;
wire [0:0] ram_block3a45_PORTADATAOUT_bus;
wire [0:0] ram_block3a45_PORTBDATAOUT_bus;
wire [0:0] ram_block3a13_PORTADATAOUT_bus;
wire [0:0] ram_block3a13_PORTBDATAOUT_bus;
wire [0:0] ram_block3a46_PORTADATAOUT_bus;
wire [0:0] ram_block3a46_PORTBDATAOUT_bus;
wire [0:0] ram_block3a14_PORTADATAOUT_bus;
wire [0:0] ram_block3a14_PORTBDATAOUT_bus;
wire [0:0] ram_block3a47_PORTADATAOUT_bus;
wire [0:0] ram_block3a47_PORTBDATAOUT_bus;
wire [0:0] ram_block3a15_PORTADATAOUT_bus;
wire [0:0] ram_block3a15_PORTBDATAOUT_bus;
wire [0:0] ram_block3a48_PORTADATAOUT_bus;
wire [0:0] ram_block3a48_PORTBDATAOUT_bus;
wire [0:0] ram_block3a16_PORTADATAOUT_bus;
wire [0:0] ram_block3a16_PORTBDATAOUT_bus;
wire [0:0] ram_block3a49_PORTADATAOUT_bus;
wire [0:0] ram_block3a49_PORTBDATAOUT_bus;
wire [0:0] ram_block3a17_PORTADATAOUT_bus;
wire [0:0] ram_block3a17_PORTBDATAOUT_bus;
wire [0:0] ram_block3a50_PORTADATAOUT_bus;
wire [0:0] ram_block3a50_PORTBDATAOUT_bus;
wire [0:0] ram_block3a18_PORTADATAOUT_bus;
wire [0:0] ram_block3a18_PORTBDATAOUT_bus;
wire [0:0] ram_block3a51_PORTADATAOUT_bus;
wire [0:0] ram_block3a51_PORTBDATAOUT_bus;
wire [0:0] ram_block3a19_PORTADATAOUT_bus;
wire [0:0] ram_block3a19_PORTBDATAOUT_bus;
wire [0:0] ram_block3a52_PORTADATAOUT_bus;
wire [0:0] ram_block3a52_PORTBDATAOUT_bus;
wire [0:0] ram_block3a20_PORTADATAOUT_bus;
wire [0:0] ram_block3a20_PORTBDATAOUT_bus;
wire [0:0] ram_block3a53_PORTADATAOUT_bus;
wire [0:0] ram_block3a53_PORTBDATAOUT_bus;
wire [0:0] ram_block3a21_PORTADATAOUT_bus;
wire [0:0] ram_block3a21_PORTBDATAOUT_bus;
wire [0:0] ram_block3a54_PORTADATAOUT_bus;
wire [0:0] ram_block3a54_PORTBDATAOUT_bus;
wire [0:0] ram_block3a22_PORTADATAOUT_bus;
wire [0:0] ram_block3a22_PORTBDATAOUT_bus;
wire [0:0] ram_block3a55_PORTADATAOUT_bus;
wire [0:0] ram_block3a55_PORTBDATAOUT_bus;
wire [0:0] ram_block3a23_PORTADATAOUT_bus;
wire [0:0] ram_block3a23_PORTBDATAOUT_bus;
wire [0:0] ram_block3a56_PORTADATAOUT_bus;
wire [0:0] ram_block3a56_PORTBDATAOUT_bus;
wire [0:0] ram_block3a24_PORTADATAOUT_bus;
wire [0:0] ram_block3a24_PORTBDATAOUT_bus;
wire [0:0] ram_block3a57_PORTADATAOUT_bus;
wire [0:0] ram_block3a57_PORTBDATAOUT_bus;
wire [0:0] ram_block3a25_PORTADATAOUT_bus;
wire [0:0] ram_block3a25_PORTBDATAOUT_bus;
wire [0:0] ram_block3a58_PORTADATAOUT_bus;
wire [0:0] ram_block3a58_PORTBDATAOUT_bus;
wire [0:0] ram_block3a26_PORTADATAOUT_bus;
wire [0:0] ram_block3a26_PORTBDATAOUT_bus;
wire [0:0] ram_block3a59_PORTADATAOUT_bus;
wire [0:0] ram_block3a59_PORTBDATAOUT_bus;
wire [0:0] ram_block3a27_PORTADATAOUT_bus;
wire [0:0] ram_block3a27_PORTBDATAOUT_bus;
wire [0:0] ram_block3a60_PORTADATAOUT_bus;
wire [0:0] ram_block3a60_PORTBDATAOUT_bus;
wire [0:0] ram_block3a28_PORTADATAOUT_bus;
wire [0:0] ram_block3a28_PORTBDATAOUT_bus;
wire [0:0] ram_block3a61_PORTADATAOUT_bus;
wire [0:0] ram_block3a61_PORTBDATAOUT_bus;
wire [0:0] ram_block3a29_PORTADATAOUT_bus;
wire [0:0] ram_block3a29_PORTBDATAOUT_bus;
wire [0:0] ram_block3a62_PORTADATAOUT_bus;
wire [0:0] ram_block3a62_PORTBDATAOUT_bus;
wire [0:0] ram_block3a30_PORTADATAOUT_bus;
wire [0:0] ram_block3a30_PORTBDATAOUT_bus;
wire [0:0] ram_block3a63_PORTADATAOUT_bus;
wire [0:0] ram_block3a63_PORTBDATAOUT_bus;
wire [0:0] ram_block3a31_PORTADATAOUT_bus;
wire [0:0] ram_block3a31_PORTBDATAOUT_bus;

assign ram_block3a321 = ram_block3a32_PORTADATAOUT_bus[0];

assign ram_block3a322 = ram_block3a32_PORTBDATAOUT_bus[0];

assign ram_block3a01 = ram_block3a0_PORTADATAOUT_bus[0];

assign ram_block3a02 = ram_block3a0_PORTBDATAOUT_bus[0];

assign ram_block3a331 = ram_block3a33_PORTADATAOUT_bus[0];

assign ram_block3a332 = ram_block3a33_PORTBDATAOUT_bus[0];

assign ram_block3a110 = ram_block3a1_PORTADATAOUT_bus[0];

assign ram_block3a111 = ram_block3a1_PORTBDATAOUT_bus[0];

assign ram_block3a341 = ram_block3a34_PORTADATAOUT_bus[0];

assign ram_block3a342 = ram_block3a34_PORTBDATAOUT_bus[0];

assign ram_block3a210 = ram_block3a2_PORTADATAOUT_bus[0];

assign ram_block3a211 = ram_block3a2_PORTBDATAOUT_bus[0];

assign ram_block3a351 = ram_block3a35_PORTADATAOUT_bus[0];

assign ram_block3a352 = ram_block3a35_PORTBDATAOUT_bus[0];

assign ram_block3a310 = ram_block3a3_PORTADATAOUT_bus[0];

assign ram_block3a311 = ram_block3a3_PORTBDATAOUT_bus[0];

assign ram_block3a361 = ram_block3a36_PORTADATAOUT_bus[0];

assign ram_block3a362 = ram_block3a36_PORTBDATAOUT_bus[0];

assign ram_block3a410 = ram_block3a4_PORTADATAOUT_bus[0];

assign ram_block3a411 = ram_block3a4_PORTBDATAOUT_bus[0];

assign ram_block3a371 = ram_block3a37_PORTADATAOUT_bus[0];

assign ram_block3a372 = ram_block3a37_PORTBDATAOUT_bus[0];

assign ram_block3a510 = ram_block3a5_PORTADATAOUT_bus[0];

assign ram_block3a511 = ram_block3a5_PORTBDATAOUT_bus[0];

assign ram_block3a381 = ram_block3a38_PORTADATAOUT_bus[0];

assign ram_block3a382 = ram_block3a38_PORTBDATAOUT_bus[0];

assign ram_block3a64 = ram_block3a6_PORTADATAOUT_bus[0];

assign ram_block3a65 = ram_block3a6_PORTBDATAOUT_bus[0];

assign ram_block3a391 = ram_block3a39_PORTADATAOUT_bus[0];

assign ram_block3a392 = ram_block3a39_PORTBDATAOUT_bus[0];

assign ram_block3a71 = ram_block3a7_PORTADATAOUT_bus[0];

assign ram_block3a72 = ram_block3a7_PORTBDATAOUT_bus[0];

assign ram_block3a401 = ram_block3a40_PORTADATAOUT_bus[0];

assign ram_block3a402 = ram_block3a40_PORTBDATAOUT_bus[0];

assign ram_block3a81 = ram_block3a8_PORTADATAOUT_bus[0];

assign ram_block3a82 = ram_block3a8_PORTBDATAOUT_bus[0];

assign ram_block3a412 = ram_block3a41_PORTADATAOUT_bus[0];

assign ram_block3a413 = ram_block3a41_PORTBDATAOUT_bus[0];

assign ram_block3a91 = ram_block3a9_PORTADATAOUT_bus[0];

assign ram_block3a92 = ram_block3a9_PORTBDATAOUT_bus[0];

assign ram_block3a421 = ram_block3a42_PORTADATAOUT_bus[0];

assign ram_block3a422 = ram_block3a42_PORTBDATAOUT_bus[0];

assign ram_block3a101 = ram_block3a10_PORTADATAOUT_bus[0];

assign ram_block3a102 = ram_block3a10_PORTBDATAOUT_bus[0];

assign ram_block3a431 = ram_block3a43_PORTADATAOUT_bus[0];

assign ram_block3a432 = ram_block3a43_PORTBDATAOUT_bus[0];

assign ram_block3a112 = ram_block3a11_PORTADATAOUT_bus[0];

assign ram_block3a113 = ram_block3a11_PORTBDATAOUT_bus[0];

assign ram_block3a441 = ram_block3a44_PORTADATAOUT_bus[0];

assign ram_block3a442 = ram_block3a44_PORTBDATAOUT_bus[0];

assign ram_block3a121 = ram_block3a12_PORTADATAOUT_bus[0];

assign ram_block3a122 = ram_block3a12_PORTBDATAOUT_bus[0];

assign ram_block3a451 = ram_block3a45_PORTADATAOUT_bus[0];

assign ram_block3a452 = ram_block3a45_PORTBDATAOUT_bus[0];

assign ram_block3a131 = ram_block3a13_PORTADATAOUT_bus[0];

assign ram_block3a132 = ram_block3a13_PORTBDATAOUT_bus[0];

assign ram_block3a461 = ram_block3a46_PORTADATAOUT_bus[0];

assign ram_block3a462 = ram_block3a46_PORTBDATAOUT_bus[0];

assign ram_block3a141 = ram_block3a14_PORTADATAOUT_bus[0];

assign ram_block3a142 = ram_block3a14_PORTBDATAOUT_bus[0];

assign ram_block3a471 = ram_block3a47_PORTADATAOUT_bus[0];

assign ram_block3a472 = ram_block3a47_PORTBDATAOUT_bus[0];

assign ram_block3a151 = ram_block3a15_PORTADATAOUT_bus[0];

assign ram_block3a152 = ram_block3a15_PORTBDATAOUT_bus[0];

assign ram_block3a481 = ram_block3a48_PORTADATAOUT_bus[0];

assign ram_block3a482 = ram_block3a48_PORTBDATAOUT_bus[0];

assign ram_block3a161 = ram_block3a16_PORTADATAOUT_bus[0];

assign ram_block3a162 = ram_block3a16_PORTBDATAOUT_bus[0];

assign ram_block3a491 = ram_block3a49_PORTADATAOUT_bus[0];

assign ram_block3a492 = ram_block3a49_PORTBDATAOUT_bus[0];

assign ram_block3a171 = ram_block3a17_PORTADATAOUT_bus[0];

assign ram_block3a172 = ram_block3a17_PORTBDATAOUT_bus[0];

assign ram_block3a501 = ram_block3a50_PORTADATAOUT_bus[0];

assign ram_block3a502 = ram_block3a50_PORTBDATAOUT_bus[0];

assign ram_block3a181 = ram_block3a18_PORTADATAOUT_bus[0];

assign ram_block3a182 = ram_block3a18_PORTBDATAOUT_bus[0];

assign ram_block3a512 = ram_block3a51_PORTADATAOUT_bus[0];

assign ram_block3a513 = ram_block3a51_PORTBDATAOUT_bus[0];

assign ram_block3a191 = ram_block3a19_PORTADATAOUT_bus[0];

assign ram_block3a192 = ram_block3a19_PORTBDATAOUT_bus[0];

assign ram_block3a521 = ram_block3a52_PORTADATAOUT_bus[0];

assign ram_block3a522 = ram_block3a52_PORTBDATAOUT_bus[0];

assign ram_block3a201 = ram_block3a20_PORTADATAOUT_bus[0];

assign ram_block3a202 = ram_block3a20_PORTBDATAOUT_bus[0];

assign ram_block3a531 = ram_block3a53_PORTADATAOUT_bus[0];

assign ram_block3a532 = ram_block3a53_PORTBDATAOUT_bus[0];

assign ram_block3a212 = ram_block3a21_PORTADATAOUT_bus[0];

assign ram_block3a213 = ram_block3a21_PORTBDATAOUT_bus[0];

assign ram_block3a541 = ram_block3a54_PORTADATAOUT_bus[0];

assign ram_block3a542 = ram_block3a54_PORTBDATAOUT_bus[0];

assign ram_block3a221 = ram_block3a22_PORTADATAOUT_bus[0];

assign ram_block3a222 = ram_block3a22_PORTBDATAOUT_bus[0];

assign ram_block3a551 = ram_block3a55_PORTADATAOUT_bus[0];

assign ram_block3a552 = ram_block3a55_PORTBDATAOUT_bus[0];

assign ram_block3a231 = ram_block3a23_PORTADATAOUT_bus[0];

assign ram_block3a232 = ram_block3a23_PORTBDATAOUT_bus[0];

assign ram_block3a561 = ram_block3a56_PORTADATAOUT_bus[0];

assign ram_block3a562 = ram_block3a56_PORTBDATAOUT_bus[0];

assign ram_block3a241 = ram_block3a24_PORTADATAOUT_bus[0];

assign ram_block3a242 = ram_block3a24_PORTBDATAOUT_bus[0];

assign ram_block3a571 = ram_block3a57_PORTADATAOUT_bus[0];

assign ram_block3a572 = ram_block3a57_PORTBDATAOUT_bus[0];

assign ram_block3a251 = ram_block3a25_PORTADATAOUT_bus[0];

assign ram_block3a252 = ram_block3a25_PORTBDATAOUT_bus[0];

assign ram_block3a581 = ram_block3a58_PORTADATAOUT_bus[0];

assign ram_block3a582 = ram_block3a58_PORTBDATAOUT_bus[0];

assign ram_block3a261 = ram_block3a26_PORTADATAOUT_bus[0];

assign ram_block3a262 = ram_block3a26_PORTBDATAOUT_bus[0];

assign ram_block3a591 = ram_block3a59_PORTADATAOUT_bus[0];

assign ram_block3a592 = ram_block3a59_PORTBDATAOUT_bus[0];

assign ram_block3a271 = ram_block3a27_PORTADATAOUT_bus[0];

assign ram_block3a272 = ram_block3a27_PORTBDATAOUT_bus[0];

assign ram_block3a601 = ram_block3a60_PORTADATAOUT_bus[0];

assign ram_block3a602 = ram_block3a60_PORTBDATAOUT_bus[0];

assign ram_block3a281 = ram_block3a28_PORTADATAOUT_bus[0];

assign ram_block3a282 = ram_block3a28_PORTBDATAOUT_bus[0];

assign ram_block3a611 = ram_block3a61_PORTADATAOUT_bus[0];

assign ram_block3a612 = ram_block3a61_PORTBDATAOUT_bus[0];

assign ram_block3a291 = ram_block3a29_PORTADATAOUT_bus[0];

assign ram_block3a292 = ram_block3a29_PORTBDATAOUT_bus[0];

assign ram_block3a621 = ram_block3a62_PORTADATAOUT_bus[0];

assign ram_block3a622 = ram_block3a62_PORTBDATAOUT_bus[0];

assign ram_block3a301 = ram_block3a30_PORTADATAOUT_bus[0];

assign ram_block3a302 = ram_block3a30_PORTBDATAOUT_bus[0];

assign ram_block3a631 = ram_block3a63_PORTADATAOUT_bus[0];

assign ram_block3a632 = ram_block3a63_PORTBDATAOUT_bus[0];

assign ram_block3a312 = ram_block3a31_PORTADATAOUT_bus[0];

assign ram_block3a313 = ram_block3a31_PORTBDATAOUT_bus[0];

decode_jsa_1 decode5(
	.ram_rom_addr_reg_13(ram_rom_addr_reg_13),
	.sdr(sdr),
	.eq_node_1(\decode5|eq_node[1]~0_combout ),
	.eq_node_0(\decode5|eq_node[0]~1_combout ),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

decode_jsa decode4(
	.ramaddr(ramaddr),
	.always1(always1),
	.ramWEN(ramWEN),
	.eq_node_1(\decode4|eq_node[1]~0_combout ),
	.eq_node_0(\decode4|eq_node[0]~1_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: M9K_X51_Y35_N0
cycloneive_ram_block ram_block3a32(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a32_PORTADATAOUT_bus),
	.portbdataout(ram_block3a32_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a32.clk0_core_clock_enable = "ena0";
defparam ram_block3a32.clk1_core_clock_enable = "ena1";
defparam ram_block3a32.data_interleave_offset_in_bits = 1;
defparam ram_block3a32.data_interleave_width_in_bits = 1;
defparam ram_block3a32.init_file = "meminit.hex";
defparam ram_block3a32.init_file_layout = "port_a";
defparam ram_block3a32.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a32.operation_mode = "bidir_dual_port";
defparam ram_block3a32.port_a_address_clear = "none";
defparam ram_block3a32.port_a_address_width = 13;
defparam ram_block3a32.port_a_byte_enable_clock = "none";
defparam ram_block3a32.port_a_data_out_clear = "none";
defparam ram_block3a32.port_a_data_out_clock = "none";
defparam ram_block3a32.port_a_data_width = 1;
defparam ram_block3a32.port_a_first_address = 0;
defparam ram_block3a32.port_a_first_bit_number = 0;
defparam ram_block3a32.port_a_last_address = 8191;
defparam ram_block3a32.port_a_logical_ram_depth = 16384;
defparam ram_block3a32.port_a_logical_ram_width = 32;
defparam ram_block3a32.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_address_clear = "none";
defparam ram_block3a32.port_b_address_clock = "clock1";
defparam ram_block3a32.port_b_address_width = 13;
defparam ram_block3a32.port_b_data_in_clock = "clock1";
defparam ram_block3a32.port_b_data_out_clear = "none";
defparam ram_block3a32.port_b_data_out_clock = "none";
defparam ram_block3a32.port_b_data_width = 1;
defparam ram_block3a32.port_b_first_address = 0;
defparam ram_block3a32.port_b_first_bit_number = 0;
defparam ram_block3a32.port_b_last_address = 8191;
defparam ram_block3a32.port_b_logical_ram_depth = 16384;
defparam ram_block3a32.port_b_logical_ram_width = 32;
defparam ram_block3a32.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_read_enable_clock = "clock1";
defparam ram_block3a32.port_b_write_enable_clock = "clock1";
defparam ram_block3a32.ram_block_type = "M9K";
defparam ram_block3a32.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y35_N0
cycloneive_ram_block ram_block3a0(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a0_PORTADATAOUT_bus),
	.portbdataout(ram_block3a0_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a0.clk0_core_clock_enable = "ena0";
defparam ram_block3a0.clk1_core_clock_enable = "ena1";
defparam ram_block3a0.data_interleave_offset_in_bits = 1;
defparam ram_block3a0.data_interleave_width_in_bits = 1;
defparam ram_block3a0.init_file = "meminit.hex";
defparam ram_block3a0.init_file_layout = "port_a";
defparam ram_block3a0.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a0.operation_mode = "bidir_dual_port";
defparam ram_block3a0.port_a_address_clear = "none";
defparam ram_block3a0.port_a_address_width = 13;
defparam ram_block3a0.port_a_byte_enable_clock = "none";
defparam ram_block3a0.port_a_data_out_clear = "none";
defparam ram_block3a0.port_a_data_out_clock = "none";
defparam ram_block3a0.port_a_data_width = 1;
defparam ram_block3a0.port_a_first_address = 0;
defparam ram_block3a0.port_a_first_bit_number = 0;
defparam ram_block3a0.port_a_last_address = 8191;
defparam ram_block3a0.port_a_logical_ram_depth = 16384;
defparam ram_block3a0.port_a_logical_ram_width = 32;
defparam ram_block3a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_address_clear = "none";
defparam ram_block3a0.port_b_address_clock = "clock1";
defparam ram_block3a0.port_b_address_width = 13;
defparam ram_block3a0.port_b_data_in_clock = "clock1";
defparam ram_block3a0.port_b_data_out_clear = "none";
defparam ram_block3a0.port_b_data_out_clock = "none";
defparam ram_block3a0.port_b_data_width = 1;
defparam ram_block3a0.port_b_first_address = 0;
defparam ram_block3a0.port_b_first_bit_number = 0;
defparam ram_block3a0.port_b_last_address = 8191;
defparam ram_block3a0.port_b_logical_ram_depth = 16384;
defparam ram_block3a0.port_b_logical_ram_width = 32;
defparam ram_block3a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_read_enable_clock = "clock1";
defparam ram_block3a0.port_b_write_enable_clock = "clock1";
defparam ram_block3a0.ram_block_type = "M9K";
defparam ram_block3a0.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004004AD3;
// synopsys translate_on

// Location: M9K_X51_Y37_N0
cycloneive_ram_block ram_block3a33(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a33_PORTADATAOUT_bus),
	.portbdataout(ram_block3a33_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a33.clk0_core_clock_enable = "ena0";
defparam ram_block3a33.clk1_core_clock_enable = "ena1";
defparam ram_block3a33.data_interleave_offset_in_bits = 1;
defparam ram_block3a33.data_interleave_width_in_bits = 1;
defparam ram_block3a33.init_file = "meminit.hex";
defparam ram_block3a33.init_file_layout = "port_a";
defparam ram_block3a33.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a33.operation_mode = "bidir_dual_port";
defparam ram_block3a33.port_a_address_clear = "none";
defparam ram_block3a33.port_a_address_width = 13;
defparam ram_block3a33.port_a_byte_enable_clock = "none";
defparam ram_block3a33.port_a_data_out_clear = "none";
defparam ram_block3a33.port_a_data_out_clock = "none";
defparam ram_block3a33.port_a_data_width = 1;
defparam ram_block3a33.port_a_first_address = 0;
defparam ram_block3a33.port_a_first_bit_number = 1;
defparam ram_block3a33.port_a_last_address = 8191;
defparam ram_block3a33.port_a_logical_ram_depth = 16384;
defparam ram_block3a33.port_a_logical_ram_width = 32;
defparam ram_block3a33.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_address_clear = "none";
defparam ram_block3a33.port_b_address_clock = "clock1";
defparam ram_block3a33.port_b_address_width = 13;
defparam ram_block3a33.port_b_data_in_clock = "clock1";
defparam ram_block3a33.port_b_data_out_clear = "none";
defparam ram_block3a33.port_b_data_out_clock = "none";
defparam ram_block3a33.port_b_data_width = 1;
defparam ram_block3a33.port_b_first_address = 0;
defparam ram_block3a33.port_b_first_bit_number = 1;
defparam ram_block3a33.port_b_last_address = 8191;
defparam ram_block3a33.port_b_logical_ram_depth = 16384;
defparam ram_block3a33.port_b_logical_ram_width = 32;
defparam ram_block3a33.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_read_enable_clock = "clock1";
defparam ram_block3a33.port_b_write_enable_clock = "clock1";
defparam ram_block3a33.ram_block_type = "M9K";
defparam ram_block3a33.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y34_N0
cycloneive_ram_block ram_block3a1(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a1_PORTADATAOUT_bus),
	.portbdataout(ram_block3a1_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a1.clk0_core_clock_enable = "ena0";
defparam ram_block3a1.clk1_core_clock_enable = "ena1";
defparam ram_block3a1.data_interleave_offset_in_bits = 1;
defparam ram_block3a1.data_interleave_width_in_bits = 1;
defparam ram_block3a1.init_file = "meminit.hex";
defparam ram_block3a1.init_file_layout = "port_a";
defparam ram_block3a1.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a1.operation_mode = "bidir_dual_port";
defparam ram_block3a1.port_a_address_clear = "none";
defparam ram_block3a1.port_a_address_width = 13;
defparam ram_block3a1.port_a_byte_enable_clock = "none";
defparam ram_block3a1.port_a_data_out_clear = "none";
defparam ram_block3a1.port_a_data_out_clock = "none";
defparam ram_block3a1.port_a_data_width = 1;
defparam ram_block3a1.port_a_first_address = 0;
defparam ram_block3a1.port_a_first_bit_number = 1;
defparam ram_block3a1.port_a_last_address = 8191;
defparam ram_block3a1.port_a_logical_ram_depth = 16384;
defparam ram_block3a1.port_a_logical_ram_width = 32;
defparam ram_block3a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_address_clear = "none";
defparam ram_block3a1.port_b_address_clock = "clock1";
defparam ram_block3a1.port_b_address_width = 13;
defparam ram_block3a1.port_b_data_in_clock = "clock1";
defparam ram_block3a1.port_b_data_out_clear = "none";
defparam ram_block3a1.port_b_data_out_clock = "none";
defparam ram_block3a1.port_b_data_width = 1;
defparam ram_block3a1.port_b_first_address = 0;
defparam ram_block3a1.port_b_first_bit_number = 1;
defparam ram_block3a1.port_b_last_address = 8191;
defparam ram_block3a1.port_b_logical_ram_depth = 16384;
defparam ram_block3a1.port_b_logical_ram_width = 32;
defparam ram_block3a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_read_enable_clock = "clock1";
defparam ram_block3a1.port_b_write_enable_clock = "clock1";
defparam ram_block3a1.ram_block_type = "M9K";
defparam ram_block3a1.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004006E40;
// synopsys translate_on

// Location: M9K_X51_Y33_N0
cycloneive_ram_block ram_block3a34(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a34_PORTADATAOUT_bus),
	.portbdataout(ram_block3a34_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a34.clk0_core_clock_enable = "ena0";
defparam ram_block3a34.clk1_core_clock_enable = "ena1";
defparam ram_block3a34.data_interleave_offset_in_bits = 1;
defparam ram_block3a34.data_interleave_width_in_bits = 1;
defparam ram_block3a34.init_file = "meminit.hex";
defparam ram_block3a34.init_file_layout = "port_a";
defparam ram_block3a34.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a34.operation_mode = "bidir_dual_port";
defparam ram_block3a34.port_a_address_clear = "none";
defparam ram_block3a34.port_a_address_width = 13;
defparam ram_block3a34.port_a_byte_enable_clock = "none";
defparam ram_block3a34.port_a_data_out_clear = "none";
defparam ram_block3a34.port_a_data_out_clock = "none";
defparam ram_block3a34.port_a_data_width = 1;
defparam ram_block3a34.port_a_first_address = 0;
defparam ram_block3a34.port_a_first_bit_number = 2;
defparam ram_block3a34.port_a_last_address = 8191;
defparam ram_block3a34.port_a_logical_ram_depth = 16384;
defparam ram_block3a34.port_a_logical_ram_width = 32;
defparam ram_block3a34.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_address_clear = "none";
defparam ram_block3a34.port_b_address_clock = "clock1";
defparam ram_block3a34.port_b_address_width = 13;
defparam ram_block3a34.port_b_data_in_clock = "clock1";
defparam ram_block3a34.port_b_data_out_clear = "none";
defparam ram_block3a34.port_b_data_out_clock = "none";
defparam ram_block3a34.port_b_data_width = 1;
defparam ram_block3a34.port_b_first_address = 0;
defparam ram_block3a34.port_b_first_bit_number = 2;
defparam ram_block3a34.port_b_last_address = 8191;
defparam ram_block3a34.port_b_logical_ram_depth = 16384;
defparam ram_block3a34.port_b_logical_ram_width = 32;
defparam ram_block3a34.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_read_enable_clock = "clock1";
defparam ram_block3a34.port_b_write_enable_clock = "clock1";
defparam ram_block3a34.ram_block_type = "M9K";
defparam ram_block3a34.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y31_N0
cycloneive_ram_block ram_block3a2(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a2_PORTADATAOUT_bus),
	.portbdataout(ram_block3a2_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a2.clk0_core_clock_enable = "ena0";
defparam ram_block3a2.clk1_core_clock_enable = "ena1";
defparam ram_block3a2.data_interleave_offset_in_bits = 1;
defparam ram_block3a2.data_interleave_width_in_bits = 1;
defparam ram_block3a2.init_file = "meminit.hex";
defparam ram_block3a2.init_file_layout = "port_a";
defparam ram_block3a2.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a2.operation_mode = "bidir_dual_port";
defparam ram_block3a2.port_a_address_clear = "none";
defparam ram_block3a2.port_a_address_width = 13;
defparam ram_block3a2.port_a_byte_enable_clock = "none";
defparam ram_block3a2.port_a_data_out_clear = "none";
defparam ram_block3a2.port_a_data_out_clock = "none";
defparam ram_block3a2.port_a_data_width = 1;
defparam ram_block3a2.port_a_first_address = 0;
defparam ram_block3a2.port_a_first_bit_number = 2;
defparam ram_block3a2.port_a_last_address = 8191;
defparam ram_block3a2.port_a_logical_ram_depth = 16384;
defparam ram_block3a2.port_a_logical_ram_width = 32;
defparam ram_block3a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_address_clear = "none";
defparam ram_block3a2.port_b_address_clock = "clock1";
defparam ram_block3a2.port_b_address_width = 13;
defparam ram_block3a2.port_b_data_in_clock = "clock1";
defparam ram_block3a2.port_b_data_out_clear = "none";
defparam ram_block3a2.port_b_data_out_clock = "none";
defparam ram_block3a2.port_b_data_width = 1;
defparam ram_block3a2.port_b_first_address = 0;
defparam ram_block3a2.port_b_first_bit_number = 2;
defparam ram_block3a2.port_b_last_address = 8191;
defparam ram_block3a2.port_b_logical_ram_depth = 16384;
defparam ram_block3a2.port_b_logical_ram_width = 32;
defparam ram_block3a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_read_enable_clock = "clock1";
defparam ram_block3a2.port_b_write_enable_clock = "clock1";
defparam ram_block3a2.ram_block_type = "M9K";
defparam ram_block3a2.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006AA4C70;
// synopsys translate_on

// Location: M9K_X64_Y33_N0
cycloneive_ram_block ram_block3a35(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a35_PORTADATAOUT_bus),
	.portbdataout(ram_block3a35_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a35.clk0_core_clock_enable = "ena0";
defparam ram_block3a35.clk1_core_clock_enable = "ena1";
defparam ram_block3a35.data_interleave_offset_in_bits = 1;
defparam ram_block3a35.data_interleave_width_in_bits = 1;
defparam ram_block3a35.init_file = "meminit.hex";
defparam ram_block3a35.init_file_layout = "port_a";
defparam ram_block3a35.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a35.operation_mode = "bidir_dual_port";
defparam ram_block3a35.port_a_address_clear = "none";
defparam ram_block3a35.port_a_address_width = 13;
defparam ram_block3a35.port_a_byte_enable_clock = "none";
defparam ram_block3a35.port_a_data_out_clear = "none";
defparam ram_block3a35.port_a_data_out_clock = "none";
defparam ram_block3a35.port_a_data_width = 1;
defparam ram_block3a35.port_a_first_address = 0;
defparam ram_block3a35.port_a_first_bit_number = 3;
defparam ram_block3a35.port_a_last_address = 8191;
defparam ram_block3a35.port_a_logical_ram_depth = 16384;
defparam ram_block3a35.port_a_logical_ram_width = 32;
defparam ram_block3a35.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_address_clear = "none";
defparam ram_block3a35.port_b_address_clock = "clock1";
defparam ram_block3a35.port_b_address_width = 13;
defparam ram_block3a35.port_b_data_in_clock = "clock1";
defparam ram_block3a35.port_b_data_out_clear = "none";
defparam ram_block3a35.port_b_data_out_clock = "none";
defparam ram_block3a35.port_b_data_width = 1;
defparam ram_block3a35.port_b_first_address = 0;
defparam ram_block3a35.port_b_first_bit_number = 3;
defparam ram_block3a35.port_b_last_address = 8191;
defparam ram_block3a35.port_b_logical_ram_depth = 16384;
defparam ram_block3a35.port_b_logical_ram_width = 32;
defparam ram_block3a35.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_read_enable_clock = "clock1";
defparam ram_block3a35.port_b_write_enable_clock = "clock1";
defparam ram_block3a35.ram_block_type = "M9K";
defparam ram_block3a35.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y33_N0
cycloneive_ram_block ram_block3a3(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a3_PORTADATAOUT_bus),
	.portbdataout(ram_block3a3_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a3.clk0_core_clock_enable = "ena0";
defparam ram_block3a3.clk1_core_clock_enable = "ena1";
defparam ram_block3a3.data_interleave_offset_in_bits = 1;
defparam ram_block3a3.data_interleave_width_in_bits = 1;
defparam ram_block3a3.init_file = "meminit.hex";
defparam ram_block3a3.init_file_layout = "port_a";
defparam ram_block3a3.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a3.operation_mode = "bidir_dual_port";
defparam ram_block3a3.port_a_address_clear = "none";
defparam ram_block3a3.port_a_address_width = 13;
defparam ram_block3a3.port_a_byte_enable_clock = "none";
defparam ram_block3a3.port_a_data_out_clear = "none";
defparam ram_block3a3.port_a_data_out_clock = "none";
defparam ram_block3a3.port_a_data_width = 1;
defparam ram_block3a3.port_a_first_address = 0;
defparam ram_block3a3.port_a_first_bit_number = 3;
defparam ram_block3a3.port_a_last_address = 8191;
defparam ram_block3a3.port_a_logical_ram_depth = 16384;
defparam ram_block3a3.port_a_logical_ram_width = 32;
defparam ram_block3a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_address_clear = "none";
defparam ram_block3a3.port_b_address_clock = "clock1";
defparam ram_block3a3.port_b_address_width = 13;
defparam ram_block3a3.port_b_data_in_clock = "clock1";
defparam ram_block3a3.port_b_data_out_clear = "none";
defparam ram_block3a3.port_b_data_out_clock = "none";
defparam ram_block3a3.port_b_data_width = 1;
defparam ram_block3a3.port_b_first_address = 0;
defparam ram_block3a3.port_b_first_bit_number = 3;
defparam ram_block3a3.port_b_last_address = 8191;
defparam ram_block3a3.port_b_logical_ram_depth = 16384;
defparam ram_block3a3.port_b_logical_ram_width = 32;
defparam ram_block3a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_read_enable_clock = "clock1";
defparam ram_block3a3.port_b_write_enable_clock = "clock1";
defparam ram_block3a3.ram_block_type = "M9K";
defparam ram_block3a3.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004CC0841;
// synopsys translate_on

// Location: M9K_X37_Y29_N0
cycloneive_ram_block ram_block3a36(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a36_PORTADATAOUT_bus),
	.portbdataout(ram_block3a36_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a36.clk0_core_clock_enable = "ena0";
defparam ram_block3a36.clk1_core_clock_enable = "ena1";
defparam ram_block3a36.data_interleave_offset_in_bits = 1;
defparam ram_block3a36.data_interleave_width_in_bits = 1;
defparam ram_block3a36.init_file = "meminit.hex";
defparam ram_block3a36.init_file_layout = "port_a";
defparam ram_block3a36.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a36.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a36.operation_mode = "bidir_dual_port";
defparam ram_block3a36.port_a_address_clear = "none";
defparam ram_block3a36.port_a_address_width = 13;
defparam ram_block3a36.port_a_byte_enable_clock = "none";
defparam ram_block3a36.port_a_data_out_clear = "none";
defparam ram_block3a36.port_a_data_out_clock = "none";
defparam ram_block3a36.port_a_data_width = 1;
defparam ram_block3a36.port_a_first_address = 0;
defparam ram_block3a36.port_a_first_bit_number = 4;
defparam ram_block3a36.port_a_last_address = 8191;
defparam ram_block3a36.port_a_logical_ram_depth = 16384;
defparam ram_block3a36.port_a_logical_ram_width = 32;
defparam ram_block3a36.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_address_clear = "none";
defparam ram_block3a36.port_b_address_clock = "clock1";
defparam ram_block3a36.port_b_address_width = 13;
defparam ram_block3a36.port_b_data_in_clock = "clock1";
defparam ram_block3a36.port_b_data_out_clear = "none";
defparam ram_block3a36.port_b_data_out_clock = "none";
defparam ram_block3a36.port_b_data_width = 1;
defparam ram_block3a36.port_b_first_address = 0;
defparam ram_block3a36.port_b_first_bit_number = 4;
defparam ram_block3a36.port_b_last_address = 8191;
defparam ram_block3a36.port_b_logical_ram_depth = 16384;
defparam ram_block3a36.port_b_logical_ram_width = 32;
defparam ram_block3a36.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_read_enable_clock = "clock1";
defparam ram_block3a36.port_b_write_enable_clock = "clock1";
defparam ram_block3a36.ram_block_type = "M9K";
defparam ram_block3a36.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y30_N0
cycloneive_ram_block ram_block3a4(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a4_PORTADATAOUT_bus),
	.portbdataout(ram_block3a4_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a4.clk0_core_clock_enable = "ena0";
defparam ram_block3a4.clk1_core_clock_enable = "ena1";
defparam ram_block3a4.data_interleave_offset_in_bits = 1;
defparam ram_block3a4.data_interleave_width_in_bits = 1;
defparam ram_block3a4.init_file = "meminit.hex";
defparam ram_block3a4.init_file_layout = "port_a";
defparam ram_block3a4.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a4.operation_mode = "bidir_dual_port";
defparam ram_block3a4.port_a_address_clear = "none";
defparam ram_block3a4.port_a_address_width = 13;
defparam ram_block3a4.port_a_byte_enable_clock = "none";
defparam ram_block3a4.port_a_data_out_clear = "none";
defparam ram_block3a4.port_a_data_out_clock = "none";
defparam ram_block3a4.port_a_data_width = 1;
defparam ram_block3a4.port_a_first_address = 0;
defparam ram_block3a4.port_a_first_bit_number = 4;
defparam ram_block3a4.port_a_last_address = 8191;
defparam ram_block3a4.port_a_logical_ram_depth = 16384;
defparam ram_block3a4.port_a_logical_ram_width = 32;
defparam ram_block3a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_address_clear = "none";
defparam ram_block3a4.port_b_address_clock = "clock1";
defparam ram_block3a4.port_b_address_width = 13;
defparam ram_block3a4.port_b_data_in_clock = "clock1";
defparam ram_block3a4.port_b_data_out_clear = "none";
defparam ram_block3a4.port_b_data_out_clock = "none";
defparam ram_block3a4.port_b_data_width = 1;
defparam ram_block3a4.port_b_first_address = 0;
defparam ram_block3a4.port_b_first_bit_number = 4;
defparam ram_block3a4.port_b_last_address = 8191;
defparam ram_block3a4.port_b_logical_ram_depth = 16384;
defparam ram_block3a4.port_b_logical_ram_width = 32;
defparam ram_block3a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_read_enable_clock = "clock1";
defparam ram_block3a4.port_b_write_enable_clock = "clock1";
defparam ram_block3a4.ram_block_type = "M9K";
defparam ram_block3a4.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004F0080A;
// synopsys translate_on

// Location: M9K_X37_Y36_N0
cycloneive_ram_block ram_block3a37(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a37_PORTADATAOUT_bus),
	.portbdataout(ram_block3a37_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a37.clk0_core_clock_enable = "ena0";
defparam ram_block3a37.clk1_core_clock_enable = "ena1";
defparam ram_block3a37.data_interleave_offset_in_bits = 1;
defparam ram_block3a37.data_interleave_width_in_bits = 1;
defparam ram_block3a37.init_file = "meminit.hex";
defparam ram_block3a37.init_file_layout = "port_a";
defparam ram_block3a37.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a37.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a37.operation_mode = "bidir_dual_port";
defparam ram_block3a37.port_a_address_clear = "none";
defparam ram_block3a37.port_a_address_width = 13;
defparam ram_block3a37.port_a_byte_enable_clock = "none";
defparam ram_block3a37.port_a_data_out_clear = "none";
defparam ram_block3a37.port_a_data_out_clock = "none";
defparam ram_block3a37.port_a_data_width = 1;
defparam ram_block3a37.port_a_first_address = 0;
defparam ram_block3a37.port_a_first_bit_number = 5;
defparam ram_block3a37.port_a_last_address = 8191;
defparam ram_block3a37.port_a_logical_ram_depth = 16384;
defparam ram_block3a37.port_a_logical_ram_width = 32;
defparam ram_block3a37.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_address_clear = "none";
defparam ram_block3a37.port_b_address_clock = "clock1";
defparam ram_block3a37.port_b_address_width = 13;
defparam ram_block3a37.port_b_data_in_clock = "clock1";
defparam ram_block3a37.port_b_data_out_clear = "none";
defparam ram_block3a37.port_b_data_out_clock = "none";
defparam ram_block3a37.port_b_data_width = 1;
defparam ram_block3a37.port_b_first_address = 0;
defparam ram_block3a37.port_b_first_bit_number = 5;
defparam ram_block3a37.port_b_last_address = 8191;
defparam ram_block3a37.port_b_logical_ram_depth = 16384;
defparam ram_block3a37.port_b_logical_ram_width = 32;
defparam ram_block3a37.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_read_enable_clock = "clock1";
defparam ram_block3a37.port_b_write_enable_clock = "clock1";
defparam ram_block3a37.ram_block_type = "M9K";
defparam ram_block3a37.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y23_N0
cycloneive_ram_block ram_block3a5(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a5_PORTADATAOUT_bus),
	.portbdataout(ram_block3a5_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a5.clk0_core_clock_enable = "ena0";
defparam ram_block3a5.clk1_core_clock_enable = "ena1";
defparam ram_block3a5.data_interleave_offset_in_bits = 1;
defparam ram_block3a5.data_interleave_width_in_bits = 1;
defparam ram_block3a5.init_file = "meminit.hex";
defparam ram_block3a5.init_file_layout = "port_a";
defparam ram_block3a5.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a5.operation_mode = "bidir_dual_port";
defparam ram_block3a5.port_a_address_clear = "none";
defparam ram_block3a5.port_a_address_width = 13;
defparam ram_block3a5.port_a_byte_enable_clock = "none";
defparam ram_block3a5.port_a_data_out_clear = "none";
defparam ram_block3a5.port_a_data_out_clock = "none";
defparam ram_block3a5.port_a_data_width = 1;
defparam ram_block3a5.port_a_first_address = 0;
defparam ram_block3a5.port_a_first_bit_number = 5;
defparam ram_block3a5.port_a_last_address = 8191;
defparam ram_block3a5.port_a_logical_ram_depth = 16384;
defparam ram_block3a5.port_a_logical_ram_width = 32;
defparam ram_block3a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_address_clear = "none";
defparam ram_block3a5.port_b_address_clock = "clock1";
defparam ram_block3a5.port_b_address_width = 13;
defparam ram_block3a5.port_b_data_in_clock = "clock1";
defparam ram_block3a5.port_b_data_out_clear = "none";
defparam ram_block3a5.port_b_data_out_clock = "none";
defparam ram_block3a5.port_b_data_width = 1;
defparam ram_block3a5.port_b_first_address = 0;
defparam ram_block3a5.port_b_first_bit_number = 5;
defparam ram_block3a5.port_b_last_address = 8191;
defparam ram_block3a5.port_b_logical_ram_depth = 16384;
defparam ram_block3a5.port_b_logical_ram_width = 32;
defparam ram_block3a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_read_enable_clock = "clock1";
defparam ram_block3a5.port_b_write_enable_clock = "clock1";
defparam ram_block3a5.ram_block_type = "M9K";
defparam ram_block3a5.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007004EBB;
// synopsys translate_on

// Location: M9K_X37_Y32_N0
cycloneive_ram_block ram_block3a38(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a38_PORTADATAOUT_bus),
	.portbdataout(ram_block3a38_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a38.clk0_core_clock_enable = "ena0";
defparam ram_block3a38.clk1_core_clock_enable = "ena1";
defparam ram_block3a38.data_interleave_offset_in_bits = 1;
defparam ram_block3a38.data_interleave_width_in_bits = 1;
defparam ram_block3a38.init_file = "meminit.hex";
defparam ram_block3a38.init_file_layout = "port_a";
defparam ram_block3a38.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a38.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a38.operation_mode = "bidir_dual_port";
defparam ram_block3a38.port_a_address_clear = "none";
defparam ram_block3a38.port_a_address_width = 13;
defparam ram_block3a38.port_a_byte_enable_clock = "none";
defparam ram_block3a38.port_a_data_out_clear = "none";
defparam ram_block3a38.port_a_data_out_clock = "none";
defparam ram_block3a38.port_a_data_width = 1;
defparam ram_block3a38.port_a_first_address = 0;
defparam ram_block3a38.port_a_first_bit_number = 6;
defparam ram_block3a38.port_a_last_address = 8191;
defparam ram_block3a38.port_a_logical_ram_depth = 16384;
defparam ram_block3a38.port_a_logical_ram_width = 32;
defparam ram_block3a38.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_address_clear = "none";
defparam ram_block3a38.port_b_address_clock = "clock1";
defparam ram_block3a38.port_b_address_width = 13;
defparam ram_block3a38.port_b_data_in_clock = "clock1";
defparam ram_block3a38.port_b_data_out_clear = "none";
defparam ram_block3a38.port_b_data_out_clock = "none";
defparam ram_block3a38.port_b_data_width = 1;
defparam ram_block3a38.port_b_first_address = 0;
defparam ram_block3a38.port_b_first_bit_number = 6;
defparam ram_block3a38.port_b_last_address = 8191;
defparam ram_block3a38.port_b_logical_ram_depth = 16384;
defparam ram_block3a38.port_b_logical_ram_width = 32;
defparam ram_block3a38.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_read_enable_clock = "clock1";
defparam ram_block3a38.port_b_write_enable_clock = "clock1";
defparam ram_block3a38.ram_block_type = "M9K";
defparam ram_block3a38.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y33_N0
cycloneive_ram_block ram_block3a6(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a6_PORTADATAOUT_bus),
	.portbdataout(ram_block3a6_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a6.clk0_core_clock_enable = "ena0";
defparam ram_block3a6.clk1_core_clock_enable = "ena1";
defparam ram_block3a6.data_interleave_offset_in_bits = 1;
defparam ram_block3a6.data_interleave_width_in_bits = 1;
defparam ram_block3a6.init_file = "meminit.hex";
defparam ram_block3a6.init_file_layout = "port_a";
defparam ram_block3a6.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a6.operation_mode = "bidir_dual_port";
defparam ram_block3a6.port_a_address_clear = "none";
defparam ram_block3a6.port_a_address_width = 13;
defparam ram_block3a6.port_a_byte_enable_clock = "none";
defparam ram_block3a6.port_a_data_out_clear = "none";
defparam ram_block3a6.port_a_data_out_clock = "none";
defparam ram_block3a6.port_a_data_width = 1;
defparam ram_block3a6.port_a_first_address = 0;
defparam ram_block3a6.port_a_first_bit_number = 6;
defparam ram_block3a6.port_a_last_address = 8191;
defparam ram_block3a6.port_a_logical_ram_depth = 16384;
defparam ram_block3a6.port_a_logical_ram_width = 32;
defparam ram_block3a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_address_clear = "none";
defparam ram_block3a6.port_b_address_clock = "clock1";
defparam ram_block3a6.port_b_address_width = 13;
defparam ram_block3a6.port_b_data_in_clock = "clock1";
defparam ram_block3a6.port_b_data_out_clear = "none";
defparam ram_block3a6.port_b_data_out_clock = "none";
defparam ram_block3a6.port_b_data_width = 1;
defparam ram_block3a6.port_b_first_address = 0;
defparam ram_block3a6.port_b_first_bit_number = 6;
defparam ram_block3a6.port_b_last_address = 8191;
defparam ram_block3a6.port_b_logical_ram_depth = 16384;
defparam ram_block3a6.port_b_logical_ram_width = 32;
defparam ram_block3a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_read_enable_clock = "clock1";
defparam ram_block3a6.port_b_write_enable_clock = "clock1";
defparam ram_block3a6.ram_block_type = "M9K";
defparam ram_block3a6.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000400210B;
// synopsys translate_on

// Location: M9K_X51_Y29_N0
cycloneive_ram_block ram_block3a39(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a39_PORTADATAOUT_bus),
	.portbdataout(ram_block3a39_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a39.clk0_core_clock_enable = "ena0";
defparam ram_block3a39.clk1_core_clock_enable = "ena1";
defparam ram_block3a39.data_interleave_offset_in_bits = 1;
defparam ram_block3a39.data_interleave_width_in_bits = 1;
defparam ram_block3a39.init_file = "meminit.hex";
defparam ram_block3a39.init_file_layout = "port_a";
defparam ram_block3a39.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a39.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a39.operation_mode = "bidir_dual_port";
defparam ram_block3a39.port_a_address_clear = "none";
defparam ram_block3a39.port_a_address_width = 13;
defparam ram_block3a39.port_a_byte_enable_clock = "none";
defparam ram_block3a39.port_a_data_out_clear = "none";
defparam ram_block3a39.port_a_data_out_clock = "none";
defparam ram_block3a39.port_a_data_width = 1;
defparam ram_block3a39.port_a_first_address = 0;
defparam ram_block3a39.port_a_first_bit_number = 7;
defparam ram_block3a39.port_a_last_address = 8191;
defparam ram_block3a39.port_a_logical_ram_depth = 16384;
defparam ram_block3a39.port_a_logical_ram_width = 32;
defparam ram_block3a39.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_address_clear = "none";
defparam ram_block3a39.port_b_address_clock = "clock1";
defparam ram_block3a39.port_b_address_width = 13;
defparam ram_block3a39.port_b_data_in_clock = "clock1";
defparam ram_block3a39.port_b_data_out_clear = "none";
defparam ram_block3a39.port_b_data_out_clock = "none";
defparam ram_block3a39.port_b_data_width = 1;
defparam ram_block3a39.port_b_first_address = 0;
defparam ram_block3a39.port_b_first_bit_number = 7;
defparam ram_block3a39.port_b_last_address = 8191;
defparam ram_block3a39.port_b_logical_ram_depth = 16384;
defparam ram_block3a39.port_b_logical_ram_width = 32;
defparam ram_block3a39.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_read_enable_clock = "clock1";
defparam ram_block3a39.port_b_write_enable_clock = "clock1";
defparam ram_block3a39.ram_block_type = "M9K";
defparam ram_block3a39.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y32_N0
cycloneive_ram_block ram_block3a7(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a7_PORTADATAOUT_bus),
	.portbdataout(ram_block3a7_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a7.clk0_core_clock_enable = "ena0";
defparam ram_block3a7.clk1_core_clock_enable = "ena1";
defparam ram_block3a7.data_interleave_offset_in_bits = 1;
defparam ram_block3a7.data_interleave_width_in_bits = 1;
defparam ram_block3a7.init_file = "meminit.hex";
defparam ram_block3a7.init_file_layout = "port_a";
defparam ram_block3a7.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a7.operation_mode = "bidir_dual_port";
defparam ram_block3a7.port_a_address_clear = "none";
defparam ram_block3a7.port_a_address_width = 13;
defparam ram_block3a7.port_a_byte_enable_clock = "none";
defparam ram_block3a7.port_a_data_out_clear = "none";
defparam ram_block3a7.port_a_data_out_clock = "none";
defparam ram_block3a7.port_a_data_width = 1;
defparam ram_block3a7.port_a_first_address = 0;
defparam ram_block3a7.port_a_first_bit_number = 7;
defparam ram_block3a7.port_a_last_address = 8191;
defparam ram_block3a7.port_a_logical_ram_depth = 16384;
defparam ram_block3a7.port_a_logical_ram_width = 32;
defparam ram_block3a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_address_clear = "none";
defparam ram_block3a7.port_b_address_clock = "clock1";
defparam ram_block3a7.port_b_address_width = 13;
defparam ram_block3a7.port_b_data_in_clock = "clock1";
defparam ram_block3a7.port_b_data_out_clear = "none";
defparam ram_block3a7.port_b_data_out_clock = "none";
defparam ram_block3a7.port_b_data_width = 1;
defparam ram_block3a7.port_b_first_address = 0;
defparam ram_block3a7.port_b_first_bit_number = 7;
defparam ram_block3a7.port_b_last_address = 8191;
defparam ram_block3a7.port_b_logical_ram_depth = 16384;
defparam ram_block3a7.port_b_logical_ram_width = 32;
defparam ram_block3a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_read_enable_clock = "clock1";
defparam ram_block3a7.port_b_write_enable_clock = "clock1";
defparam ram_block3a7.ram_block_type = "M9K";
defparam ram_block3a7.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000400000E;
// synopsys translate_on

// Location: M9K_X78_Y32_N0
cycloneive_ram_block ram_block3a40(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a40_PORTADATAOUT_bus),
	.portbdataout(ram_block3a40_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a40.clk0_core_clock_enable = "ena0";
defparam ram_block3a40.clk1_core_clock_enable = "ena1";
defparam ram_block3a40.data_interleave_offset_in_bits = 1;
defparam ram_block3a40.data_interleave_width_in_bits = 1;
defparam ram_block3a40.init_file = "meminit.hex";
defparam ram_block3a40.init_file_layout = "port_a";
defparam ram_block3a40.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a40.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a40.operation_mode = "bidir_dual_port";
defparam ram_block3a40.port_a_address_clear = "none";
defparam ram_block3a40.port_a_address_width = 13;
defparam ram_block3a40.port_a_byte_enable_clock = "none";
defparam ram_block3a40.port_a_data_out_clear = "none";
defparam ram_block3a40.port_a_data_out_clock = "none";
defparam ram_block3a40.port_a_data_width = 1;
defparam ram_block3a40.port_a_first_address = 0;
defparam ram_block3a40.port_a_first_bit_number = 8;
defparam ram_block3a40.port_a_last_address = 8191;
defparam ram_block3a40.port_a_logical_ram_depth = 16384;
defparam ram_block3a40.port_a_logical_ram_width = 32;
defparam ram_block3a40.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_address_clear = "none";
defparam ram_block3a40.port_b_address_clock = "clock1";
defparam ram_block3a40.port_b_address_width = 13;
defparam ram_block3a40.port_b_data_in_clock = "clock1";
defparam ram_block3a40.port_b_data_out_clear = "none";
defparam ram_block3a40.port_b_data_out_clock = "none";
defparam ram_block3a40.port_b_data_width = 1;
defparam ram_block3a40.port_b_first_address = 0;
defparam ram_block3a40.port_b_first_bit_number = 8;
defparam ram_block3a40.port_b_last_address = 8191;
defparam ram_block3a40.port_b_logical_ram_depth = 16384;
defparam ram_block3a40.port_b_logical_ram_width = 32;
defparam ram_block3a40.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_read_enable_clock = "clock1";
defparam ram_block3a40.port_b_write_enable_clock = "clock1";
defparam ram_block3a40.ram_block_type = "M9K";
defparam ram_block3a40.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y43_N0
cycloneive_ram_block ram_block3a8(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a8_PORTADATAOUT_bus),
	.portbdataout(ram_block3a8_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a8.clk0_core_clock_enable = "ena0";
defparam ram_block3a8.clk1_core_clock_enable = "ena1";
defparam ram_block3a8.data_interleave_offset_in_bits = 1;
defparam ram_block3a8.data_interleave_width_in_bits = 1;
defparam ram_block3a8.init_file = "meminit.hex";
defparam ram_block3a8.init_file_layout = "port_a";
defparam ram_block3a8.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a8.operation_mode = "bidir_dual_port";
defparam ram_block3a8.port_a_address_clear = "none";
defparam ram_block3a8.port_a_address_width = 13;
defparam ram_block3a8.port_a_byte_enable_clock = "none";
defparam ram_block3a8.port_a_data_out_clear = "none";
defparam ram_block3a8.port_a_data_out_clock = "none";
defparam ram_block3a8.port_a_data_width = 1;
defparam ram_block3a8.port_a_first_address = 0;
defparam ram_block3a8.port_a_first_bit_number = 8;
defparam ram_block3a8.port_a_last_address = 8191;
defparam ram_block3a8.port_a_logical_ram_depth = 16384;
defparam ram_block3a8.port_a_logical_ram_width = 32;
defparam ram_block3a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_address_clear = "none";
defparam ram_block3a8.port_b_address_clock = "clock1";
defparam ram_block3a8.port_b_address_width = 13;
defparam ram_block3a8.port_b_data_in_clock = "clock1";
defparam ram_block3a8.port_b_data_out_clear = "none";
defparam ram_block3a8.port_b_data_out_clock = "none";
defparam ram_block3a8.port_b_data_width = 1;
defparam ram_block3a8.port_b_first_address = 0;
defparam ram_block3a8.port_b_first_bit_number = 8;
defparam ram_block3a8.port_b_last_address = 8191;
defparam ram_block3a8.port_b_logical_ram_depth = 16384;
defparam ram_block3a8.port_b_logical_ram_width = 32;
defparam ram_block3a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_read_enable_clock = "clock1";
defparam ram_block3a8.port_b_write_enable_clock = "clock1";
defparam ram_block3a8.ram_block_type = "M9K";
defparam ram_block3a8.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004003902;
// synopsys translate_on

// Location: M9K_X51_Y24_N0
cycloneive_ram_block ram_block3a41(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a41_PORTADATAOUT_bus),
	.portbdataout(ram_block3a41_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a41.clk0_core_clock_enable = "ena0";
defparam ram_block3a41.clk1_core_clock_enable = "ena1";
defparam ram_block3a41.data_interleave_offset_in_bits = 1;
defparam ram_block3a41.data_interleave_width_in_bits = 1;
defparam ram_block3a41.init_file = "meminit.hex";
defparam ram_block3a41.init_file_layout = "port_a";
defparam ram_block3a41.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a41.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a41.operation_mode = "bidir_dual_port";
defparam ram_block3a41.port_a_address_clear = "none";
defparam ram_block3a41.port_a_address_width = 13;
defparam ram_block3a41.port_a_byte_enable_clock = "none";
defparam ram_block3a41.port_a_data_out_clear = "none";
defparam ram_block3a41.port_a_data_out_clock = "none";
defparam ram_block3a41.port_a_data_width = 1;
defparam ram_block3a41.port_a_first_address = 0;
defparam ram_block3a41.port_a_first_bit_number = 9;
defparam ram_block3a41.port_a_last_address = 8191;
defparam ram_block3a41.port_a_logical_ram_depth = 16384;
defparam ram_block3a41.port_a_logical_ram_width = 32;
defparam ram_block3a41.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_address_clear = "none";
defparam ram_block3a41.port_b_address_clock = "clock1";
defparam ram_block3a41.port_b_address_width = 13;
defparam ram_block3a41.port_b_data_in_clock = "clock1";
defparam ram_block3a41.port_b_data_out_clear = "none";
defparam ram_block3a41.port_b_data_out_clock = "none";
defparam ram_block3a41.port_b_data_width = 1;
defparam ram_block3a41.port_b_first_address = 0;
defparam ram_block3a41.port_b_first_bit_number = 9;
defparam ram_block3a41.port_b_last_address = 8191;
defparam ram_block3a41.port_b_logical_ram_depth = 16384;
defparam ram_block3a41.port_b_logical_ram_width = 32;
defparam ram_block3a41.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_read_enable_clock = "clock1";
defparam ram_block3a41.port_b_write_enable_clock = "clock1";
defparam ram_block3a41.ram_block_type = "M9K";
defparam ram_block3a41.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y28_N0
cycloneive_ram_block ram_block3a9(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a9_PORTADATAOUT_bus),
	.portbdataout(ram_block3a9_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a9.clk0_core_clock_enable = "ena0";
defparam ram_block3a9.clk1_core_clock_enable = "ena1";
defparam ram_block3a9.data_interleave_offset_in_bits = 1;
defparam ram_block3a9.data_interleave_width_in_bits = 1;
defparam ram_block3a9.init_file = "meminit.hex";
defparam ram_block3a9.init_file_layout = "port_a";
defparam ram_block3a9.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a9.operation_mode = "bidir_dual_port";
defparam ram_block3a9.port_a_address_clear = "none";
defparam ram_block3a9.port_a_address_width = 13;
defparam ram_block3a9.port_a_byte_enable_clock = "none";
defparam ram_block3a9.port_a_data_out_clear = "none";
defparam ram_block3a9.port_a_data_out_clock = "none";
defparam ram_block3a9.port_a_data_width = 1;
defparam ram_block3a9.port_a_first_address = 0;
defparam ram_block3a9.port_a_first_bit_number = 9;
defparam ram_block3a9.port_a_last_address = 8191;
defparam ram_block3a9.port_a_logical_ram_depth = 16384;
defparam ram_block3a9.port_a_logical_ram_width = 32;
defparam ram_block3a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_address_clear = "none";
defparam ram_block3a9.port_b_address_clock = "clock1";
defparam ram_block3a9.port_b_address_width = 13;
defparam ram_block3a9.port_b_data_in_clock = "clock1";
defparam ram_block3a9.port_b_data_out_clear = "none";
defparam ram_block3a9.port_b_data_out_clock = "none";
defparam ram_block3a9.port_b_data_width = 1;
defparam ram_block3a9.port_b_first_address = 0;
defparam ram_block3a9.port_b_first_bit_number = 9;
defparam ram_block3a9.port_b_last_address = 8191;
defparam ram_block3a9.port_b_logical_ram_depth = 16384;
defparam ram_block3a9.port_b_logical_ram_width = 32;
defparam ram_block3a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_read_enable_clock = "clock1";
defparam ram_block3a9.port_b_write_enable_clock = "clock1";
defparam ram_block3a9.ram_block_type = "M9K";
defparam ram_block3a9.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004000903;
// synopsys translate_on

// Location: M9K_X64_Y39_N0
cycloneive_ram_block ram_block3a42(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a42_PORTADATAOUT_bus),
	.portbdataout(ram_block3a42_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a42.clk0_core_clock_enable = "ena0";
defparam ram_block3a42.clk1_core_clock_enable = "ena1";
defparam ram_block3a42.data_interleave_offset_in_bits = 1;
defparam ram_block3a42.data_interleave_width_in_bits = 1;
defparam ram_block3a42.init_file = "meminit.hex";
defparam ram_block3a42.init_file_layout = "port_a";
defparam ram_block3a42.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a42.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a42.operation_mode = "bidir_dual_port";
defparam ram_block3a42.port_a_address_clear = "none";
defparam ram_block3a42.port_a_address_width = 13;
defparam ram_block3a42.port_a_byte_enable_clock = "none";
defparam ram_block3a42.port_a_data_out_clear = "none";
defparam ram_block3a42.port_a_data_out_clock = "none";
defparam ram_block3a42.port_a_data_width = 1;
defparam ram_block3a42.port_a_first_address = 0;
defparam ram_block3a42.port_a_first_bit_number = 10;
defparam ram_block3a42.port_a_last_address = 8191;
defparam ram_block3a42.port_a_logical_ram_depth = 16384;
defparam ram_block3a42.port_a_logical_ram_width = 32;
defparam ram_block3a42.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_address_clear = "none";
defparam ram_block3a42.port_b_address_clock = "clock1";
defparam ram_block3a42.port_b_address_width = 13;
defparam ram_block3a42.port_b_data_in_clock = "clock1";
defparam ram_block3a42.port_b_data_out_clear = "none";
defparam ram_block3a42.port_b_data_out_clock = "none";
defparam ram_block3a42.port_b_data_width = 1;
defparam ram_block3a42.port_b_first_address = 0;
defparam ram_block3a42.port_b_first_bit_number = 10;
defparam ram_block3a42.port_b_last_address = 8191;
defparam ram_block3a42.port_b_logical_ram_depth = 16384;
defparam ram_block3a42.port_b_logical_ram_width = 32;
defparam ram_block3a42.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_read_enable_clock = "clock1";
defparam ram_block3a42.port_b_write_enable_clock = "clock1";
defparam ram_block3a42.ram_block_type = "M9K";
defparam ram_block3a42.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y38_N0
cycloneive_ram_block ram_block3a10(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a10_PORTADATAOUT_bus),
	.portbdataout(ram_block3a10_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a10.clk0_core_clock_enable = "ena0";
defparam ram_block3a10.clk1_core_clock_enable = "ena1";
defparam ram_block3a10.data_interleave_offset_in_bits = 1;
defparam ram_block3a10.data_interleave_width_in_bits = 1;
defparam ram_block3a10.init_file = "meminit.hex";
defparam ram_block3a10.init_file_layout = "port_a";
defparam ram_block3a10.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a10.operation_mode = "bidir_dual_port";
defparam ram_block3a10.port_a_address_clear = "none";
defparam ram_block3a10.port_a_address_width = 13;
defparam ram_block3a10.port_a_byte_enable_clock = "none";
defparam ram_block3a10.port_a_data_out_clear = "none";
defparam ram_block3a10.port_a_data_out_clock = "none";
defparam ram_block3a10.port_a_data_width = 1;
defparam ram_block3a10.port_a_first_address = 0;
defparam ram_block3a10.port_a_first_bit_number = 10;
defparam ram_block3a10.port_a_last_address = 8191;
defparam ram_block3a10.port_a_logical_ram_depth = 16384;
defparam ram_block3a10.port_a_logical_ram_width = 32;
defparam ram_block3a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_address_clear = "none";
defparam ram_block3a10.port_b_address_clock = "clock1";
defparam ram_block3a10.port_b_address_width = 13;
defparam ram_block3a10.port_b_data_in_clock = "clock1";
defparam ram_block3a10.port_b_data_out_clear = "none";
defparam ram_block3a10.port_b_data_out_clock = "none";
defparam ram_block3a10.port_b_data_width = 1;
defparam ram_block3a10.port_b_first_address = 0;
defparam ram_block3a10.port_b_first_bit_number = 10;
defparam ram_block3a10.port_b_last_address = 8191;
defparam ram_block3a10.port_b_logical_ram_depth = 16384;
defparam ram_block3a10.port_b_logical_ram_width = 32;
defparam ram_block3a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_read_enable_clock = "clock1";
defparam ram_block3a10.port_b_write_enable_clock = "clock1";
defparam ram_block3a10.ram_block_type = "M9K";
defparam ram_block3a10.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004000102;
// synopsys translate_on

// Location: M9K_X78_Y35_N0
cycloneive_ram_block ram_block3a43(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a43_PORTADATAOUT_bus),
	.portbdataout(ram_block3a43_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a43.clk0_core_clock_enable = "ena0";
defparam ram_block3a43.clk1_core_clock_enable = "ena1";
defparam ram_block3a43.data_interleave_offset_in_bits = 1;
defparam ram_block3a43.data_interleave_width_in_bits = 1;
defparam ram_block3a43.init_file = "meminit.hex";
defparam ram_block3a43.init_file_layout = "port_a";
defparam ram_block3a43.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a43.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a43.operation_mode = "bidir_dual_port";
defparam ram_block3a43.port_a_address_clear = "none";
defparam ram_block3a43.port_a_address_width = 13;
defparam ram_block3a43.port_a_byte_enable_clock = "none";
defparam ram_block3a43.port_a_data_out_clear = "none";
defparam ram_block3a43.port_a_data_out_clock = "none";
defparam ram_block3a43.port_a_data_width = 1;
defparam ram_block3a43.port_a_first_address = 0;
defparam ram_block3a43.port_a_first_bit_number = 11;
defparam ram_block3a43.port_a_last_address = 8191;
defparam ram_block3a43.port_a_logical_ram_depth = 16384;
defparam ram_block3a43.port_a_logical_ram_width = 32;
defparam ram_block3a43.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_address_clear = "none";
defparam ram_block3a43.port_b_address_clock = "clock1";
defparam ram_block3a43.port_b_address_width = 13;
defparam ram_block3a43.port_b_data_in_clock = "clock1";
defparam ram_block3a43.port_b_data_out_clear = "none";
defparam ram_block3a43.port_b_data_out_clock = "none";
defparam ram_block3a43.port_b_data_width = 1;
defparam ram_block3a43.port_b_first_address = 0;
defparam ram_block3a43.port_b_first_bit_number = 11;
defparam ram_block3a43.port_b_last_address = 8191;
defparam ram_block3a43.port_b_logical_ram_depth = 16384;
defparam ram_block3a43.port_b_logical_ram_width = 32;
defparam ram_block3a43.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_read_enable_clock = "clock1";
defparam ram_block3a43.port_b_write_enable_clock = "clock1";
defparam ram_block3a43.ram_block_type = "M9K";
defparam ram_block3a43.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y35_N0
cycloneive_ram_block ram_block3a11(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a11_PORTADATAOUT_bus),
	.portbdataout(ram_block3a11_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a11.clk0_core_clock_enable = "ena0";
defparam ram_block3a11.clk1_core_clock_enable = "ena1";
defparam ram_block3a11.data_interleave_offset_in_bits = 1;
defparam ram_block3a11.data_interleave_width_in_bits = 1;
defparam ram_block3a11.init_file = "meminit.hex";
defparam ram_block3a11.init_file_layout = "port_a";
defparam ram_block3a11.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a11.operation_mode = "bidir_dual_port";
defparam ram_block3a11.port_a_address_clear = "none";
defparam ram_block3a11.port_a_address_width = 13;
defparam ram_block3a11.port_a_byte_enable_clock = "none";
defparam ram_block3a11.port_a_data_out_clear = "none";
defparam ram_block3a11.port_a_data_out_clock = "none";
defparam ram_block3a11.port_a_data_width = 1;
defparam ram_block3a11.port_a_first_address = 0;
defparam ram_block3a11.port_a_first_bit_number = 11;
defparam ram_block3a11.port_a_last_address = 8191;
defparam ram_block3a11.port_a_logical_ram_depth = 16384;
defparam ram_block3a11.port_a_logical_ram_width = 32;
defparam ram_block3a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_address_clear = "none";
defparam ram_block3a11.port_b_address_clock = "clock1";
defparam ram_block3a11.port_b_address_width = 13;
defparam ram_block3a11.port_b_data_in_clock = "clock1";
defparam ram_block3a11.port_b_data_out_clear = "none";
defparam ram_block3a11.port_b_data_out_clock = "none";
defparam ram_block3a11.port_b_data_width = 1;
defparam ram_block3a11.port_b_first_address = 0;
defparam ram_block3a11.port_b_first_bit_number = 11;
defparam ram_block3a11.port_b_last_address = 8191;
defparam ram_block3a11.port_b_logical_ram_depth = 16384;
defparam ram_block3a11.port_b_logical_ram_width = 32;
defparam ram_block3a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_read_enable_clock = "clock1";
defparam ram_block3a11.port_b_write_enable_clock = "clock1";
defparam ram_block3a11.ram_block_type = "M9K";
defparam ram_block3a11.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004005410;
// synopsys translate_on

// Location: M9K_X64_Y37_N0
cycloneive_ram_block ram_block3a44(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a44_PORTADATAOUT_bus),
	.portbdataout(ram_block3a44_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a44.clk0_core_clock_enable = "ena0";
defparam ram_block3a44.clk1_core_clock_enable = "ena1";
defparam ram_block3a44.data_interleave_offset_in_bits = 1;
defparam ram_block3a44.data_interleave_width_in_bits = 1;
defparam ram_block3a44.init_file = "meminit.hex";
defparam ram_block3a44.init_file_layout = "port_a";
defparam ram_block3a44.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a44.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a44.operation_mode = "bidir_dual_port";
defparam ram_block3a44.port_a_address_clear = "none";
defparam ram_block3a44.port_a_address_width = 13;
defparam ram_block3a44.port_a_byte_enable_clock = "none";
defparam ram_block3a44.port_a_data_out_clear = "none";
defparam ram_block3a44.port_a_data_out_clock = "none";
defparam ram_block3a44.port_a_data_width = 1;
defparam ram_block3a44.port_a_first_address = 0;
defparam ram_block3a44.port_a_first_bit_number = 12;
defparam ram_block3a44.port_a_last_address = 8191;
defparam ram_block3a44.port_a_logical_ram_depth = 16384;
defparam ram_block3a44.port_a_logical_ram_width = 32;
defparam ram_block3a44.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_address_clear = "none";
defparam ram_block3a44.port_b_address_clock = "clock1";
defparam ram_block3a44.port_b_address_width = 13;
defparam ram_block3a44.port_b_data_in_clock = "clock1";
defparam ram_block3a44.port_b_data_out_clear = "none";
defparam ram_block3a44.port_b_data_out_clock = "none";
defparam ram_block3a44.port_b_data_width = 1;
defparam ram_block3a44.port_b_first_address = 0;
defparam ram_block3a44.port_b_first_bit_number = 12;
defparam ram_block3a44.port_b_last_address = 8191;
defparam ram_block3a44.port_b_logical_ram_depth = 16384;
defparam ram_block3a44.port_b_logical_ram_width = 32;
defparam ram_block3a44.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_read_enable_clock = "clock1";
defparam ram_block3a44.port_b_write_enable_clock = "clock1";
defparam ram_block3a44.ram_block_type = "M9K";
defparam ram_block3a44.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y30_N0
cycloneive_ram_block ram_block3a12(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a12_PORTADATAOUT_bus),
	.portbdataout(ram_block3a12_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a12.clk0_core_clock_enable = "ena0";
defparam ram_block3a12.clk1_core_clock_enable = "ena1";
defparam ram_block3a12.data_interleave_offset_in_bits = 1;
defparam ram_block3a12.data_interleave_width_in_bits = 1;
defparam ram_block3a12.init_file = "meminit.hex";
defparam ram_block3a12.init_file_layout = "port_a";
defparam ram_block3a12.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a12.operation_mode = "bidir_dual_port";
defparam ram_block3a12.port_a_address_clear = "none";
defparam ram_block3a12.port_a_address_width = 13;
defparam ram_block3a12.port_a_byte_enable_clock = "none";
defparam ram_block3a12.port_a_data_out_clear = "none";
defparam ram_block3a12.port_a_data_out_clock = "none";
defparam ram_block3a12.port_a_data_width = 1;
defparam ram_block3a12.port_a_first_address = 0;
defparam ram_block3a12.port_a_first_bit_number = 12;
defparam ram_block3a12.port_a_last_address = 8191;
defparam ram_block3a12.port_a_logical_ram_depth = 16384;
defparam ram_block3a12.port_a_logical_ram_width = 32;
defparam ram_block3a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_address_clear = "none";
defparam ram_block3a12.port_b_address_clock = "clock1";
defparam ram_block3a12.port_b_address_width = 13;
defparam ram_block3a12.port_b_data_in_clock = "clock1";
defparam ram_block3a12.port_b_data_out_clear = "none";
defparam ram_block3a12.port_b_data_out_clock = "none";
defparam ram_block3a12.port_b_data_width = 1;
defparam ram_block3a12.port_b_first_address = 0;
defparam ram_block3a12.port_b_first_bit_number = 12;
defparam ram_block3a12.port_b_last_address = 8191;
defparam ram_block3a12.port_b_logical_ram_depth = 16384;
defparam ram_block3a12.port_b_logical_ram_width = 32;
defparam ram_block3a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_read_enable_clock = "clock1";
defparam ram_block3a12.port_b_write_enable_clock = "clock1";
defparam ram_block3a12.ram_block_type = "M9K";
defparam ram_block3a12.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004001893;
// synopsys translate_on

// Location: M9K_X64_Y24_N0
cycloneive_ram_block ram_block3a45(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a45_PORTADATAOUT_bus),
	.portbdataout(ram_block3a45_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a45.clk0_core_clock_enable = "ena0";
defparam ram_block3a45.clk1_core_clock_enable = "ena1";
defparam ram_block3a45.data_interleave_offset_in_bits = 1;
defparam ram_block3a45.data_interleave_width_in_bits = 1;
defparam ram_block3a45.init_file = "meminit.hex";
defparam ram_block3a45.init_file_layout = "port_a";
defparam ram_block3a45.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a45.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a45.operation_mode = "bidir_dual_port";
defparam ram_block3a45.port_a_address_clear = "none";
defparam ram_block3a45.port_a_address_width = 13;
defparam ram_block3a45.port_a_byte_enable_clock = "none";
defparam ram_block3a45.port_a_data_out_clear = "none";
defparam ram_block3a45.port_a_data_out_clock = "none";
defparam ram_block3a45.port_a_data_width = 1;
defparam ram_block3a45.port_a_first_address = 0;
defparam ram_block3a45.port_a_first_bit_number = 13;
defparam ram_block3a45.port_a_last_address = 8191;
defparam ram_block3a45.port_a_logical_ram_depth = 16384;
defparam ram_block3a45.port_a_logical_ram_width = 32;
defparam ram_block3a45.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_address_clear = "none";
defparam ram_block3a45.port_b_address_clock = "clock1";
defparam ram_block3a45.port_b_address_width = 13;
defparam ram_block3a45.port_b_data_in_clock = "clock1";
defparam ram_block3a45.port_b_data_out_clear = "none";
defparam ram_block3a45.port_b_data_out_clock = "none";
defparam ram_block3a45.port_b_data_width = 1;
defparam ram_block3a45.port_b_first_address = 0;
defparam ram_block3a45.port_b_first_bit_number = 13;
defparam ram_block3a45.port_b_last_address = 8191;
defparam ram_block3a45.port_b_logical_ram_depth = 16384;
defparam ram_block3a45.port_b_logical_ram_width = 32;
defparam ram_block3a45.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_read_enable_clock = "clock1";
defparam ram_block3a45.port_b_write_enable_clock = "clock1";
defparam ram_block3a45.ram_block_type = "M9K";
defparam ram_block3a45.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y27_N0
cycloneive_ram_block ram_block3a13(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a13_PORTADATAOUT_bus),
	.portbdataout(ram_block3a13_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a13.clk0_core_clock_enable = "ena0";
defparam ram_block3a13.clk1_core_clock_enable = "ena1";
defparam ram_block3a13.data_interleave_offset_in_bits = 1;
defparam ram_block3a13.data_interleave_width_in_bits = 1;
defparam ram_block3a13.init_file = "meminit.hex";
defparam ram_block3a13.init_file_layout = "port_a";
defparam ram_block3a13.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a13.operation_mode = "bidir_dual_port";
defparam ram_block3a13.port_a_address_clear = "none";
defparam ram_block3a13.port_a_address_width = 13;
defparam ram_block3a13.port_a_byte_enable_clock = "none";
defparam ram_block3a13.port_a_data_out_clear = "none";
defparam ram_block3a13.port_a_data_out_clock = "none";
defparam ram_block3a13.port_a_data_width = 1;
defparam ram_block3a13.port_a_first_address = 0;
defparam ram_block3a13.port_a_first_bit_number = 13;
defparam ram_block3a13.port_a_last_address = 8191;
defparam ram_block3a13.port_a_logical_ram_depth = 16384;
defparam ram_block3a13.port_a_logical_ram_width = 32;
defparam ram_block3a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_address_clear = "none";
defparam ram_block3a13.port_b_address_clock = "clock1";
defparam ram_block3a13.port_b_address_width = 13;
defparam ram_block3a13.port_b_data_in_clock = "clock1";
defparam ram_block3a13.port_b_data_out_clear = "none";
defparam ram_block3a13.port_b_data_out_clock = "none";
defparam ram_block3a13.port_b_data_width = 1;
defparam ram_block3a13.port_b_first_address = 0;
defparam ram_block3a13.port_b_first_bit_number = 13;
defparam ram_block3a13.port_b_last_address = 8191;
defparam ram_block3a13.port_b_logical_ram_depth = 16384;
defparam ram_block3a13.port_b_logical_ram_width = 32;
defparam ram_block3a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_read_enable_clock = "clock1";
defparam ram_block3a13.port_b_write_enable_clock = "clock1";
defparam ram_block3a13.ram_block_type = "M9K";
defparam ram_block3a13.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000040068A2;
// synopsys translate_on

// Location: M9K_X51_Y28_N0
cycloneive_ram_block ram_block3a46(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a46_PORTADATAOUT_bus),
	.portbdataout(ram_block3a46_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a46.clk0_core_clock_enable = "ena0";
defparam ram_block3a46.clk1_core_clock_enable = "ena1";
defparam ram_block3a46.data_interleave_offset_in_bits = 1;
defparam ram_block3a46.data_interleave_width_in_bits = 1;
defparam ram_block3a46.init_file = "meminit.hex";
defparam ram_block3a46.init_file_layout = "port_a";
defparam ram_block3a46.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a46.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a46.operation_mode = "bidir_dual_port";
defparam ram_block3a46.port_a_address_clear = "none";
defparam ram_block3a46.port_a_address_width = 13;
defparam ram_block3a46.port_a_byte_enable_clock = "none";
defparam ram_block3a46.port_a_data_out_clear = "none";
defparam ram_block3a46.port_a_data_out_clock = "none";
defparam ram_block3a46.port_a_data_width = 1;
defparam ram_block3a46.port_a_first_address = 0;
defparam ram_block3a46.port_a_first_bit_number = 14;
defparam ram_block3a46.port_a_last_address = 8191;
defparam ram_block3a46.port_a_logical_ram_depth = 16384;
defparam ram_block3a46.port_a_logical_ram_width = 32;
defparam ram_block3a46.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_address_clear = "none";
defparam ram_block3a46.port_b_address_clock = "clock1";
defparam ram_block3a46.port_b_address_width = 13;
defparam ram_block3a46.port_b_data_in_clock = "clock1";
defparam ram_block3a46.port_b_data_out_clear = "none";
defparam ram_block3a46.port_b_data_out_clock = "none";
defparam ram_block3a46.port_b_data_width = 1;
defparam ram_block3a46.port_b_first_address = 0;
defparam ram_block3a46.port_b_first_bit_number = 14;
defparam ram_block3a46.port_b_last_address = 8191;
defparam ram_block3a46.port_b_logical_ram_depth = 16384;
defparam ram_block3a46.port_b_logical_ram_width = 32;
defparam ram_block3a46.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_read_enable_clock = "clock1";
defparam ram_block3a46.port_b_write_enable_clock = "clock1";
defparam ram_block3a46.ram_block_type = "M9K";
defparam ram_block3a46.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y21_N0
cycloneive_ram_block ram_block3a14(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a14_PORTADATAOUT_bus),
	.portbdataout(ram_block3a14_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a14.clk0_core_clock_enable = "ena0";
defparam ram_block3a14.clk1_core_clock_enable = "ena1";
defparam ram_block3a14.data_interleave_offset_in_bits = 1;
defparam ram_block3a14.data_interleave_width_in_bits = 1;
defparam ram_block3a14.init_file = "meminit.hex";
defparam ram_block3a14.init_file_layout = "port_a";
defparam ram_block3a14.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a14.operation_mode = "bidir_dual_port";
defparam ram_block3a14.port_a_address_clear = "none";
defparam ram_block3a14.port_a_address_width = 13;
defparam ram_block3a14.port_a_byte_enable_clock = "none";
defparam ram_block3a14.port_a_data_out_clear = "none";
defparam ram_block3a14.port_a_data_out_clock = "none";
defparam ram_block3a14.port_a_data_width = 1;
defparam ram_block3a14.port_a_first_address = 0;
defparam ram_block3a14.port_a_first_bit_number = 14;
defparam ram_block3a14.port_a_last_address = 8191;
defparam ram_block3a14.port_a_logical_ram_depth = 16384;
defparam ram_block3a14.port_a_logical_ram_width = 32;
defparam ram_block3a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_address_clear = "none";
defparam ram_block3a14.port_b_address_clock = "clock1";
defparam ram_block3a14.port_b_address_width = 13;
defparam ram_block3a14.port_b_data_in_clock = "clock1";
defparam ram_block3a14.port_b_data_out_clear = "none";
defparam ram_block3a14.port_b_data_out_clock = "none";
defparam ram_block3a14.port_b_data_width = 1;
defparam ram_block3a14.port_b_first_address = 0;
defparam ram_block3a14.port_b_first_bit_number = 14;
defparam ram_block3a14.port_b_last_address = 8191;
defparam ram_block3a14.port_b_logical_ram_depth = 16384;
defparam ram_block3a14.port_b_logical_ram_width = 32;
defparam ram_block3a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_read_enable_clock = "clock1";
defparam ram_block3a14.port_b_write_enable_clock = "clock1";
defparam ram_block3a14.ram_block_type = "M9K";
defparam ram_block3a14.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004007E01;
// synopsys translate_on

// Location: M9K_X51_Y26_N0
cycloneive_ram_block ram_block3a47(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a47_PORTADATAOUT_bus),
	.portbdataout(ram_block3a47_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a47.clk0_core_clock_enable = "ena0";
defparam ram_block3a47.clk1_core_clock_enable = "ena1";
defparam ram_block3a47.data_interleave_offset_in_bits = 1;
defparam ram_block3a47.data_interleave_width_in_bits = 1;
defparam ram_block3a47.init_file = "meminit.hex";
defparam ram_block3a47.init_file_layout = "port_a";
defparam ram_block3a47.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a47.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a47.operation_mode = "bidir_dual_port";
defparam ram_block3a47.port_a_address_clear = "none";
defparam ram_block3a47.port_a_address_width = 13;
defparam ram_block3a47.port_a_byte_enable_clock = "none";
defparam ram_block3a47.port_a_data_out_clear = "none";
defparam ram_block3a47.port_a_data_out_clock = "none";
defparam ram_block3a47.port_a_data_width = 1;
defparam ram_block3a47.port_a_first_address = 0;
defparam ram_block3a47.port_a_first_bit_number = 15;
defparam ram_block3a47.port_a_last_address = 8191;
defparam ram_block3a47.port_a_logical_ram_depth = 16384;
defparam ram_block3a47.port_a_logical_ram_width = 32;
defparam ram_block3a47.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_address_clear = "none";
defparam ram_block3a47.port_b_address_clock = "clock1";
defparam ram_block3a47.port_b_address_width = 13;
defparam ram_block3a47.port_b_data_in_clock = "clock1";
defparam ram_block3a47.port_b_data_out_clear = "none";
defparam ram_block3a47.port_b_data_out_clock = "none";
defparam ram_block3a47.port_b_data_width = 1;
defparam ram_block3a47.port_b_first_address = 0;
defparam ram_block3a47.port_b_first_bit_number = 15;
defparam ram_block3a47.port_b_last_address = 8191;
defparam ram_block3a47.port_b_logical_ram_depth = 16384;
defparam ram_block3a47.port_b_logical_ram_width = 32;
defparam ram_block3a47.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_read_enable_clock = "clock1";
defparam ram_block3a47.port_b_write_enable_clock = "clock1";
defparam ram_block3a47.ram_block_type = "M9K";
defparam ram_block3a47.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y26_N0
cycloneive_ram_block ram_block3a15(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a15_PORTADATAOUT_bus),
	.portbdataout(ram_block3a15_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a15.clk0_core_clock_enable = "ena0";
defparam ram_block3a15.clk1_core_clock_enable = "ena1";
defparam ram_block3a15.data_interleave_offset_in_bits = 1;
defparam ram_block3a15.data_interleave_width_in_bits = 1;
defparam ram_block3a15.init_file = "meminit.hex";
defparam ram_block3a15.init_file_layout = "port_a";
defparam ram_block3a15.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a15.operation_mode = "bidir_dual_port";
defparam ram_block3a15.port_a_address_clear = "none";
defparam ram_block3a15.port_a_address_width = 13;
defparam ram_block3a15.port_a_byte_enable_clock = "none";
defparam ram_block3a15.port_a_data_out_clear = "none";
defparam ram_block3a15.port_a_data_out_clock = "none";
defparam ram_block3a15.port_a_data_width = 1;
defparam ram_block3a15.port_a_first_address = 0;
defparam ram_block3a15.port_a_first_bit_number = 15;
defparam ram_block3a15.port_a_last_address = 8191;
defparam ram_block3a15.port_a_logical_ram_depth = 16384;
defparam ram_block3a15.port_a_logical_ram_width = 32;
defparam ram_block3a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_address_clear = "none";
defparam ram_block3a15.port_b_address_clock = "clock1";
defparam ram_block3a15.port_b_address_width = 13;
defparam ram_block3a15.port_b_data_in_clock = "clock1";
defparam ram_block3a15.port_b_data_out_clear = "none";
defparam ram_block3a15.port_b_data_out_clock = "none";
defparam ram_block3a15.port_b_data_width = 1;
defparam ram_block3a15.port_b_first_address = 0;
defparam ram_block3a15.port_b_first_bit_number = 15;
defparam ram_block3a15.port_b_last_address = 8191;
defparam ram_block3a15.port_b_logical_ram_depth = 16384;
defparam ram_block3a15.port_b_logical_ram_width = 32;
defparam ram_block3a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_read_enable_clock = "clock1";
defparam ram_block3a15.port_b_write_enable_clock = "clock1";
defparam ram_block3a15.ram_block_type = "M9K";
defparam ram_block3a15.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004000901;
// synopsys translate_on

// Location: M9K_X64_Y36_N0
cycloneive_ram_block ram_block3a48(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a48_PORTADATAOUT_bus),
	.portbdataout(ram_block3a48_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a48.clk0_core_clock_enable = "ena0";
defparam ram_block3a48.clk1_core_clock_enable = "ena1";
defparam ram_block3a48.data_interleave_offset_in_bits = 1;
defparam ram_block3a48.data_interleave_width_in_bits = 1;
defparam ram_block3a48.init_file = "meminit.hex";
defparam ram_block3a48.init_file_layout = "port_a";
defparam ram_block3a48.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a48.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a48.operation_mode = "bidir_dual_port";
defparam ram_block3a48.port_a_address_clear = "none";
defparam ram_block3a48.port_a_address_width = 13;
defparam ram_block3a48.port_a_byte_enable_clock = "none";
defparam ram_block3a48.port_a_data_out_clear = "none";
defparam ram_block3a48.port_a_data_out_clock = "none";
defparam ram_block3a48.port_a_data_width = 1;
defparam ram_block3a48.port_a_first_address = 0;
defparam ram_block3a48.port_a_first_bit_number = 16;
defparam ram_block3a48.port_a_last_address = 8191;
defparam ram_block3a48.port_a_logical_ram_depth = 16384;
defparam ram_block3a48.port_a_logical_ram_width = 32;
defparam ram_block3a48.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_address_clear = "none";
defparam ram_block3a48.port_b_address_clock = "clock1";
defparam ram_block3a48.port_b_address_width = 13;
defparam ram_block3a48.port_b_data_in_clock = "clock1";
defparam ram_block3a48.port_b_data_out_clear = "none";
defparam ram_block3a48.port_b_data_out_clock = "none";
defparam ram_block3a48.port_b_data_width = 1;
defparam ram_block3a48.port_b_first_address = 0;
defparam ram_block3a48.port_b_first_bit_number = 16;
defparam ram_block3a48.port_b_last_address = 8191;
defparam ram_block3a48.port_b_logical_ram_depth = 16384;
defparam ram_block3a48.port_b_logical_ram_width = 32;
defparam ram_block3a48.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_read_enable_clock = "clock1";
defparam ram_block3a48.port_b_write_enable_clock = "clock1";
defparam ram_block3a48.ram_block_type = "M9K";
defparam ram_block3a48.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y44_N0
cycloneive_ram_block ram_block3a16(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a16_PORTADATAOUT_bus),
	.portbdataout(ram_block3a16_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a16.clk0_core_clock_enable = "ena0";
defparam ram_block3a16.clk1_core_clock_enable = "ena1";
defparam ram_block3a16.data_interleave_offset_in_bits = 1;
defparam ram_block3a16.data_interleave_width_in_bits = 1;
defparam ram_block3a16.init_file = "meminit.hex";
defparam ram_block3a16.init_file_layout = "port_a";
defparam ram_block3a16.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a16.operation_mode = "bidir_dual_port";
defparam ram_block3a16.port_a_address_clear = "none";
defparam ram_block3a16.port_a_address_width = 13;
defparam ram_block3a16.port_a_byte_enable_clock = "none";
defparam ram_block3a16.port_a_data_out_clear = "none";
defparam ram_block3a16.port_a_data_out_clock = "none";
defparam ram_block3a16.port_a_data_width = 1;
defparam ram_block3a16.port_a_first_address = 0;
defparam ram_block3a16.port_a_first_bit_number = 16;
defparam ram_block3a16.port_a_last_address = 8191;
defparam ram_block3a16.port_a_logical_ram_depth = 16384;
defparam ram_block3a16.port_a_logical_ram_width = 32;
defparam ram_block3a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_address_clear = "none";
defparam ram_block3a16.port_b_address_clock = "clock1";
defparam ram_block3a16.port_b_address_width = 13;
defparam ram_block3a16.port_b_data_in_clock = "clock1";
defparam ram_block3a16.port_b_data_out_clear = "none";
defparam ram_block3a16.port_b_data_out_clock = "none";
defparam ram_block3a16.port_b_data_width = 1;
defparam ram_block3a16.port_b_first_address = 0;
defparam ram_block3a16.port_b_first_bit_number = 16;
defparam ram_block3a16.port_b_last_address = 8191;
defparam ram_block3a16.port_b_logical_ram_depth = 16384;
defparam ram_block3a16.port_b_logical_ram_width = 32;
defparam ram_block3a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_read_enable_clock = "clock1";
defparam ram_block3a16.port_b_write_enable_clock = "clock1";
defparam ram_block3a16.ram_block_type = "M9K";
defparam ram_block3a16.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005558145;
// synopsys translate_on

// Location: M9K_X51_Y36_N0
cycloneive_ram_block ram_block3a49(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a49_PORTADATAOUT_bus),
	.portbdataout(ram_block3a49_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a49.clk0_core_clock_enable = "ena0";
defparam ram_block3a49.clk1_core_clock_enable = "ena1";
defparam ram_block3a49.data_interleave_offset_in_bits = 1;
defparam ram_block3a49.data_interleave_width_in_bits = 1;
defparam ram_block3a49.init_file = "meminit.hex";
defparam ram_block3a49.init_file_layout = "port_a";
defparam ram_block3a49.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a49.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a49.operation_mode = "bidir_dual_port";
defparam ram_block3a49.port_a_address_clear = "none";
defparam ram_block3a49.port_a_address_width = 13;
defparam ram_block3a49.port_a_byte_enable_clock = "none";
defparam ram_block3a49.port_a_data_out_clear = "none";
defparam ram_block3a49.port_a_data_out_clock = "none";
defparam ram_block3a49.port_a_data_width = 1;
defparam ram_block3a49.port_a_first_address = 0;
defparam ram_block3a49.port_a_first_bit_number = 17;
defparam ram_block3a49.port_a_last_address = 8191;
defparam ram_block3a49.port_a_logical_ram_depth = 16384;
defparam ram_block3a49.port_a_logical_ram_width = 32;
defparam ram_block3a49.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_address_clear = "none";
defparam ram_block3a49.port_b_address_clock = "clock1";
defparam ram_block3a49.port_b_address_width = 13;
defparam ram_block3a49.port_b_data_in_clock = "clock1";
defparam ram_block3a49.port_b_data_out_clear = "none";
defparam ram_block3a49.port_b_data_out_clock = "none";
defparam ram_block3a49.port_b_data_width = 1;
defparam ram_block3a49.port_b_first_address = 0;
defparam ram_block3a49.port_b_first_bit_number = 17;
defparam ram_block3a49.port_b_last_address = 8191;
defparam ram_block3a49.port_b_logical_ram_depth = 16384;
defparam ram_block3a49.port_b_logical_ram_width = 32;
defparam ram_block3a49.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_read_enable_clock = "clock1";
defparam ram_block3a49.port_b_write_enable_clock = "clock1";
defparam ram_block3a49.ram_block_type = "M9K";
defparam ram_block3a49.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y38_N0
cycloneive_ram_block ram_block3a17(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a17_PORTADATAOUT_bus),
	.portbdataout(ram_block3a17_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a17.clk0_core_clock_enable = "ena0";
defparam ram_block3a17.clk1_core_clock_enable = "ena1";
defparam ram_block3a17.data_interleave_offset_in_bits = 1;
defparam ram_block3a17.data_interleave_width_in_bits = 1;
defparam ram_block3a17.init_file = "meminit.hex";
defparam ram_block3a17.init_file_layout = "port_a";
defparam ram_block3a17.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a17.operation_mode = "bidir_dual_port";
defparam ram_block3a17.port_a_address_clear = "none";
defparam ram_block3a17.port_a_address_width = 13;
defparam ram_block3a17.port_a_byte_enable_clock = "none";
defparam ram_block3a17.port_a_data_out_clear = "none";
defparam ram_block3a17.port_a_data_out_clock = "none";
defparam ram_block3a17.port_a_data_width = 1;
defparam ram_block3a17.port_a_first_address = 0;
defparam ram_block3a17.port_a_first_bit_number = 17;
defparam ram_block3a17.port_a_last_address = 8191;
defparam ram_block3a17.port_a_logical_ram_depth = 16384;
defparam ram_block3a17.port_a_logical_ram_width = 32;
defparam ram_block3a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_address_clear = "none";
defparam ram_block3a17.port_b_address_clock = "clock1";
defparam ram_block3a17.port_b_address_width = 13;
defparam ram_block3a17.port_b_data_in_clock = "clock1";
defparam ram_block3a17.port_b_data_out_clear = "none";
defparam ram_block3a17.port_b_data_out_clock = "none";
defparam ram_block3a17.port_b_data_width = 1;
defparam ram_block3a17.port_b_first_address = 0;
defparam ram_block3a17.port_b_first_bit_number = 17;
defparam ram_block3a17.port_b_last_address = 8191;
defparam ram_block3a17.port_b_logical_ram_depth = 16384;
defparam ram_block3a17.port_b_logical_ram_width = 32;
defparam ram_block3a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_read_enable_clock = "clock1";
defparam ram_block3a17.port_b_write_enable_clock = "clock1";
defparam ram_block3a17.ram_block_type = "M9K";
defparam ram_block3a17.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005994FBA;
// synopsys translate_on

// Location: M9K_X64_Y25_N0
cycloneive_ram_block ram_block3a50(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a50_PORTADATAOUT_bus),
	.portbdataout(ram_block3a50_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a50.clk0_core_clock_enable = "ena0";
defparam ram_block3a50.clk1_core_clock_enable = "ena1";
defparam ram_block3a50.data_interleave_offset_in_bits = 1;
defparam ram_block3a50.data_interleave_width_in_bits = 1;
defparam ram_block3a50.init_file = "meminit.hex";
defparam ram_block3a50.init_file_layout = "port_a";
defparam ram_block3a50.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a50.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a50.operation_mode = "bidir_dual_port";
defparam ram_block3a50.port_a_address_clear = "none";
defparam ram_block3a50.port_a_address_width = 13;
defparam ram_block3a50.port_a_byte_enable_clock = "none";
defparam ram_block3a50.port_a_data_out_clear = "none";
defparam ram_block3a50.port_a_data_out_clock = "none";
defparam ram_block3a50.port_a_data_width = 1;
defparam ram_block3a50.port_a_first_address = 0;
defparam ram_block3a50.port_a_first_bit_number = 18;
defparam ram_block3a50.port_a_last_address = 8191;
defparam ram_block3a50.port_a_logical_ram_depth = 16384;
defparam ram_block3a50.port_a_logical_ram_width = 32;
defparam ram_block3a50.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_address_clear = "none";
defparam ram_block3a50.port_b_address_clock = "clock1";
defparam ram_block3a50.port_b_address_width = 13;
defparam ram_block3a50.port_b_data_in_clock = "clock1";
defparam ram_block3a50.port_b_data_out_clear = "none";
defparam ram_block3a50.port_b_data_out_clock = "none";
defparam ram_block3a50.port_b_data_width = 1;
defparam ram_block3a50.port_b_first_address = 0;
defparam ram_block3a50.port_b_first_bit_number = 18;
defparam ram_block3a50.port_b_last_address = 8191;
defparam ram_block3a50.port_b_logical_ram_depth = 16384;
defparam ram_block3a50.port_b_logical_ram_width = 32;
defparam ram_block3a50.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_read_enable_clock = "clock1";
defparam ram_block3a50.port_b_write_enable_clock = "clock1";
defparam ram_block3a50.ram_block_type = "M9K";
defparam ram_block3a50.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y28_N0
cycloneive_ram_block ram_block3a18(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a18_PORTADATAOUT_bus),
	.portbdataout(ram_block3a18_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a18.clk0_core_clock_enable = "ena0";
defparam ram_block3a18.clk1_core_clock_enable = "ena1";
defparam ram_block3a18.data_interleave_offset_in_bits = 1;
defparam ram_block3a18.data_interleave_width_in_bits = 1;
defparam ram_block3a18.init_file = "meminit.hex";
defparam ram_block3a18.init_file_layout = "port_a";
defparam ram_block3a18.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a18.operation_mode = "bidir_dual_port";
defparam ram_block3a18.port_a_address_clear = "none";
defparam ram_block3a18.port_a_address_width = 13;
defparam ram_block3a18.port_a_byte_enable_clock = "none";
defparam ram_block3a18.port_a_data_out_clear = "none";
defparam ram_block3a18.port_a_data_out_clock = "none";
defparam ram_block3a18.port_a_data_width = 1;
defparam ram_block3a18.port_a_first_address = 0;
defparam ram_block3a18.port_a_first_bit_number = 18;
defparam ram_block3a18.port_a_last_address = 8191;
defparam ram_block3a18.port_a_logical_ram_depth = 16384;
defparam ram_block3a18.port_a_logical_ram_width = 32;
defparam ram_block3a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_address_clear = "none";
defparam ram_block3a18.port_b_address_clock = "clock1";
defparam ram_block3a18.port_b_address_width = 13;
defparam ram_block3a18.port_b_data_in_clock = "clock1";
defparam ram_block3a18.port_b_data_out_clear = "none";
defparam ram_block3a18.port_b_data_out_clock = "none";
defparam ram_block3a18.port_b_data_width = 1;
defparam ram_block3a18.port_b_first_address = 0;
defparam ram_block3a18.port_b_first_bit_number = 18;
defparam ram_block3a18.port_b_last_address = 8191;
defparam ram_block3a18.port_b_logical_ram_depth = 16384;
defparam ram_block3a18.port_b_logical_ram_width = 32;
defparam ram_block3a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_read_enable_clock = "clock1";
defparam ram_block3a18.port_b_write_enable_clock = "clock1";
defparam ram_block3a18.ram_block_type = "M9K";
defparam ram_block3a18.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000061E814C;
// synopsys translate_on

// Location: M9K_X64_Y29_N0
cycloneive_ram_block ram_block3a51(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a51_PORTADATAOUT_bus),
	.portbdataout(ram_block3a51_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a51.clk0_core_clock_enable = "ena0";
defparam ram_block3a51.clk1_core_clock_enable = "ena1";
defparam ram_block3a51.data_interleave_offset_in_bits = 1;
defparam ram_block3a51.data_interleave_width_in_bits = 1;
defparam ram_block3a51.init_file = "meminit.hex";
defparam ram_block3a51.init_file_layout = "port_a";
defparam ram_block3a51.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a51.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a51.operation_mode = "bidir_dual_port";
defparam ram_block3a51.port_a_address_clear = "none";
defparam ram_block3a51.port_a_address_width = 13;
defparam ram_block3a51.port_a_byte_enable_clock = "none";
defparam ram_block3a51.port_a_data_out_clear = "none";
defparam ram_block3a51.port_a_data_out_clock = "none";
defparam ram_block3a51.port_a_data_width = 1;
defparam ram_block3a51.port_a_first_address = 0;
defparam ram_block3a51.port_a_first_bit_number = 19;
defparam ram_block3a51.port_a_last_address = 8191;
defparam ram_block3a51.port_a_logical_ram_depth = 16384;
defparam ram_block3a51.port_a_logical_ram_width = 32;
defparam ram_block3a51.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_address_clear = "none";
defparam ram_block3a51.port_b_address_clock = "clock1";
defparam ram_block3a51.port_b_address_width = 13;
defparam ram_block3a51.port_b_data_in_clock = "clock1";
defparam ram_block3a51.port_b_data_out_clear = "none";
defparam ram_block3a51.port_b_data_out_clock = "none";
defparam ram_block3a51.port_b_data_width = 1;
defparam ram_block3a51.port_b_first_address = 0;
defparam ram_block3a51.port_b_first_bit_number = 19;
defparam ram_block3a51.port_b_last_address = 8191;
defparam ram_block3a51.port_b_logical_ram_depth = 16384;
defparam ram_block3a51.port_b_logical_ram_width = 32;
defparam ram_block3a51.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_read_enable_clock = "clock1";
defparam ram_block3a51.port_b_write_enable_clock = "clock1";
defparam ram_block3a51.ram_block_type = "M9K";
defparam ram_block3a51.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y21_N0
cycloneive_ram_block ram_block3a19(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a19_PORTADATAOUT_bus),
	.portbdataout(ram_block3a19_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a19.clk0_core_clock_enable = "ena0";
defparam ram_block3a19.clk1_core_clock_enable = "ena1";
defparam ram_block3a19.data_interleave_offset_in_bits = 1;
defparam ram_block3a19.data_interleave_width_in_bits = 1;
defparam ram_block3a19.init_file = "meminit.hex";
defparam ram_block3a19.init_file_layout = "port_a";
defparam ram_block3a19.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a19.operation_mode = "bidir_dual_port";
defparam ram_block3a19.port_a_address_clear = "none";
defparam ram_block3a19.port_a_address_width = 13;
defparam ram_block3a19.port_a_byte_enable_clock = "none";
defparam ram_block3a19.port_a_data_out_clear = "none";
defparam ram_block3a19.port_a_data_out_clock = "none";
defparam ram_block3a19.port_a_data_width = 1;
defparam ram_block3a19.port_a_first_address = 0;
defparam ram_block3a19.port_a_first_bit_number = 19;
defparam ram_block3a19.port_a_last_address = 8191;
defparam ram_block3a19.port_a_logical_ram_depth = 16384;
defparam ram_block3a19.port_a_logical_ram_width = 32;
defparam ram_block3a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_address_clear = "none";
defparam ram_block3a19.port_b_address_clock = "clock1";
defparam ram_block3a19.port_b_address_width = 13;
defparam ram_block3a19.port_b_data_in_clock = "clock1";
defparam ram_block3a19.port_b_data_out_clear = "none";
defparam ram_block3a19.port_b_data_out_clock = "none";
defparam ram_block3a19.port_b_data_width = 1;
defparam ram_block3a19.port_b_first_address = 0;
defparam ram_block3a19.port_b_first_bit_number = 19;
defparam ram_block3a19.port_b_last_address = 8191;
defparam ram_block3a19.port_b_logical_ram_depth = 16384;
defparam ram_block3a19.port_b_logical_ram_width = 32;
defparam ram_block3a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_read_enable_clock = "clock1";
defparam ram_block3a19.port_b_write_enable_clock = "clock1";
defparam ram_block3a19.ram_block_type = "M9K";
defparam ram_block3a19.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007E08800;
// synopsys translate_on

// Location: M9K_X51_Y40_N0
cycloneive_ram_block ram_block3a52(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a52_PORTADATAOUT_bus),
	.portbdataout(ram_block3a52_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a52.clk0_core_clock_enable = "ena0";
defparam ram_block3a52.clk1_core_clock_enable = "ena1";
defparam ram_block3a52.data_interleave_offset_in_bits = 1;
defparam ram_block3a52.data_interleave_width_in_bits = 1;
defparam ram_block3a52.init_file = "meminit.hex";
defparam ram_block3a52.init_file_layout = "port_a";
defparam ram_block3a52.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a52.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a52.operation_mode = "bidir_dual_port";
defparam ram_block3a52.port_a_address_clear = "none";
defparam ram_block3a52.port_a_address_width = 13;
defparam ram_block3a52.port_a_byte_enable_clock = "none";
defparam ram_block3a52.port_a_data_out_clear = "none";
defparam ram_block3a52.port_a_data_out_clock = "none";
defparam ram_block3a52.port_a_data_width = 1;
defparam ram_block3a52.port_a_first_address = 0;
defparam ram_block3a52.port_a_first_bit_number = 20;
defparam ram_block3a52.port_a_last_address = 8191;
defparam ram_block3a52.port_a_logical_ram_depth = 16384;
defparam ram_block3a52.port_a_logical_ram_width = 32;
defparam ram_block3a52.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_address_clear = "none";
defparam ram_block3a52.port_b_address_clock = "clock1";
defparam ram_block3a52.port_b_address_width = 13;
defparam ram_block3a52.port_b_data_in_clock = "clock1";
defparam ram_block3a52.port_b_data_out_clear = "none";
defparam ram_block3a52.port_b_data_out_clock = "none";
defparam ram_block3a52.port_b_data_width = 1;
defparam ram_block3a52.port_b_first_address = 0;
defparam ram_block3a52.port_b_first_bit_number = 20;
defparam ram_block3a52.port_b_last_address = 8191;
defparam ram_block3a52.port_b_logical_ram_depth = 16384;
defparam ram_block3a52.port_b_logical_ram_width = 32;
defparam ram_block3a52.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_read_enable_clock = "clock1";
defparam ram_block3a52.port_b_write_enable_clock = "clock1";
defparam ram_block3a52.ram_block_type = "M9K";
defparam ram_block3a52.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y39_N0
cycloneive_ram_block ram_block3a20(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a20_PORTADATAOUT_bus),
	.portbdataout(ram_block3a20_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a20.clk0_core_clock_enable = "ena0";
defparam ram_block3a20.clk1_core_clock_enable = "ena1";
defparam ram_block3a20.data_interleave_offset_in_bits = 1;
defparam ram_block3a20.data_interleave_width_in_bits = 1;
defparam ram_block3a20.init_file = "meminit.hex";
defparam ram_block3a20.init_file_layout = "port_a";
defparam ram_block3a20.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a20.operation_mode = "bidir_dual_port";
defparam ram_block3a20.port_a_address_clear = "none";
defparam ram_block3a20.port_a_address_width = 13;
defparam ram_block3a20.port_a_byte_enable_clock = "none";
defparam ram_block3a20.port_a_data_out_clear = "none";
defparam ram_block3a20.port_a_data_out_clock = "none";
defparam ram_block3a20.port_a_data_width = 1;
defparam ram_block3a20.port_a_first_address = 0;
defparam ram_block3a20.port_a_first_bit_number = 20;
defparam ram_block3a20.port_a_last_address = 8191;
defparam ram_block3a20.port_a_logical_ram_depth = 16384;
defparam ram_block3a20.port_a_logical_ram_width = 32;
defparam ram_block3a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_address_clear = "none";
defparam ram_block3a20.port_b_address_clock = "clock1";
defparam ram_block3a20.port_b_address_width = 13;
defparam ram_block3a20.port_b_data_in_clock = "clock1";
defparam ram_block3a20.port_b_data_out_clear = "none";
defparam ram_block3a20.port_b_data_out_clock = "none";
defparam ram_block3a20.port_b_data_width = 1;
defparam ram_block3a20.port_b_first_address = 0;
defparam ram_block3a20.port_b_first_bit_number = 20;
defparam ram_block3a20.port_b_last_address = 8191;
defparam ram_block3a20.port_b_logical_ram_depth = 16384;
defparam ram_block3a20.port_b_logical_ram_width = 32;
defparam ram_block3a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_read_enable_clock = "clock1";
defparam ram_block3a20.port_b_write_enable_clock = "clock1";
defparam ram_block3a20.ram_block_type = "M9K";
defparam ram_block3a20.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000400000C;
// synopsys translate_on

// Location: M9K_X51_Y42_N0
cycloneive_ram_block ram_block3a53(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a53_PORTADATAOUT_bus),
	.portbdataout(ram_block3a53_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a53.clk0_core_clock_enable = "ena0";
defparam ram_block3a53.clk1_core_clock_enable = "ena1";
defparam ram_block3a53.data_interleave_offset_in_bits = 1;
defparam ram_block3a53.data_interleave_width_in_bits = 1;
defparam ram_block3a53.init_file = "meminit.hex";
defparam ram_block3a53.init_file_layout = "port_a";
defparam ram_block3a53.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a53.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a53.operation_mode = "bidir_dual_port";
defparam ram_block3a53.port_a_address_clear = "none";
defparam ram_block3a53.port_a_address_width = 13;
defparam ram_block3a53.port_a_byte_enable_clock = "none";
defparam ram_block3a53.port_a_data_out_clear = "none";
defparam ram_block3a53.port_a_data_out_clock = "none";
defparam ram_block3a53.port_a_data_width = 1;
defparam ram_block3a53.port_a_first_address = 0;
defparam ram_block3a53.port_a_first_bit_number = 21;
defparam ram_block3a53.port_a_last_address = 8191;
defparam ram_block3a53.port_a_logical_ram_depth = 16384;
defparam ram_block3a53.port_a_logical_ram_width = 32;
defparam ram_block3a53.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_address_clear = "none";
defparam ram_block3a53.port_b_address_clock = "clock1";
defparam ram_block3a53.port_b_address_width = 13;
defparam ram_block3a53.port_b_data_in_clock = "clock1";
defparam ram_block3a53.port_b_data_out_clear = "none";
defparam ram_block3a53.port_b_data_out_clock = "none";
defparam ram_block3a53.port_b_data_width = 1;
defparam ram_block3a53.port_b_first_address = 0;
defparam ram_block3a53.port_b_first_bit_number = 21;
defparam ram_block3a53.port_b_last_address = 8191;
defparam ram_block3a53.port_b_logical_ram_depth = 16384;
defparam ram_block3a53.port_b_logical_ram_width = 32;
defparam ram_block3a53.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_read_enable_clock = "clock1";
defparam ram_block3a53.port_b_write_enable_clock = "clock1";
defparam ram_block3a53.ram_block_type = "M9K";
defparam ram_block3a53.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y22_N0
cycloneive_ram_block ram_block3a21(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a21_PORTADATAOUT_bus),
	.portbdataout(ram_block3a21_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a21.clk0_core_clock_enable = "ena0";
defparam ram_block3a21.clk1_core_clock_enable = "ena1";
defparam ram_block3a21.data_interleave_offset_in_bits = 1;
defparam ram_block3a21.data_interleave_width_in_bits = 1;
defparam ram_block3a21.init_file = "meminit.hex";
defparam ram_block3a21.init_file_layout = "port_a";
defparam ram_block3a21.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a21.operation_mode = "bidir_dual_port";
defparam ram_block3a21.port_a_address_clear = "none";
defparam ram_block3a21.port_a_address_width = 13;
defparam ram_block3a21.port_a_byte_enable_clock = "none";
defparam ram_block3a21.port_a_data_out_clear = "none";
defparam ram_block3a21.port_a_data_out_clock = "none";
defparam ram_block3a21.port_a_data_width = 1;
defparam ram_block3a21.port_a_first_address = 0;
defparam ram_block3a21.port_a_first_bit_number = 21;
defparam ram_block3a21.port_a_last_address = 8191;
defparam ram_block3a21.port_a_logical_ram_depth = 16384;
defparam ram_block3a21.port_a_logical_ram_width = 32;
defparam ram_block3a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_address_clear = "none";
defparam ram_block3a21.port_b_address_clock = "clock1";
defparam ram_block3a21.port_b_address_width = 13;
defparam ram_block3a21.port_b_data_in_clock = "clock1";
defparam ram_block3a21.port_b_data_out_clear = "none";
defparam ram_block3a21.port_b_data_out_clock = "none";
defparam ram_block3a21.port_b_data_width = 1;
defparam ram_block3a21.port_b_first_address = 0;
defparam ram_block3a21.port_b_first_bit_number = 21;
defparam ram_block3a21.port_b_last_address = 8191;
defparam ram_block3a21.port_b_logical_ram_depth = 16384;
defparam ram_block3a21.port_b_logical_ram_width = 32;
defparam ram_block3a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_read_enable_clock = "clock1";
defparam ram_block3a21.port_b_write_enable_clock = "clock1";
defparam ram_block3a21.ram_block_type = "M9K";
defparam ram_block3a21.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FF7DF0;
// synopsys translate_on

// Location: M9K_X64_Y40_N0
cycloneive_ram_block ram_block3a54(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a54_PORTADATAOUT_bus),
	.portbdataout(ram_block3a54_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a54.clk0_core_clock_enable = "ena0";
defparam ram_block3a54.clk1_core_clock_enable = "ena1";
defparam ram_block3a54.data_interleave_offset_in_bits = 1;
defparam ram_block3a54.data_interleave_width_in_bits = 1;
defparam ram_block3a54.init_file = "meminit.hex";
defparam ram_block3a54.init_file_layout = "port_a";
defparam ram_block3a54.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a54.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a54.operation_mode = "bidir_dual_port";
defparam ram_block3a54.port_a_address_clear = "none";
defparam ram_block3a54.port_a_address_width = 13;
defparam ram_block3a54.port_a_byte_enable_clock = "none";
defparam ram_block3a54.port_a_data_out_clear = "none";
defparam ram_block3a54.port_a_data_out_clock = "none";
defparam ram_block3a54.port_a_data_width = 1;
defparam ram_block3a54.port_a_first_address = 0;
defparam ram_block3a54.port_a_first_bit_number = 22;
defparam ram_block3a54.port_a_last_address = 8191;
defparam ram_block3a54.port_a_logical_ram_depth = 16384;
defparam ram_block3a54.port_a_logical_ram_width = 32;
defparam ram_block3a54.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_address_clear = "none";
defparam ram_block3a54.port_b_address_clock = "clock1";
defparam ram_block3a54.port_b_address_width = 13;
defparam ram_block3a54.port_b_data_in_clock = "clock1";
defparam ram_block3a54.port_b_data_out_clear = "none";
defparam ram_block3a54.port_b_data_out_clock = "none";
defparam ram_block3a54.port_b_data_width = 1;
defparam ram_block3a54.port_b_first_address = 0;
defparam ram_block3a54.port_b_first_bit_number = 22;
defparam ram_block3a54.port_b_last_address = 8191;
defparam ram_block3a54.port_b_logical_ram_depth = 16384;
defparam ram_block3a54.port_b_logical_ram_width = 32;
defparam ram_block3a54.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_read_enable_clock = "clock1";
defparam ram_block3a54.port_b_write_enable_clock = "clock1";
defparam ram_block3a54.ram_block_type = "M9K";
defparam ram_block3a54.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y42_N0
cycloneive_ram_block ram_block3a22(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a22_PORTADATAOUT_bus),
	.portbdataout(ram_block3a22_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a22.clk0_core_clock_enable = "ena0";
defparam ram_block3a22.clk1_core_clock_enable = "ena1";
defparam ram_block3a22.data_interleave_offset_in_bits = 1;
defparam ram_block3a22.data_interleave_width_in_bits = 1;
defparam ram_block3a22.init_file = "meminit.hex";
defparam ram_block3a22.init_file_layout = "port_a";
defparam ram_block3a22.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a22.operation_mode = "bidir_dual_port";
defparam ram_block3a22.port_a_address_clear = "none";
defparam ram_block3a22.port_a_address_width = 13;
defparam ram_block3a22.port_a_byte_enable_clock = "none";
defparam ram_block3a22.port_a_data_out_clear = "none";
defparam ram_block3a22.port_a_data_out_clock = "none";
defparam ram_block3a22.port_a_data_width = 1;
defparam ram_block3a22.port_a_first_address = 0;
defparam ram_block3a22.port_a_first_bit_number = 22;
defparam ram_block3a22.port_a_last_address = 8191;
defparam ram_block3a22.port_a_logical_ram_depth = 16384;
defparam ram_block3a22.port_a_logical_ram_width = 32;
defparam ram_block3a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_address_clear = "none";
defparam ram_block3a22.port_b_address_clock = "clock1";
defparam ram_block3a22.port_b_address_width = 13;
defparam ram_block3a22.port_b_data_in_clock = "clock1";
defparam ram_block3a22.port_b_data_out_clear = "none";
defparam ram_block3a22.port_b_data_out_clock = "none";
defparam ram_block3a22.port_b_data_width = 1;
defparam ram_block3a22.port_b_first_address = 0;
defparam ram_block3a22.port_b_first_bit_number = 22;
defparam ram_block3a22.port_b_last_address = 8191;
defparam ram_block3a22.port_b_logical_ram_depth = 16384;
defparam ram_block3a22.port_b_logical_ram_width = 32;
defparam ram_block3a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_read_enable_clock = "clock1";
defparam ram_block3a22.port_b_write_enable_clock = "clock1";
defparam ram_block3a22.ram_block_type = "M9K";
defparam ram_block3a22.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004008100;
// synopsys translate_on

// Location: M9K_X51_Y25_N0
cycloneive_ram_block ram_block3a55(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a55_PORTADATAOUT_bus),
	.portbdataout(ram_block3a55_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a55.clk0_core_clock_enable = "ena0";
defparam ram_block3a55.clk1_core_clock_enable = "ena1";
defparam ram_block3a55.data_interleave_offset_in_bits = 1;
defparam ram_block3a55.data_interleave_width_in_bits = 1;
defparam ram_block3a55.init_file = "meminit.hex";
defparam ram_block3a55.init_file_layout = "port_a";
defparam ram_block3a55.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a55.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a55.operation_mode = "bidir_dual_port";
defparam ram_block3a55.port_a_address_clear = "none";
defparam ram_block3a55.port_a_address_width = 13;
defparam ram_block3a55.port_a_byte_enable_clock = "none";
defparam ram_block3a55.port_a_data_out_clear = "none";
defparam ram_block3a55.port_a_data_out_clock = "none";
defparam ram_block3a55.port_a_data_width = 1;
defparam ram_block3a55.port_a_first_address = 0;
defparam ram_block3a55.port_a_first_bit_number = 23;
defparam ram_block3a55.port_a_last_address = 8191;
defparam ram_block3a55.port_a_logical_ram_depth = 16384;
defparam ram_block3a55.port_a_logical_ram_width = 32;
defparam ram_block3a55.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_address_clear = "none";
defparam ram_block3a55.port_b_address_clock = "clock1";
defparam ram_block3a55.port_b_address_width = 13;
defparam ram_block3a55.port_b_data_in_clock = "clock1";
defparam ram_block3a55.port_b_data_out_clear = "none";
defparam ram_block3a55.port_b_data_out_clock = "none";
defparam ram_block3a55.port_b_data_width = 1;
defparam ram_block3a55.port_b_first_address = 0;
defparam ram_block3a55.port_b_first_bit_number = 23;
defparam ram_block3a55.port_b_last_address = 8191;
defparam ram_block3a55.port_b_logical_ram_depth = 16384;
defparam ram_block3a55.port_b_logical_ram_width = 32;
defparam ram_block3a55.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_read_enable_clock = "clock1";
defparam ram_block3a55.port_b_write_enable_clock = "clock1";
defparam ram_block3a55.ram_block_type = "M9K";
defparam ram_block3a55.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y36_N0
cycloneive_ram_block ram_block3a23(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a23_PORTADATAOUT_bus),
	.portbdataout(ram_block3a23_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a23.clk0_core_clock_enable = "ena0";
defparam ram_block3a23.clk1_core_clock_enable = "ena1";
defparam ram_block3a23.data_interleave_offset_in_bits = 1;
defparam ram_block3a23.data_interleave_width_in_bits = 1;
defparam ram_block3a23.init_file = "meminit.hex";
defparam ram_block3a23.init_file_layout = "port_a";
defparam ram_block3a23.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a23.operation_mode = "bidir_dual_port";
defparam ram_block3a23.port_a_address_clear = "none";
defparam ram_block3a23.port_a_address_width = 13;
defparam ram_block3a23.port_a_byte_enable_clock = "none";
defparam ram_block3a23.port_a_data_out_clear = "none";
defparam ram_block3a23.port_a_data_out_clock = "none";
defparam ram_block3a23.port_a_data_width = 1;
defparam ram_block3a23.port_a_first_address = 0;
defparam ram_block3a23.port_a_first_bit_number = 23;
defparam ram_block3a23.port_a_last_address = 8191;
defparam ram_block3a23.port_a_logical_ram_depth = 16384;
defparam ram_block3a23.port_a_logical_ram_width = 32;
defparam ram_block3a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_address_clear = "none";
defparam ram_block3a23.port_b_address_clock = "clock1";
defparam ram_block3a23.port_b_address_width = 13;
defparam ram_block3a23.port_b_data_in_clock = "clock1";
defparam ram_block3a23.port_b_data_out_clear = "none";
defparam ram_block3a23.port_b_data_out_clock = "none";
defparam ram_block3a23.port_b_data_width = 1;
defparam ram_block3a23.port_b_first_address = 0;
defparam ram_block3a23.port_b_first_bit_number = 23;
defparam ram_block3a23.port_b_last_address = 8191;
defparam ram_block3a23.port_b_logical_ram_depth = 16384;
defparam ram_block3a23.port_b_logical_ram_width = 32;
defparam ram_block3a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_read_enable_clock = "clock1";
defparam ram_block3a23.port_b_write_enable_clock = "clock1";
defparam ram_block3a23.ram_block_type = "M9K";
defparam ram_block3a23.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FF8600;
// synopsys translate_on

// Location: M9K_X78_Y34_N0
cycloneive_ram_block ram_block3a56(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a56_PORTADATAOUT_bus),
	.portbdataout(ram_block3a56_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a56.clk0_core_clock_enable = "ena0";
defparam ram_block3a56.clk1_core_clock_enable = "ena1";
defparam ram_block3a56.data_interleave_offset_in_bits = 1;
defparam ram_block3a56.data_interleave_width_in_bits = 1;
defparam ram_block3a56.init_file = "meminit.hex";
defparam ram_block3a56.init_file_layout = "port_a";
defparam ram_block3a56.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a56.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a56.operation_mode = "bidir_dual_port";
defparam ram_block3a56.port_a_address_clear = "none";
defparam ram_block3a56.port_a_address_width = 13;
defparam ram_block3a56.port_a_byte_enable_clock = "none";
defparam ram_block3a56.port_a_data_out_clear = "none";
defparam ram_block3a56.port_a_data_out_clock = "none";
defparam ram_block3a56.port_a_data_width = 1;
defparam ram_block3a56.port_a_first_address = 0;
defparam ram_block3a56.port_a_first_bit_number = 24;
defparam ram_block3a56.port_a_last_address = 8191;
defparam ram_block3a56.port_a_logical_ram_depth = 16384;
defparam ram_block3a56.port_a_logical_ram_width = 32;
defparam ram_block3a56.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_address_clear = "none";
defparam ram_block3a56.port_b_address_clock = "clock1";
defparam ram_block3a56.port_b_address_width = 13;
defparam ram_block3a56.port_b_data_in_clock = "clock1";
defparam ram_block3a56.port_b_data_out_clear = "none";
defparam ram_block3a56.port_b_data_out_clock = "none";
defparam ram_block3a56.port_b_data_width = 1;
defparam ram_block3a56.port_b_first_address = 0;
defparam ram_block3a56.port_b_first_bit_number = 24;
defparam ram_block3a56.port_b_last_address = 8191;
defparam ram_block3a56.port_b_logical_ram_depth = 16384;
defparam ram_block3a56.port_b_logical_ram_width = 32;
defparam ram_block3a56.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_read_enable_clock = "clock1";
defparam ram_block3a56.port_b_write_enable_clock = "clock1";
defparam ram_block3a56.ram_block_type = "M9K";
defparam ram_block3a56.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y34_N0
cycloneive_ram_block ram_block3a24(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a24_PORTADATAOUT_bus),
	.portbdataout(ram_block3a24_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a24.clk0_core_clock_enable = "ena0";
defparam ram_block3a24.clk1_core_clock_enable = "ena1";
defparam ram_block3a24.data_interleave_offset_in_bits = 1;
defparam ram_block3a24.data_interleave_width_in_bits = 1;
defparam ram_block3a24.init_file = "meminit.hex";
defparam ram_block3a24.init_file_layout = "port_a";
defparam ram_block3a24.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a24.operation_mode = "bidir_dual_port";
defparam ram_block3a24.port_a_address_clear = "none";
defparam ram_block3a24.port_a_address_width = 13;
defparam ram_block3a24.port_a_byte_enable_clock = "none";
defparam ram_block3a24.port_a_data_out_clear = "none";
defparam ram_block3a24.port_a_data_out_clock = "none";
defparam ram_block3a24.port_a_data_width = 1;
defparam ram_block3a24.port_a_first_address = 0;
defparam ram_block3a24.port_a_first_bit_number = 24;
defparam ram_block3a24.port_a_last_address = 8191;
defparam ram_block3a24.port_a_logical_ram_depth = 16384;
defparam ram_block3a24.port_a_logical_ram_width = 32;
defparam ram_block3a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_address_clear = "none";
defparam ram_block3a24.port_b_address_clock = "clock1";
defparam ram_block3a24.port_b_address_width = 13;
defparam ram_block3a24.port_b_data_in_clock = "clock1";
defparam ram_block3a24.port_b_data_out_clear = "none";
defparam ram_block3a24.port_b_data_out_clock = "none";
defparam ram_block3a24.port_b_data_width = 1;
defparam ram_block3a24.port_b_first_address = 0;
defparam ram_block3a24.port_b_first_bit_number = 24;
defparam ram_block3a24.port_b_last_address = 8191;
defparam ram_block3a24.port_b_logical_ram_depth = 16384;
defparam ram_block3a24.port_b_logical_ram_width = 32;
defparam ram_block3a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_read_enable_clock = "clock1";
defparam ram_block3a24.port_b_write_enable_clock = "clock1";
defparam ram_block3a24.ram_block_type = "M9K";
defparam ram_block3a24.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004000000;
// synopsys translate_on

// Location: M9K_X78_Y31_N0
cycloneive_ram_block ram_block3a57(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a57_PORTADATAOUT_bus),
	.portbdataout(ram_block3a57_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a57.clk0_core_clock_enable = "ena0";
defparam ram_block3a57.clk1_core_clock_enable = "ena1";
defparam ram_block3a57.data_interleave_offset_in_bits = 1;
defparam ram_block3a57.data_interleave_width_in_bits = 1;
defparam ram_block3a57.init_file = "meminit.hex";
defparam ram_block3a57.init_file_layout = "port_a";
defparam ram_block3a57.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a57.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a57.operation_mode = "bidir_dual_port";
defparam ram_block3a57.port_a_address_clear = "none";
defparam ram_block3a57.port_a_address_width = 13;
defparam ram_block3a57.port_a_byte_enable_clock = "none";
defparam ram_block3a57.port_a_data_out_clear = "none";
defparam ram_block3a57.port_a_data_out_clock = "none";
defparam ram_block3a57.port_a_data_width = 1;
defparam ram_block3a57.port_a_first_address = 0;
defparam ram_block3a57.port_a_first_bit_number = 25;
defparam ram_block3a57.port_a_last_address = 8191;
defparam ram_block3a57.port_a_logical_ram_depth = 16384;
defparam ram_block3a57.port_a_logical_ram_width = 32;
defparam ram_block3a57.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_address_clear = "none";
defparam ram_block3a57.port_b_address_clock = "clock1";
defparam ram_block3a57.port_b_address_width = 13;
defparam ram_block3a57.port_b_data_in_clock = "clock1";
defparam ram_block3a57.port_b_data_out_clear = "none";
defparam ram_block3a57.port_b_data_out_clock = "none";
defparam ram_block3a57.port_b_data_width = 1;
defparam ram_block3a57.port_b_first_address = 0;
defparam ram_block3a57.port_b_first_bit_number = 25;
defparam ram_block3a57.port_b_last_address = 8191;
defparam ram_block3a57.port_b_logical_ram_depth = 16384;
defparam ram_block3a57.port_b_logical_ram_width = 32;
defparam ram_block3a57.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_read_enable_clock = "clock1";
defparam ram_block3a57.port_b_write_enable_clock = "clock1";
defparam ram_block3a57.ram_block_type = "M9K";
defparam ram_block3a57.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y30_N0
cycloneive_ram_block ram_block3a25(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a25_PORTADATAOUT_bus),
	.portbdataout(ram_block3a25_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a25.clk0_core_clock_enable = "ena0";
defparam ram_block3a25.clk1_core_clock_enable = "ena1";
defparam ram_block3a25.data_interleave_offset_in_bits = 1;
defparam ram_block3a25.data_interleave_width_in_bits = 1;
defparam ram_block3a25.init_file = "meminit.hex";
defparam ram_block3a25.init_file_layout = "port_a";
defparam ram_block3a25.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a25.operation_mode = "bidir_dual_port";
defparam ram_block3a25.port_a_address_clear = "none";
defparam ram_block3a25.port_a_address_width = 13;
defparam ram_block3a25.port_a_byte_enable_clock = "none";
defparam ram_block3a25.port_a_data_out_clear = "none";
defparam ram_block3a25.port_a_data_out_clock = "none";
defparam ram_block3a25.port_a_data_width = 1;
defparam ram_block3a25.port_a_first_address = 0;
defparam ram_block3a25.port_a_first_bit_number = 25;
defparam ram_block3a25.port_a_last_address = 8191;
defparam ram_block3a25.port_a_logical_ram_depth = 16384;
defparam ram_block3a25.port_a_logical_ram_width = 32;
defparam ram_block3a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_address_clear = "none";
defparam ram_block3a25.port_b_address_clock = "clock1";
defparam ram_block3a25.port_b_address_width = 13;
defparam ram_block3a25.port_b_data_in_clock = "clock1";
defparam ram_block3a25.port_b_data_out_clear = "none";
defparam ram_block3a25.port_b_data_out_clock = "none";
defparam ram_block3a25.port_b_data_width = 1;
defparam ram_block3a25.port_b_first_address = 0;
defparam ram_block3a25.port_b_first_bit_number = 25;
defparam ram_block3a25.port_b_last_address = 8191;
defparam ram_block3a25.port_b_logical_ram_depth = 16384;
defparam ram_block3a25.port_b_logical_ram_width = 32;
defparam ram_block3a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_read_enable_clock = "clock1";
defparam ram_block3a25.port_b_write_enable_clock = "clock1";
defparam ram_block3a25.ram_block_type = "M9K";
defparam ram_block3a25.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FF8000;
// synopsys translate_on

// Location: M9K_X37_Y34_N0
cycloneive_ram_block ram_block3a58(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a58_PORTADATAOUT_bus),
	.portbdataout(ram_block3a58_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a58.clk0_core_clock_enable = "ena0";
defparam ram_block3a58.clk1_core_clock_enable = "ena1";
defparam ram_block3a58.data_interleave_offset_in_bits = 1;
defparam ram_block3a58.data_interleave_width_in_bits = 1;
defparam ram_block3a58.init_file = "meminit.hex";
defparam ram_block3a58.init_file_layout = "port_a";
defparam ram_block3a58.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a58.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a58.operation_mode = "bidir_dual_port";
defparam ram_block3a58.port_a_address_clear = "none";
defparam ram_block3a58.port_a_address_width = 13;
defparam ram_block3a58.port_a_byte_enable_clock = "none";
defparam ram_block3a58.port_a_data_out_clear = "none";
defparam ram_block3a58.port_a_data_out_clock = "none";
defparam ram_block3a58.port_a_data_width = 1;
defparam ram_block3a58.port_a_first_address = 0;
defparam ram_block3a58.port_a_first_bit_number = 26;
defparam ram_block3a58.port_a_last_address = 8191;
defparam ram_block3a58.port_a_logical_ram_depth = 16384;
defparam ram_block3a58.port_a_logical_ram_width = 32;
defparam ram_block3a58.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_address_clear = "none";
defparam ram_block3a58.port_b_address_clock = "clock1";
defparam ram_block3a58.port_b_address_width = 13;
defparam ram_block3a58.port_b_data_in_clock = "clock1";
defparam ram_block3a58.port_b_data_out_clear = "none";
defparam ram_block3a58.port_b_data_out_clock = "none";
defparam ram_block3a58.port_b_data_width = 1;
defparam ram_block3a58.port_b_first_address = 0;
defparam ram_block3a58.port_b_first_bit_number = 26;
defparam ram_block3a58.port_b_last_address = 8191;
defparam ram_block3a58.port_b_logical_ram_depth = 16384;
defparam ram_block3a58.port_b_logical_ram_width = 32;
defparam ram_block3a58.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_read_enable_clock = "clock1";
defparam ram_block3a58.port_b_write_enable_clock = "clock1";
defparam ram_block3a58.ram_block_type = "M9K";
defparam ram_block3a58.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y31_N0
cycloneive_ram_block ram_block3a26(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a26_PORTADATAOUT_bus),
	.portbdataout(ram_block3a26_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a26.clk0_core_clock_enable = "ena0";
defparam ram_block3a26.clk1_core_clock_enable = "ena1";
defparam ram_block3a26.data_interleave_offset_in_bits = 1;
defparam ram_block3a26.data_interleave_width_in_bits = 1;
defparam ram_block3a26.init_file = "meminit.hex";
defparam ram_block3a26.init_file_layout = "port_a";
defparam ram_block3a26.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a26.operation_mode = "bidir_dual_port";
defparam ram_block3a26.port_a_address_clear = "none";
defparam ram_block3a26.port_a_address_width = 13;
defparam ram_block3a26.port_a_byte_enable_clock = "none";
defparam ram_block3a26.port_a_data_out_clear = "none";
defparam ram_block3a26.port_a_data_out_clock = "none";
defparam ram_block3a26.port_a_data_width = 1;
defparam ram_block3a26.port_a_first_address = 0;
defparam ram_block3a26.port_a_first_bit_number = 26;
defparam ram_block3a26.port_a_last_address = 8191;
defparam ram_block3a26.port_a_logical_ram_depth = 16384;
defparam ram_block3a26.port_a_logical_ram_width = 32;
defparam ram_block3a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_address_clear = "none";
defparam ram_block3a26.port_b_address_clock = "clock1";
defparam ram_block3a26.port_b_address_width = 13;
defparam ram_block3a26.port_b_data_in_clock = "clock1";
defparam ram_block3a26.port_b_data_out_clear = "none";
defparam ram_block3a26.port_b_data_out_clock = "none";
defparam ram_block3a26.port_b_data_width = 1;
defparam ram_block3a26.port_b_first_address = 0;
defparam ram_block3a26.port_b_first_bit_number = 26;
defparam ram_block3a26.port_b_last_address = 8191;
defparam ram_block3a26.port_b_logical_ram_depth = 16384;
defparam ram_block3a26.port_b_logical_ram_width = 32;
defparam ram_block3a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_read_enable_clock = "clock1";
defparam ram_block3a26.port_b_write_enable_clock = "clock1";
defparam ram_block3a26.ram_block_type = "M9K";
defparam ram_block3a26.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FF810F;
// synopsys translate_on

// Location: M9K_X64_Y32_N0
cycloneive_ram_block ram_block3a59(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a59_PORTADATAOUT_bus),
	.portbdataout(ram_block3a59_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a59.clk0_core_clock_enable = "ena0";
defparam ram_block3a59.clk1_core_clock_enable = "ena1";
defparam ram_block3a59.data_interleave_offset_in_bits = 1;
defparam ram_block3a59.data_interleave_width_in_bits = 1;
defparam ram_block3a59.init_file = "meminit.hex";
defparam ram_block3a59.init_file_layout = "port_a";
defparam ram_block3a59.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a59.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a59.operation_mode = "bidir_dual_port";
defparam ram_block3a59.port_a_address_clear = "none";
defparam ram_block3a59.port_a_address_width = 13;
defparam ram_block3a59.port_a_byte_enable_clock = "none";
defparam ram_block3a59.port_a_data_out_clear = "none";
defparam ram_block3a59.port_a_data_out_clock = "none";
defparam ram_block3a59.port_a_data_width = 1;
defparam ram_block3a59.port_a_first_address = 0;
defparam ram_block3a59.port_a_first_bit_number = 27;
defparam ram_block3a59.port_a_last_address = 8191;
defparam ram_block3a59.port_a_logical_ram_depth = 16384;
defparam ram_block3a59.port_a_logical_ram_width = 32;
defparam ram_block3a59.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_address_clear = "none";
defparam ram_block3a59.port_b_address_clock = "clock1";
defparam ram_block3a59.port_b_address_width = 13;
defparam ram_block3a59.port_b_data_in_clock = "clock1";
defparam ram_block3a59.port_b_data_out_clear = "none";
defparam ram_block3a59.port_b_data_out_clock = "none";
defparam ram_block3a59.port_b_data_width = 1;
defparam ram_block3a59.port_b_first_address = 0;
defparam ram_block3a59.port_b_first_bit_number = 27;
defparam ram_block3a59.port_b_last_address = 8191;
defparam ram_block3a59.port_b_logical_ram_depth = 16384;
defparam ram_block3a59.port_b_logical_ram_width = 32;
defparam ram_block3a59.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_read_enable_clock = "clock1";
defparam ram_block3a59.port_b_write_enable_clock = "clock1";
defparam ram_block3a59.ram_block_type = "M9K";
defparam ram_block3a59.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y31_N0
cycloneive_ram_block ram_block3a27(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a27_PORTADATAOUT_bus),
	.portbdataout(ram_block3a27_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a27.clk0_core_clock_enable = "ena0";
defparam ram_block3a27.clk1_core_clock_enable = "ena1";
defparam ram_block3a27.data_interleave_offset_in_bits = 1;
defparam ram_block3a27.data_interleave_width_in_bits = 1;
defparam ram_block3a27.init_file = "meminit.hex";
defparam ram_block3a27.init_file_layout = "port_a";
defparam ram_block3a27.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a27.operation_mode = "bidir_dual_port";
defparam ram_block3a27.port_a_address_clear = "none";
defparam ram_block3a27.port_a_address_width = 13;
defparam ram_block3a27.port_a_byte_enable_clock = "none";
defparam ram_block3a27.port_a_data_out_clear = "none";
defparam ram_block3a27.port_a_data_out_clock = "none";
defparam ram_block3a27.port_a_data_width = 1;
defparam ram_block3a27.port_a_first_address = 0;
defparam ram_block3a27.port_a_first_bit_number = 27;
defparam ram_block3a27.port_a_last_address = 8191;
defparam ram_block3a27.port_a_logical_ram_depth = 16384;
defparam ram_block3a27.port_a_logical_ram_width = 32;
defparam ram_block3a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_address_clear = "none";
defparam ram_block3a27.port_b_address_clock = "clock1";
defparam ram_block3a27.port_b_address_width = 13;
defparam ram_block3a27.port_b_data_in_clock = "clock1";
defparam ram_block3a27.port_b_data_out_clear = "none";
defparam ram_block3a27.port_b_data_out_clock = "none";
defparam ram_block3a27.port_b_data_width = 1;
defparam ram_block3a27.port_b_first_address = 0;
defparam ram_block3a27.port_b_first_bit_number = 27;
defparam ram_block3a27.port_b_last_address = 8191;
defparam ram_block3a27.port_b_logical_ram_depth = 16384;
defparam ram_block3a27.port_b_logical_ram_width = 32;
defparam ram_block3a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_read_enable_clock = "clock1";
defparam ram_block3a27.port_b_write_enable_clock = "clock1";
defparam ram_block3a27.ram_block_type = "M9K";
defparam ram_block3a27.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FF8800;
// synopsys translate_on

// Location: M9K_X51_Y41_N0
cycloneive_ram_block ram_block3a60(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a60_PORTADATAOUT_bus),
	.portbdataout(ram_block3a60_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a60.clk0_core_clock_enable = "ena0";
defparam ram_block3a60.clk1_core_clock_enable = "ena1";
defparam ram_block3a60.data_interleave_offset_in_bits = 1;
defparam ram_block3a60.data_interleave_width_in_bits = 1;
defparam ram_block3a60.init_file = "meminit.hex";
defparam ram_block3a60.init_file_layout = "port_a";
defparam ram_block3a60.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a60.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a60.operation_mode = "bidir_dual_port";
defparam ram_block3a60.port_a_address_clear = "none";
defparam ram_block3a60.port_a_address_width = 13;
defparam ram_block3a60.port_a_byte_enable_clock = "none";
defparam ram_block3a60.port_a_data_out_clear = "none";
defparam ram_block3a60.port_a_data_out_clock = "none";
defparam ram_block3a60.port_a_data_width = 1;
defparam ram_block3a60.port_a_first_address = 0;
defparam ram_block3a60.port_a_first_bit_number = 28;
defparam ram_block3a60.port_a_last_address = 8191;
defparam ram_block3a60.port_a_logical_ram_depth = 16384;
defparam ram_block3a60.port_a_logical_ram_width = 32;
defparam ram_block3a60.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_address_clear = "none";
defparam ram_block3a60.port_b_address_clock = "clock1";
defparam ram_block3a60.port_b_address_width = 13;
defparam ram_block3a60.port_b_data_in_clock = "clock1";
defparam ram_block3a60.port_b_data_out_clear = "none";
defparam ram_block3a60.port_b_data_out_clock = "none";
defparam ram_block3a60.port_b_data_width = 1;
defparam ram_block3a60.port_b_first_address = 0;
defparam ram_block3a60.port_b_first_bit_number = 28;
defparam ram_block3a60.port_b_last_address = 8191;
defparam ram_block3a60.port_b_logical_ram_depth = 16384;
defparam ram_block3a60.port_b_logical_ram_width = 32;
defparam ram_block3a60.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_read_enable_clock = "clock1";
defparam ram_block3a60.port_b_write_enable_clock = "clock1";
defparam ram_block3a60.ram_block_type = "M9K";
defparam ram_block3a60.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y38_N0
cycloneive_ram_block ram_block3a28(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a28_PORTADATAOUT_bus),
	.portbdataout(ram_block3a28_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a28.clk0_core_clock_enable = "ena0";
defparam ram_block3a28.clk1_core_clock_enable = "ena1";
defparam ram_block3a28.data_interleave_offset_in_bits = 1;
defparam ram_block3a28.data_interleave_width_in_bits = 1;
defparam ram_block3a28.init_file = "meminit.hex";
defparam ram_block3a28.init_file_layout = "port_a";
defparam ram_block3a28.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a28.operation_mode = "bidir_dual_port";
defparam ram_block3a28.port_a_address_clear = "none";
defparam ram_block3a28.port_a_address_width = 13;
defparam ram_block3a28.port_a_byte_enable_clock = "none";
defparam ram_block3a28.port_a_data_out_clear = "none";
defparam ram_block3a28.port_a_data_out_clock = "none";
defparam ram_block3a28.port_a_data_width = 1;
defparam ram_block3a28.port_a_first_address = 0;
defparam ram_block3a28.port_a_first_bit_number = 28;
defparam ram_block3a28.port_a_last_address = 8191;
defparam ram_block3a28.port_a_logical_ram_depth = 16384;
defparam ram_block3a28.port_a_logical_ram_width = 32;
defparam ram_block3a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_address_clear = "none";
defparam ram_block3a28.port_b_address_clock = "clock1";
defparam ram_block3a28.port_b_address_width = 13;
defparam ram_block3a28.port_b_data_in_clock = "clock1";
defparam ram_block3a28.port_b_data_out_clear = "none";
defparam ram_block3a28.port_b_data_out_clock = "none";
defparam ram_block3a28.port_b_data_width = 1;
defparam ram_block3a28.port_b_first_address = 0;
defparam ram_block3a28.port_b_first_bit_number = 28;
defparam ram_block3a28.port_b_last_address = 8191;
defparam ram_block3a28.port_b_logical_ram_depth = 16384;
defparam ram_block3a28.port_b_logical_ram_width = 32;
defparam ram_block3a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_read_enable_clock = "clock1";
defparam ram_block3a28.port_b_write_enable_clock = "clock1";
defparam ram_block3a28.ram_block_type = "M9K";
defparam ram_block3a28.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000400084F;
// synopsys translate_on

// Location: M9K_X64_Y23_N0
cycloneive_ram_block ram_block3a61(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a61_PORTADATAOUT_bus),
	.portbdataout(ram_block3a61_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a61.clk0_core_clock_enable = "ena0";
defparam ram_block3a61.clk1_core_clock_enable = "ena1";
defparam ram_block3a61.data_interleave_offset_in_bits = 1;
defparam ram_block3a61.data_interleave_width_in_bits = 1;
defparam ram_block3a61.init_file = "meminit.hex";
defparam ram_block3a61.init_file_layout = "port_a";
defparam ram_block3a61.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a61.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a61.operation_mode = "bidir_dual_port";
defparam ram_block3a61.port_a_address_clear = "none";
defparam ram_block3a61.port_a_address_width = 13;
defparam ram_block3a61.port_a_byte_enable_clock = "none";
defparam ram_block3a61.port_a_data_out_clear = "none";
defparam ram_block3a61.port_a_data_out_clock = "none";
defparam ram_block3a61.port_a_data_width = 1;
defparam ram_block3a61.port_a_first_address = 0;
defparam ram_block3a61.port_a_first_bit_number = 29;
defparam ram_block3a61.port_a_last_address = 8191;
defparam ram_block3a61.port_a_logical_ram_depth = 16384;
defparam ram_block3a61.port_a_logical_ram_width = 32;
defparam ram_block3a61.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_address_clear = "none";
defparam ram_block3a61.port_b_address_clock = "clock1";
defparam ram_block3a61.port_b_address_width = 13;
defparam ram_block3a61.port_b_data_in_clock = "clock1";
defparam ram_block3a61.port_b_data_out_clear = "none";
defparam ram_block3a61.port_b_data_out_clock = "none";
defparam ram_block3a61.port_b_data_width = 1;
defparam ram_block3a61.port_b_first_address = 0;
defparam ram_block3a61.port_b_first_bit_number = 29;
defparam ram_block3a61.port_b_last_address = 8191;
defparam ram_block3a61.port_b_logical_ram_depth = 16384;
defparam ram_block3a61.port_b_logical_ram_width = 32;
defparam ram_block3a61.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_read_enable_clock = "clock1";
defparam ram_block3a61.port_b_write_enable_clock = "clock1";
defparam ram_block3a61.ram_block_type = "M9K";
defparam ram_block3a61.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y37_N0
cycloneive_ram_block ram_block3a29(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a29_PORTADATAOUT_bus),
	.portbdataout(ram_block3a29_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a29.clk0_core_clock_enable = "ena0";
defparam ram_block3a29.clk1_core_clock_enable = "ena1";
defparam ram_block3a29.data_interleave_offset_in_bits = 1;
defparam ram_block3a29.data_interleave_width_in_bits = 1;
defparam ram_block3a29.init_file = "meminit.hex";
defparam ram_block3a29.init_file_layout = "port_a";
defparam ram_block3a29.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a29.operation_mode = "bidir_dual_port";
defparam ram_block3a29.port_a_address_clear = "none";
defparam ram_block3a29.port_a_address_width = 13;
defparam ram_block3a29.port_a_byte_enable_clock = "none";
defparam ram_block3a29.port_a_data_out_clear = "none";
defparam ram_block3a29.port_a_data_out_clock = "none";
defparam ram_block3a29.port_a_data_width = 1;
defparam ram_block3a29.port_a_first_address = 0;
defparam ram_block3a29.port_a_first_bit_number = 29;
defparam ram_block3a29.port_a_last_address = 8191;
defparam ram_block3a29.port_a_logical_ram_depth = 16384;
defparam ram_block3a29.port_a_logical_ram_width = 32;
defparam ram_block3a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_address_clear = "none";
defparam ram_block3a29.port_b_address_clock = "clock1";
defparam ram_block3a29.port_b_address_width = 13;
defparam ram_block3a29.port_b_data_in_clock = "clock1";
defparam ram_block3a29.port_b_data_out_clear = "none";
defparam ram_block3a29.port_b_data_out_clock = "none";
defparam ram_block3a29.port_b_data_width = 1;
defparam ram_block3a29.port_b_first_address = 0;
defparam ram_block3a29.port_b_first_bit_number = 29;
defparam ram_block3a29.port_b_last_address = 8191;
defparam ram_block3a29.port_b_logical_ram_depth = 16384;
defparam ram_block3a29.port_b_logical_ram_width = 32;
defparam ram_block3a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_read_enable_clock = "clock1";
defparam ram_block3a29.port_b_write_enable_clock = "clock1";
defparam ram_block3a29.ram_block_type = "M9K";
defparam ram_block3a29.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FF894F;
// synopsys translate_on

// Location: M9K_X64_Y41_N0
cycloneive_ram_block ram_block3a62(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a62_PORTADATAOUT_bus),
	.portbdataout(ram_block3a62_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a62.clk0_core_clock_enable = "ena0";
defparam ram_block3a62.clk1_core_clock_enable = "ena1";
defparam ram_block3a62.data_interleave_offset_in_bits = 1;
defparam ram_block3a62.data_interleave_width_in_bits = 1;
defparam ram_block3a62.init_file = "meminit.hex";
defparam ram_block3a62.init_file_layout = "port_a";
defparam ram_block3a62.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a62.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a62.operation_mode = "bidir_dual_port";
defparam ram_block3a62.port_a_address_clear = "none";
defparam ram_block3a62.port_a_address_width = 13;
defparam ram_block3a62.port_a_byte_enable_clock = "none";
defparam ram_block3a62.port_a_data_out_clear = "none";
defparam ram_block3a62.port_a_data_out_clock = "none";
defparam ram_block3a62.port_a_data_width = 1;
defparam ram_block3a62.port_a_first_address = 0;
defparam ram_block3a62.port_a_first_bit_number = 30;
defparam ram_block3a62.port_a_last_address = 8191;
defparam ram_block3a62.port_a_logical_ram_depth = 16384;
defparam ram_block3a62.port_a_logical_ram_width = 32;
defparam ram_block3a62.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_address_clear = "none";
defparam ram_block3a62.port_b_address_clock = "clock1";
defparam ram_block3a62.port_b_address_width = 13;
defparam ram_block3a62.port_b_data_in_clock = "clock1";
defparam ram_block3a62.port_b_data_out_clear = "none";
defparam ram_block3a62.port_b_data_out_clock = "none";
defparam ram_block3a62.port_b_data_width = 1;
defparam ram_block3a62.port_b_first_address = 0;
defparam ram_block3a62.port_b_first_bit_number = 30;
defparam ram_block3a62.port_b_last_address = 8191;
defparam ram_block3a62.port_b_logical_ram_depth = 16384;
defparam ram_block3a62.port_b_logical_ram_width = 32;
defparam ram_block3a62.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_read_enable_clock = "clock1";
defparam ram_block3a62.port_b_write_enable_clock = "clock1";
defparam ram_block3a62.ram_block_type = "M9K";
defparam ram_block3a62.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y43_N0
cycloneive_ram_block ram_block3a30(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a30_PORTADATAOUT_bus),
	.portbdataout(ram_block3a30_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a30.clk0_core_clock_enable = "ena0";
defparam ram_block3a30.clk1_core_clock_enable = "ena1";
defparam ram_block3a30.data_interleave_offset_in_bits = 1;
defparam ram_block3a30.data_interleave_width_in_bits = 1;
defparam ram_block3a30.init_file = "meminit.hex";
defparam ram_block3a30.init_file_layout = "port_a";
defparam ram_block3a30.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a30.operation_mode = "bidir_dual_port";
defparam ram_block3a30.port_a_address_clear = "none";
defparam ram_block3a30.port_a_address_width = 13;
defparam ram_block3a30.port_a_byte_enable_clock = "none";
defparam ram_block3a30.port_a_data_out_clear = "none";
defparam ram_block3a30.port_a_data_out_clock = "none";
defparam ram_block3a30.port_a_data_width = 1;
defparam ram_block3a30.port_a_first_address = 0;
defparam ram_block3a30.port_a_first_bit_number = 30;
defparam ram_block3a30.port_a_last_address = 8191;
defparam ram_block3a30.port_a_logical_ram_depth = 16384;
defparam ram_block3a30.port_a_logical_ram_width = 32;
defparam ram_block3a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_address_clear = "none";
defparam ram_block3a30.port_b_address_clock = "clock1";
defparam ram_block3a30.port_b_address_width = 13;
defparam ram_block3a30.port_b_data_in_clock = "clock1";
defparam ram_block3a30.port_b_data_out_clear = "none";
defparam ram_block3a30.port_b_data_out_clock = "none";
defparam ram_block3a30.port_b_data_width = 1;
defparam ram_block3a30.port_b_first_address = 0;
defparam ram_block3a30.port_b_first_bit_number = 30;
defparam ram_block3a30.port_b_last_address = 8191;
defparam ram_block3a30.port_b_logical_ram_depth = 16384;
defparam ram_block3a30.port_b_logical_ram_width = 32;
defparam ram_block3a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_read_enable_clock = "clock1";
defparam ram_block3a30.port_b_write_enable_clock = "clock1";
defparam ram_block3a30.ram_block_type = "M9K";
defparam ram_block3a30.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004000000;
// synopsys translate_on

// Location: M9K_X51_Y27_N0
cycloneive_ram_block ram_block3a63(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a63_PORTADATAOUT_bus),
	.portbdataout(ram_block3a63_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a63.clk0_core_clock_enable = "ena0";
defparam ram_block3a63.clk1_core_clock_enable = "ena1";
defparam ram_block3a63.data_interleave_offset_in_bits = 1;
defparam ram_block3a63.data_interleave_width_in_bits = 1;
defparam ram_block3a63.init_file = "meminit.hex";
defparam ram_block3a63.init_file_layout = "port_a";
defparam ram_block3a63.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a63.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a63.operation_mode = "bidir_dual_port";
defparam ram_block3a63.port_a_address_clear = "none";
defparam ram_block3a63.port_a_address_width = 13;
defparam ram_block3a63.port_a_byte_enable_clock = "none";
defparam ram_block3a63.port_a_data_out_clear = "none";
defparam ram_block3a63.port_a_data_out_clock = "none";
defparam ram_block3a63.port_a_data_width = 1;
defparam ram_block3a63.port_a_first_address = 0;
defparam ram_block3a63.port_a_first_bit_number = 31;
defparam ram_block3a63.port_a_last_address = 8191;
defparam ram_block3a63.port_a_logical_ram_depth = 16384;
defparam ram_block3a63.port_a_logical_ram_width = 32;
defparam ram_block3a63.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_address_clear = "none";
defparam ram_block3a63.port_b_address_clock = "clock1";
defparam ram_block3a63.port_b_address_width = 13;
defparam ram_block3a63.port_b_data_in_clock = "clock1";
defparam ram_block3a63.port_b_data_out_clear = "none";
defparam ram_block3a63.port_b_data_out_clock = "none";
defparam ram_block3a63.port_b_data_width = 1;
defparam ram_block3a63.port_b_first_address = 0;
defparam ram_block3a63.port_b_first_bit_number = 31;
defparam ram_block3a63.port_b_last_address = 8191;
defparam ram_block3a63.port_b_logical_ram_depth = 16384;
defparam ram_block3a63.port_b_logical_ram_width = 32;
defparam ram_block3a63.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_read_enable_clock = "clock1";
defparam ram_block3a63.port_b_write_enable_clock = "clock1";
defparam ram_block3a63.ram_block_type = "M9K";
defparam ram_block3a63.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y30_N0
cycloneive_ram_block ram_block3a31(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a31_PORTADATAOUT_bus),
	.portbdataout(ram_block3a31_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a31.clk0_core_clock_enable = "ena0";
defparam ram_block3a31.clk1_core_clock_enable = "ena1";
defparam ram_block3a31.data_interleave_offset_in_bits = 1;
defparam ram_block3a31.data_interleave_width_in_bits = 1;
defparam ram_block3a31.init_file = "meminit.hex";
defparam ram_block3a31.init_file_layout = "port_a";
defparam ram_block3a31.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a31.operation_mode = "bidir_dual_port";
defparam ram_block3a31.port_a_address_clear = "none";
defparam ram_block3a31.port_a_address_width = 13;
defparam ram_block3a31.port_a_byte_enable_clock = "none";
defparam ram_block3a31.port_a_data_out_clear = "none";
defparam ram_block3a31.port_a_data_out_clock = "none";
defparam ram_block3a31.port_a_data_width = 1;
defparam ram_block3a31.port_a_first_address = 0;
defparam ram_block3a31.port_a_first_bit_number = 31;
defparam ram_block3a31.port_a_last_address = 8191;
defparam ram_block3a31.port_a_logical_ram_depth = 16384;
defparam ram_block3a31.port_a_logical_ram_width = 32;
defparam ram_block3a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_address_clear = "none";
defparam ram_block3a31.port_b_address_clock = "clock1";
defparam ram_block3a31.port_b_address_width = 13;
defparam ram_block3a31.port_b_data_in_clock = "clock1";
defparam ram_block3a31.port_b_data_out_clear = "none";
defparam ram_block3a31.port_b_data_out_clock = "none";
defparam ram_block3a31.port_b_data_width = 1;
defparam ram_block3a31.port_b_first_address = 0;
defparam ram_block3a31.port_b_first_bit_number = 31;
defparam ram_block3a31.port_b_last_address = 8191;
defparam ram_block3a31.port_b_logical_ram_depth = 16384;
defparam ram_block3a31.port_b_logical_ram_width = 32;
defparam ram_block3a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_read_enable_clock = "clock1";
defparam ram_block3a31.port_b_write_enable_clock = "clock1";
defparam ram_block3a31.ram_block_type = "M9K";
defparam ram_block3a31.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FF8000;
// synopsys translate_on

// Location: FF_X55_Y35_N5
dffeas \address_reg_a[0] (
	.clk(clock0),
	.d(gnd),
	.asdata(ramaddr1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_a_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_a[0] .is_wysiwyg = "true";
defparam \address_reg_a[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N21
dffeas \address_reg_b[0] (
	.clk(clock1),
	.d(\address_reg_b[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_b_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_b[0] .is_wysiwyg = "true";
defparam \address_reg_b[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N20
cycloneive_lcell_comb \address_reg_b[0]~feeder (
// Equation(s):
// \address_reg_b[0]~feeder_combout  = ram_rom_addr_reg_13

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_13),
	.cin(gnd),
	.combout(\address_reg_b[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \address_reg_b[0]~feeder .lut_mask = 16'hFF00;
defparam \address_reg_b[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa (
	ramaddr,
	always1,
	ramWEN,
	eq_node_1,
	eq_node_0,
	devpor,
	devclrn,
	devoe);
input 	ramaddr;
input 	always1;
input 	ramWEN;
output 	eq_node_1;
output 	eq_node_0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X55_Y32_N8
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (!\ramaddr~29_combout  & (!\ramWEN~0_combout  & always11))

	.dataa(gnd),
	.datab(ramaddr),
	.datac(ramWEN),
	.datad(always1),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h0300;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N14
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (\ramaddr~29_combout  & (!\ramWEN~0_combout  & always11))

	.dataa(gnd),
	.datab(ramaddr),
	.datac(ramWEN),
	.datad(always1),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h0C00;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa_1 (
	ram_rom_addr_reg_13,
	sdr,
	eq_node_1,
	eq_node_0,
	irf_reg_2_1,
	state_5,
	devpor,
	devclrn,
	devoe);
input 	ram_rom_addr_reg_13;
input 	sdr;
output 	eq_node_1;
output 	eq_node_0;
input 	irf_reg_2_1;
input 	state_5;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X47_Y34_N30
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q  & (ram_rom_addr_reg_13 & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5] & sdr)))

	.dataa(irf_reg_2_1),
	.datab(ram_rom_addr_reg_13),
	.datac(state_5),
	.datad(sdr),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h8000;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N16
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q  & (!ram_rom_addr_reg_13 & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5] & sdr)))

	.dataa(irf_reg_2_1),
	.datab(ram_rom_addr_reg_13),
	.datac(state_5),
	.datad(sdr),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h2000;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_mod_ram_rom (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg1,
	ram_rom_data_reg_0,
	ram_rom_addr_reg_13,
	ram_rom_addr_reg_0,
	ram_rom_addr_reg_1,
	ram_rom_addr_reg_2,
	ram_rom_addr_reg_3,
	ram_rom_addr_reg_4,
	ram_rom_addr_reg_5,
	ram_rom_addr_reg_6,
	ram_rom_addr_reg_7,
	ram_rom_addr_reg_8,
	ram_rom_addr_reg_9,
	ram_rom_addr_reg_10,
	ram_rom_addr_reg_11,
	ram_rom_addr_reg_12,
	ram_rom_data_reg_1,
	ram_rom_data_reg_2,
	ram_rom_data_reg_3,
	ram_rom_data_reg_4,
	ram_rom_data_reg_5,
	ram_rom_data_reg_6,
	ram_rom_data_reg_7,
	ram_rom_data_reg_8,
	ram_rom_data_reg_9,
	ram_rom_data_reg_10,
	ram_rom_data_reg_11,
	ram_rom_data_reg_12,
	ram_rom_data_reg_13,
	ram_rom_data_reg_14,
	ram_rom_data_reg_15,
	ram_rom_data_reg_16,
	ram_rom_data_reg_17,
	ram_rom_data_reg_18,
	ram_rom_data_reg_19,
	ram_rom_data_reg_20,
	ram_rom_data_reg_21,
	ram_rom_data_reg_22,
	ram_rom_data_reg_23,
	ram_rom_data_reg_24,
	ram_rom_data_reg_25,
	ram_rom_data_reg_26,
	ram_rom_data_reg_27,
	ram_rom_data_reg_28,
	ram_rom_data_reg_29,
	ram_rom_data_reg_30,
	ram_rom_data_reg_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	sdr,
	address_reg_b_0,
	altera_internal_jtag,
	state_4,
	ir_in,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_4_1,
	node_ena_1,
	clr,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	raw_tck,
	devpor,
	devclrn,
	devoe);
input 	ram_block3a32;
input 	ram_block3a0;
input 	ram_block3a33;
input 	ram_block3a1;
input 	ram_block3a34;
input 	ram_block3a2;
input 	ram_block3a35;
input 	ram_block3a3;
input 	ram_block3a36;
input 	ram_block3a4;
input 	ram_block3a37;
input 	ram_block3a5;
input 	ram_block3a38;
input 	ram_block3a6;
input 	ram_block3a39;
input 	ram_block3a7;
input 	ram_block3a40;
input 	ram_block3a8;
input 	ram_block3a41;
input 	ram_block3a9;
input 	ram_block3a42;
input 	ram_block3a10;
input 	ram_block3a43;
input 	ram_block3a11;
input 	ram_block3a44;
input 	ram_block3a12;
input 	ram_block3a45;
input 	ram_block3a13;
input 	ram_block3a46;
input 	ram_block3a14;
input 	ram_block3a47;
input 	ram_block3a15;
input 	ram_block3a48;
input 	ram_block3a16;
input 	ram_block3a49;
input 	ram_block3a17;
input 	ram_block3a50;
input 	ram_block3a18;
input 	ram_block3a51;
input 	ram_block3a19;
input 	ram_block3a52;
input 	ram_block3a20;
input 	ram_block3a53;
input 	ram_block3a21;
input 	ram_block3a54;
input 	ram_block3a22;
input 	ram_block3a55;
input 	ram_block3a23;
input 	ram_block3a56;
input 	ram_block3a24;
input 	ram_block3a57;
input 	ram_block3a25;
input 	ram_block3a58;
input 	ram_block3a26;
input 	ram_block3a59;
input 	ram_block3a27;
input 	ram_block3a60;
input 	ram_block3a28;
input 	ram_block3a61;
input 	ram_block3a29;
input 	ram_block3a62;
input 	ram_block3a30;
input 	ram_block3a63;
input 	ram_block3a31;
output 	is_in_use_reg1;
output 	ram_rom_data_reg_0;
output 	ram_rom_addr_reg_13;
output 	ram_rom_addr_reg_0;
output 	ram_rom_addr_reg_1;
output 	ram_rom_addr_reg_2;
output 	ram_rom_addr_reg_3;
output 	ram_rom_addr_reg_4;
output 	ram_rom_addr_reg_5;
output 	ram_rom_addr_reg_6;
output 	ram_rom_addr_reg_7;
output 	ram_rom_addr_reg_8;
output 	ram_rom_addr_reg_9;
output 	ram_rom_addr_reg_10;
output 	ram_rom_addr_reg_11;
output 	ram_rom_addr_reg_12;
output 	ram_rom_data_reg_1;
output 	ram_rom_data_reg_2;
output 	ram_rom_data_reg_3;
output 	ram_rom_data_reg_4;
output 	ram_rom_data_reg_5;
output 	ram_rom_data_reg_6;
output 	ram_rom_data_reg_7;
output 	ram_rom_data_reg_8;
output 	ram_rom_data_reg_9;
output 	ram_rom_data_reg_10;
output 	ram_rom_data_reg_11;
output 	ram_rom_data_reg_12;
output 	ram_rom_data_reg_13;
output 	ram_rom_data_reg_14;
output 	ram_rom_data_reg_15;
output 	ram_rom_data_reg_16;
output 	ram_rom_data_reg_17;
output 	ram_rom_data_reg_18;
output 	ram_rom_data_reg_19;
output 	ram_rom_data_reg_20;
output 	ram_rom_data_reg_21;
output 	ram_rom_data_reg_22;
output 	ram_rom_data_reg_23;
output 	ram_rom_data_reg_24;
output 	ram_rom_data_reg_25;
output 	ram_rom_data_reg_26;
output 	ram_rom_data_reg_27;
output 	ram_rom_data_reg_28;
output 	ram_rom_data_reg_29;
output 	ram_rom_data_reg_30;
output 	ram_rom_data_reg_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
output 	sdr;
input 	address_reg_b_0;
input 	altera_internal_jtag;
input 	state_4;
input 	[4:0] ir_in;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	raw_tck;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~6_combout ;
wire \Add1~9 ;
wire \Add1~10_combout ;
wire \ram_rom_data_shift_cntr_reg[3]~8_combout ;
wire \is_in_use_reg~0_combout ;
wire \ram_rom_data_reg[0]~0_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~4_combout ;
wire \Add1~3 ;
wire \Add1~4_combout ;
wire \ram_rom_data_shift_cntr_reg[2]~9_combout ;
wire \Add1~5 ;
wire \Add1~7 ;
wire \Add1~8_combout ;
wire \ram_rom_data_shift_cntr_reg[4]~7_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~12_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~10_combout ;
wire \Equal1~0_combout ;
wire \ram_rom_data_shift_cntr_reg[2]~11_combout ;
wire \Add1~0_combout ;
wire \ram_rom_data_shift_cntr_reg[0]~6_combout ;
wire \Add1~1 ;
wire \Add1~2_combout ;
wire \ram_rom_data_shift_cntr_reg[1]~5_combout ;
wire \Equal1~1_combout ;
wire \process_0~2_combout ;
wire \ram_rom_data_reg[21]~32_combout ;
wire \ram_rom_addr_reg[0]~15 ;
wire \ram_rom_addr_reg[1]~17 ;
wire \ram_rom_addr_reg[2]~19 ;
wire \ram_rom_addr_reg[3]~21 ;
wire \ram_rom_addr_reg[4]~23 ;
wire \ram_rom_addr_reg[5]~25 ;
wire \ram_rom_addr_reg[6]~27 ;
wire \ram_rom_addr_reg[7]~29 ;
wire \ram_rom_addr_reg[8]~31 ;
wire \ram_rom_addr_reg[9]~33 ;
wire \ram_rom_addr_reg[10]~35 ;
wire \ram_rom_addr_reg[11]~37 ;
wire \ram_rom_addr_reg[12]~39 ;
wire \ram_rom_addr_reg[13]~40_combout ;
wire \process_0~3_combout ;
wire \ram_rom_addr_reg[6]~42_combout ;
wire \ram_rom_addr_reg[6]~43_combout ;
wire \ram_rom_addr_reg[0]~14_combout ;
wire \ram_rom_addr_reg[1]~16_combout ;
wire \ram_rom_addr_reg[2]~18_combout ;
wire \ram_rom_addr_reg[3]~20_combout ;
wire \ram_rom_addr_reg[4]~22_combout ;
wire \ram_rom_addr_reg[5]~24_combout ;
wire \ram_rom_addr_reg[6]~26_combout ;
wire \ram_rom_addr_reg[7]~28_combout ;
wire \ram_rom_addr_reg[8]~30_combout ;
wire \ram_rom_addr_reg[9]~32_combout ;
wire \ram_rom_addr_reg[10]~34_combout ;
wire \ram_rom_addr_reg[11]~36_combout ;
wire \ram_rom_addr_reg[12]~38_combout ;
wire \ram_rom_data_reg[1]~1_combout ;
wire \ram_rom_data_reg[2]~2_combout ;
wire \ram_rom_data_reg[3]~3_combout ;
wire \ram_rom_data_reg[4]~4_combout ;
wire \ram_rom_data_reg[5]~5_combout ;
wire \ram_rom_data_reg[6]~6_combout ;
wire \ram_rom_data_reg[7]~7_combout ;
wire \ram_rom_data_reg[8]~8_combout ;
wire \ram_rom_data_reg[9]~9_combout ;
wire \ram_rom_data_reg[10]~10_combout ;
wire \ram_rom_data_reg[11]~11_combout ;
wire \ram_rom_data_reg[12]~12_combout ;
wire \ram_rom_data_reg[13]~13_combout ;
wire \ram_rom_data_reg[14]~14_combout ;
wire \ram_rom_data_reg[15]~15_combout ;
wire \ram_rom_data_reg[16]~16_combout ;
wire \ram_rom_data_reg[17]~17_combout ;
wire \ram_rom_data_reg[18]~18_combout ;
wire \ram_rom_data_reg[19]~19_combout ;
wire \ram_rom_data_reg[20]~20_combout ;
wire \ram_rom_data_reg[21]~21_combout ;
wire \ram_rom_data_reg[22]~22_combout ;
wire \ram_rom_data_reg[23]~23_combout ;
wire \ram_rom_data_reg[24]~24_combout ;
wire \ram_rom_data_reg[25]~25_combout ;
wire \ram_rom_data_reg[26]~26_combout ;
wire \ram_rom_data_reg[27]~27_combout ;
wire \ram_rom_data_reg[28]~28_combout ;
wire \ram_rom_data_reg[29]~29_combout ;
wire \ram_rom_data_reg[30]~30_combout ;
wire \ram_rom_data_reg[31]~31_combout ;
wire \process_0~0_combout ;
wire \process_0~1_combout ;
wire \ir_loaded_address_reg[1]~feeder_combout ;
wire \ir_loaded_address_reg[3]~feeder_combout ;
wire \bypass_reg_out~0_combout ;
wire \bypass_reg_out~q ;
wire \tdo~0_combout ;
wire [5:0] ram_rom_data_shift_cntr_reg;
wire [3:0] \ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR ;


sld_rom_sr \ram_rom_logic_gen:name_gen:info_rom_sr (
	.WORD_SR_0(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.sdr(sdr),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.TCK(raw_tck),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X47_Y35_N18
cycloneive_lcell_comb \Add1~6 (
	.dataa(ram_rom_data_shift_cntr_reg[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h5A5F;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N20
cycloneive_lcell_comb \Add1~8 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'hC30C;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N22
cycloneive_lcell_comb \Add1~10 (
	.dataa(ram_rom_data_shift_cntr_reg[5]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h5A5A;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X47_Y35_N11
dffeas \ram_rom_data_shift_cntr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[3]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N10
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[3]~8 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[2]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[3]),
	.datad(\Add1~6_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3]~8 .lut_mask = 16'hD5C0;
defparam \ram_rom_data_shift_cntr_reg[3]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N9
dffeas is_in_use_reg(
	.clk(raw_tck),
	.d(\is_in_use_reg~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(ir_in[0]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(is_in_use_reg1),
	.prn(vcc));
// synopsys translate_off
defparam is_in_use_reg.is_wysiwyg = "true";
defparam is_in_use_reg.power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N25
dffeas \ram_rom_data_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[0]~0_combout ),
	.asdata(ram_rom_data_reg_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N27
dffeas \ram_rom_addr_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[13]~40_combout ),
	.asdata(altera_internal_jtag),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[6]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N1
dffeas \ram_rom_addr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[0]~14_combout ),
	.asdata(ram_rom_addr_reg_1),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[6]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N3
dffeas \ram_rom_addr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[1]~16_combout ),
	.asdata(ram_rom_addr_reg_2),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[6]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N5
dffeas \ram_rom_addr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[2]~18_combout ),
	.asdata(ram_rom_addr_reg_3),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[6]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N7
dffeas \ram_rom_addr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[3]~20_combout ),
	.asdata(ram_rom_addr_reg_4),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[6]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N9
dffeas \ram_rom_addr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[4]~22_combout ),
	.asdata(ram_rom_addr_reg_5),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[6]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N11
dffeas \ram_rom_addr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[5]~24_combout ),
	.asdata(ram_rom_addr_reg_6),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[6]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N13
dffeas \ram_rom_addr_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[6]~26_combout ),
	.asdata(ram_rom_addr_reg_7),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[6]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N15
dffeas \ram_rom_addr_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[7]~28_combout ),
	.asdata(ram_rom_addr_reg_8),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[6]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N17
dffeas \ram_rom_addr_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[8]~30_combout ),
	.asdata(ram_rom_addr_reg_9),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[6]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N19
dffeas \ram_rom_addr_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[9]~32_combout ),
	.asdata(ram_rom_addr_reg_10),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[6]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N21
dffeas \ram_rom_addr_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[10]~34_combout ),
	.asdata(ram_rom_addr_reg_11),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[6]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N23
dffeas \ram_rom_addr_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[11]~36_combout ),
	.asdata(ram_rom_addr_reg_12),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[6]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X48_Y34_N25
dffeas \ram_rom_addr_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[12]~38_combout ),
	.asdata(ram_rom_addr_reg_13),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[6]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N11
dffeas \ram_rom_data_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[1]~1_combout ),
	.asdata(ram_rom_data_reg_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N21
dffeas \ram_rom_data_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[2]~2_combout ),
	.asdata(ram_rom_data_reg_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N27
dffeas \ram_rom_data_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[3]~3_combout ),
	.asdata(ram_rom_data_reg_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N13
dffeas \ram_rom_data_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[4]~4_combout ),
	.asdata(ram_rom_data_reg_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N23
dffeas \ram_rom_data_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[5]~5_combout ),
	.asdata(ram_rom_data_reg_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N9
dffeas \ram_rom_data_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[6]~6_combout ),
	.asdata(ram_rom_data_reg_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N31
dffeas \ram_rom_data_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[7]~7_combout ),
	.asdata(ram_rom_data_reg_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N17
dffeas \ram_rom_data_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[8]~8_combout ),
	.asdata(ram_rom_data_reg_9),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N15
dffeas \ram_rom_data_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[9]~9_combout ),
	.asdata(ram_rom_data_reg_10),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N25
dffeas \ram_rom_data_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[10]~10_combout ),
	.asdata(ram_rom_data_reg_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N27
dffeas \ram_rom_data_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[11]~11_combout ),
	.asdata(ram_rom_data_reg_12),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N9
dffeas \ram_rom_data_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[12]~12_combout ),
	.asdata(ram_rom_data_reg_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N7
dffeas \ram_rom_data_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[13]~13_combout ),
	.asdata(ram_rom_data_reg_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N5
dffeas \ram_rom_data_reg[14] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[14]~14_combout ),
	.asdata(ram_rom_data_reg_15),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_14),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[14] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N11
dffeas \ram_rom_data_reg[15] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[15]~15_combout ),
	.asdata(ram_rom_data_reg_16),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_15),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[15] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N13
dffeas \ram_rom_data_reg[16] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[16]~16_combout ),
	.asdata(ram_rom_data_reg_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_16),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[16] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N23
dffeas \ram_rom_data_reg[17] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[17]~17_combout ),
	.asdata(ram_rom_data_reg_18),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_17),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[17] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N17
dffeas \ram_rom_data_reg[18] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[18]~18_combout ),
	.asdata(ram_rom_data_reg_19),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_18),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[18] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N15
dffeas \ram_rom_data_reg[19] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[19]~19_combout ),
	.asdata(ram_rom_data_reg_20),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_19),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[19] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N13
dffeas \ram_rom_data_reg[20] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[20]~20_combout ),
	.asdata(ram_rom_data_reg_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_20),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[20] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N15
dffeas \ram_rom_data_reg[21] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[21]~21_combout ),
	.asdata(ram_rom_data_reg_22),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_21),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[21] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N21
dffeas \ram_rom_data_reg[22] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[22]~22_combout ),
	.asdata(ram_rom_data_reg_23),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_22),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[22] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N19
dffeas \ram_rom_data_reg[23] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[23]~23_combout ),
	.asdata(ram_rom_data_reg_24),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_23),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[23] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N17
dffeas \ram_rom_data_reg[24] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[24]~24_combout ),
	.asdata(ram_rom_data_reg_25),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_24),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[24] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N27
dffeas \ram_rom_data_reg[25] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[25]~25_combout ),
	.asdata(ram_rom_data_reg_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_25),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[25] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N9
dffeas \ram_rom_data_reg[26] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[26]~26_combout ),
	.asdata(ram_rom_data_reg_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_26),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[26] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N31
dffeas \ram_rom_data_reg[27] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[27]~27_combout ),
	.asdata(ram_rom_data_reg_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_27),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[27] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N25
dffeas \ram_rom_data_reg[28] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[28]~28_combout ),
	.asdata(ram_rom_data_reg_29),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_28),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[28] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N23
dffeas \ram_rom_data_reg[29] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[29]~29_combout ),
	.asdata(ram_rom_data_reg_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_29),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[29] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y38_N29
dffeas \ram_rom_data_reg[30] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[30]~30_combout ),
	.asdata(ram_rom_data_reg_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_30),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[30] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N29
dffeas \ram_rom_data_reg[31] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[31]~31_combout ),
	.asdata(altera_internal_jtag),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[21]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_31),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[31] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y34_N5
dffeas \ir_loaded_address_reg[0] (
	.clk(raw_tck),
	.d(gnd),
	.asdata(ram_rom_addr_reg_0),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[0] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y34_N27
dffeas \ir_loaded_address_reg[1] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[1] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y34_N21
dffeas \ir_loaded_address_reg[2] (
	.clk(raw_tck),
	.d(gnd),
	.asdata(ram_rom_addr_reg_2),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[2] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y34_N23
dffeas \ir_loaded_address_reg[3] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[3] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N2
cycloneive_lcell_comb \tdo~1 (
	.dataa(gnd),
	.datab(ir_in[0]),
	.datac(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.datad(\tdo~0_combout ),
	.cin(gnd),
	.combout(tdo),
	.cout());
// synopsys translate_off
defparam \tdo~1 .lut_mask = 16'hF3C0;
defparam \tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N0
cycloneive_lcell_comb \sdr~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(node_ena_1),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(sdr),
	.cout());
// synopsys translate_off
defparam \sdr~0 .lut_mask = 16'h00F0;
defparam \sdr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N8
cycloneive_lcell_comb \is_in_use_reg~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(is_in_use_reg1),
	.datad(irf_reg_4_1),
	.cin(gnd),
	.combout(\is_in_use_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \is_in_use_reg~0 .lut_mask = 16'h00F0;
defparam \is_in_use_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N24
cycloneive_lcell_comb \ram_rom_data_reg[0]~0 (
	.dataa(ram_block3a32),
	.datab(ram_block3a0),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[0]~0 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N6
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~4 (
	.dataa(irf_reg_1_1),
	.datab(sdr),
	.datac(irf_reg_2_1),
	.datad(state_4),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~4 .lut_mask = 16'hC800;
defparam \ram_rom_data_shift_cntr_reg[5]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N14
cycloneive_lcell_comb \Add1~2 (
	.dataa(ram_rom_data_shift_cntr_reg[1]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h5A5F;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N16
cycloneive_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'hC30C;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N0
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[2]~9 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[2]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[2]),
	.datad(\Add1~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2]~9 .lut_mask = 16'hD5C0;
defparam \ram_rom_data_shift_cntr_reg[2]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y35_N1
dffeas \ram_rom_data_shift_cntr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[2]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N28
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[4]~7 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[2]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[4]),
	.datad(\Add1~8_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4]~7 .lut_mask = 16'hD5C0;
defparam \ram_rom_data_shift_cntr_reg[4]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y35_N29
dffeas \ram_rom_data_shift_cntr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[4]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N6
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~12 (
	.dataa(ram_rom_data_shift_cntr_reg[1]),
	.datab(\Equal1~0_combout ),
	.datac(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datad(ram_rom_data_shift_cntr_reg[0]),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~12 .lut_mask = 16'h8F0F;
defparam \ram_rom_data_shift_cntr_reg[5]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N26
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~10 (
	.dataa(\Add1~10_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[2]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[5]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~10 .lut_mask = 16'hC0EA;
defparam \ram_rom_data_shift_cntr_reg[5]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y35_N27
dffeas \ram_rom_data_shift_cntr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[5]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N24
cycloneive_lcell_comb \Equal1~0 (
	.dataa(ram_rom_data_shift_cntr_reg[3]),
	.datab(ram_rom_data_shift_cntr_reg[4]),
	.datac(ram_rom_data_shift_cntr_reg[5]),
	.datad(ram_rom_data_shift_cntr_reg[2]),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~0 .lut_mask = 16'h0800;
defparam \Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N4
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[2]~11 (
	.dataa(ram_rom_data_shift_cntr_reg[1]),
	.datab(\Equal1~0_combout ),
	.datac(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datad(ram_rom_data_shift_cntr_reg[0]),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[2]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2]~11 .lut_mask = 16'h070F;
defparam \ram_rom_data_shift_cntr_reg[2]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N12
cycloneive_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h33CC;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N2
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[0]~6 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[2]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[0]),
	.datad(\Add1~0_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0]~6 .lut_mask = 16'hD5C0;
defparam \ram_rom_data_shift_cntr_reg[0]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y35_N3
dffeas \ram_rom_data_shift_cntr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[0]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N8
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[1]~5 (
	.dataa(\Equal1~1_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(\Add1~2_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1]~5 .lut_mask = 16'h5C10;
defparam \ram_rom_data_shift_cntr_reg[1]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y35_N9
dffeas \ram_rom_data_shift_cntr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[1]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N30
cycloneive_lcell_comb \Equal1~1 (
	.dataa(gnd),
	.datab(\Equal1~0_combout ),
	.datac(gnd),
	.datad(ram_rom_data_shift_cntr_reg[0]),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~1 .lut_mask = 16'hCC00;
defparam \Equal1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N20
cycloneive_lcell_comb \process_0~2 (
	.dataa(irf_reg_1_1),
	.datab(ram_rom_data_shift_cntr_reg[1]),
	.datac(\Equal1~1_combout ),
	.datad(ir_in[3]),
	.cin(gnd),
	.combout(\process_0~2_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~2 .lut_mask = 16'h007F;
defparam \process_0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N30
cycloneive_lcell_comb \ram_rom_data_reg[21]~32 (
	.dataa(gnd),
	.datab(\process_0~2_combout ),
	.datac(gnd),
	.datad(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_reg[21]~32_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[21]~32 .lut_mask = 16'hFF33;
defparam \ram_rom_data_reg[21]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N0
cycloneive_lcell_comb \ram_rom_addr_reg[0]~14 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[0]~14_combout ),
	.cout(\ram_rom_addr_reg[0]~15 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[0]~14 .lut_mask = 16'h33CC;
defparam \ram_rom_addr_reg[0]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N2
cycloneive_lcell_comb \ram_rom_addr_reg[1]~16 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[0]~15 ),
	.combout(\ram_rom_addr_reg[1]~16_combout ),
	.cout(\ram_rom_addr_reg[1]~17 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[1]~16 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[1]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N4
cycloneive_lcell_comb \ram_rom_addr_reg[2]~18 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[1]~17 ),
	.combout(\ram_rom_addr_reg[2]~18_combout ),
	.cout(\ram_rom_addr_reg[2]~19 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[2]~18 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[2]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N6
cycloneive_lcell_comb \ram_rom_addr_reg[3]~20 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[2]~19 ),
	.combout(\ram_rom_addr_reg[3]~20_combout ),
	.cout(\ram_rom_addr_reg[3]~21 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[3]~20 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[3]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N8
cycloneive_lcell_comb \ram_rom_addr_reg[4]~22 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[3]~21 ),
	.combout(\ram_rom_addr_reg[4]~22_combout ),
	.cout(\ram_rom_addr_reg[4]~23 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[4]~22 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[4]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N10
cycloneive_lcell_comb \ram_rom_addr_reg[5]~24 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[4]~23 ),
	.combout(\ram_rom_addr_reg[5]~24_combout ),
	.cout(\ram_rom_addr_reg[5]~25 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[5]~24 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[5]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N12
cycloneive_lcell_comb \ram_rom_addr_reg[6]~26 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[5]~25 ),
	.combout(\ram_rom_addr_reg[6]~26_combout ),
	.cout(\ram_rom_addr_reg[6]~27 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[6]~26 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[6]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N14
cycloneive_lcell_comb \ram_rom_addr_reg[7]~28 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[6]~27 ),
	.combout(\ram_rom_addr_reg[7]~28_combout ),
	.cout(\ram_rom_addr_reg[7]~29 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[7]~28 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[7]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N16
cycloneive_lcell_comb \ram_rom_addr_reg[8]~30 (
	.dataa(ram_rom_addr_reg_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[7]~29 ),
	.combout(\ram_rom_addr_reg[8]~30_combout ),
	.cout(\ram_rom_addr_reg[8]~31 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[8]~30 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[8]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N18
cycloneive_lcell_comb \ram_rom_addr_reg[9]~32 (
	.dataa(ram_rom_addr_reg_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[8]~31 ),
	.combout(\ram_rom_addr_reg[9]~32_combout ),
	.cout(\ram_rom_addr_reg[9]~33 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[9]~32 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[9]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N20
cycloneive_lcell_comb \ram_rom_addr_reg[10]~34 (
	.dataa(ram_rom_addr_reg_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[9]~33 ),
	.combout(\ram_rom_addr_reg[10]~34_combout ),
	.cout(\ram_rom_addr_reg[10]~35 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[10]~34 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[10]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N22
cycloneive_lcell_comb \ram_rom_addr_reg[11]~36 (
	.dataa(ram_rom_addr_reg_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[10]~35 ),
	.combout(\ram_rom_addr_reg[11]~36_combout ),
	.cout(\ram_rom_addr_reg[11]~37 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[11]~36 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[11]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N24
cycloneive_lcell_comb \ram_rom_addr_reg[12]~38 (
	.dataa(ram_rom_addr_reg_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[11]~37 ),
	.combout(\ram_rom_addr_reg[12]~38_combout ),
	.cout(\ram_rom_addr_reg[12]~39 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[12]~38 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[12]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X48_Y34_N26
cycloneive_lcell_comb \ram_rom_addr_reg[13]~40 (
	.dataa(ram_rom_addr_reg_13),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\ram_rom_addr_reg[12]~39 ),
	.combout(\ram_rom_addr_reg[13]~40_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[13]~40 .lut_mask = 16'h5A5A;
defparam \ram_rom_addr_reg[13]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N28
cycloneive_lcell_comb \process_0~3 (
	.dataa(state_4),
	.datab(virtual_ir_scan_reg),
	.datac(node_ena_1),
	.datad(ir_in[3]),
	.cin(gnd),
	.combout(\process_0~3_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~3 .lut_mask = 16'h2000;
defparam \process_0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N18
cycloneive_lcell_comb \ram_rom_addr_reg[6]~42 (
	.dataa(irf_reg_1_1),
	.datab(\process_0~3_combout ),
	.datac(\Equal1~1_combout ),
	.datad(ram_rom_data_shift_cntr_reg[1]),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[6]~42_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[6]~42 .lut_mask = 16'hCCEC;
defparam \ram_rom_addr_reg[6]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N24
cycloneive_lcell_comb \ram_rom_addr_reg[6]~43 (
	.dataa(irf_reg_2_1),
	.datab(\ram_rom_addr_reg[6]~42_combout ),
	.datac(state_8),
	.datad(sdr),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[6]~43_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[6]~43 .lut_mask = 16'hECCC;
defparam \ram_rom_addr_reg[6]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N10
cycloneive_lcell_comb \ram_rom_data_reg[1]~1 (
	.dataa(ram_block3a33),
	.datab(ram_block3a1),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[1]~1 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N20
cycloneive_lcell_comb \ram_rom_data_reg[2]~2 (
	.dataa(ram_block3a2),
	.datab(ram_block3a34),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[2]~2 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N26
cycloneive_lcell_comb \ram_rom_data_reg[3]~3 (
	.dataa(ram_block3a35),
	.datab(ram_block3a3),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[3]~3 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N12
cycloneive_lcell_comb \ram_rom_data_reg[4]~4 (
	.dataa(ram_block3a4),
	.datab(ram_block3a36),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[4]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[4]~4 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N22
cycloneive_lcell_comb \ram_rom_data_reg[5]~5 (
	.dataa(ram_block3a37),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a5),
	.cin(gnd),
	.combout(\ram_rom_data_reg[5]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[5]~5 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[5]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N8
cycloneive_lcell_comb \ram_rom_data_reg[6]~6 (
	.dataa(ram_block3a38),
	.datab(ram_block3a6),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[6]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[6]~6 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[6]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N30
cycloneive_lcell_comb \ram_rom_data_reg[7]~7 (
	.dataa(ram_block3a7),
	.datab(ram_block3a39),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[7]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[7]~7 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[7]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N16
cycloneive_lcell_comb \ram_rom_data_reg[8]~8 (
	.dataa(ram_block3a8),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a40),
	.cin(gnd),
	.combout(\ram_rom_data_reg[8]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[8]~8 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[8]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N14
cycloneive_lcell_comb \ram_rom_data_reg[9]~9 (
	.dataa(ram_block3a41),
	.datab(ram_block3a9),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[9]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[9]~9 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[9]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N24
cycloneive_lcell_comb \ram_rom_data_reg[10]~10 (
	.dataa(ram_block3a10),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a42),
	.cin(gnd),
	.combout(\ram_rom_data_reg[10]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[10]~10 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[10]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N26
cycloneive_lcell_comb \ram_rom_data_reg[11]~11 (
	.dataa(ram_block3a11),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a43),
	.cin(gnd),
	.combout(\ram_rom_data_reg[11]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[11]~11 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[11]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N8
cycloneive_lcell_comb \ram_rom_data_reg[12]~12 (
	.dataa(ram_block3a12),
	.datab(ram_block3a44),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[12]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[12]~12 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[12]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N6
cycloneive_lcell_comb \ram_rom_data_reg[13]~13 (
	.dataa(ram_block3a45),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a13),
	.cin(gnd),
	.combout(\ram_rom_data_reg[13]~13_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[13]~13 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[13]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N4
cycloneive_lcell_comb \ram_rom_data_reg[14]~14 (
	.dataa(ram_block3a46),
	.datab(ram_block3a14),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[14]~14_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[14]~14 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[14]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N10
cycloneive_lcell_comb \ram_rom_data_reg[15]~15 (
	.dataa(ram_block3a15),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a47),
	.cin(gnd),
	.combout(\ram_rom_data_reg[15]~15_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[15]~15 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[15]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N12
cycloneive_lcell_comb \ram_rom_data_reg[16]~16 (
	.dataa(ram_block3a48),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a16),
	.cin(gnd),
	.combout(\ram_rom_data_reg[16]~16_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[16]~16 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[16]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N22
cycloneive_lcell_comb \ram_rom_data_reg[17]~17 (
	.dataa(ram_block3a17),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a49),
	.cin(gnd),
	.combout(\ram_rom_data_reg[17]~17_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[17]~17 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[17]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N16
cycloneive_lcell_comb \ram_rom_data_reg[18]~18 (
	.dataa(ram_block3a18),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a50),
	.cin(gnd),
	.combout(\ram_rom_data_reg[18]~18_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[18]~18 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[18]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N14
cycloneive_lcell_comb \ram_rom_data_reg[19]~19 (
	.dataa(ram_block3a19),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a51),
	.cin(gnd),
	.combout(\ram_rom_data_reg[19]~19_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[19]~19 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[19]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N12
cycloneive_lcell_comb \ram_rom_data_reg[20]~20 (
	.dataa(ram_block3a52),
	.datab(ram_block3a20),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[20]~20_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[20]~20 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[20]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N14
cycloneive_lcell_comb \ram_rom_data_reg[21]~21 (
	.dataa(ram_block3a53),
	.datab(ram_block3a21),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[21]~21_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[21]~21 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[21]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N20
cycloneive_lcell_comb \ram_rom_data_reg[22]~22 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a22),
	.datac(gnd),
	.datad(ram_block3a54),
	.cin(gnd),
	.combout(\ram_rom_data_reg[22]~22_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[22]~22 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[22]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N18
cycloneive_lcell_comb \ram_rom_data_reg[23]~23 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a23),
	.datac(gnd),
	.datad(ram_block3a55),
	.cin(gnd),
	.combout(\ram_rom_data_reg[23]~23_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[23]~23 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[23]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N16
cycloneive_lcell_comb \ram_rom_data_reg[24]~24 (
	.dataa(ram_block3a24),
	.datab(ram_block3a56),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[24]~24_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[24]~24 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[24]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N26
cycloneive_lcell_comb \ram_rom_data_reg[25]~25 (
	.dataa(ram_block3a57),
	.datab(ram_block3a25),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[25]~25_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[25]~25 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[25]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N8
cycloneive_lcell_comb \ram_rom_data_reg[26]~26 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a26),
	.datac(gnd),
	.datad(ram_block3a58),
	.cin(gnd),
	.combout(\ram_rom_data_reg[26]~26_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[26]~26 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[26]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N30
cycloneive_lcell_comb \ram_rom_data_reg[27]~27 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a27),
	.datac(gnd),
	.datad(ram_block3a59),
	.cin(gnd),
	.combout(\ram_rom_data_reg[27]~27_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[27]~27 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[27]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N24
cycloneive_lcell_comb \ram_rom_data_reg[28]~28 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a28),
	.datac(gnd),
	.datad(ram_block3a60),
	.cin(gnd),
	.combout(\ram_rom_data_reg[28]~28_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[28]~28 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[28]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N22
cycloneive_lcell_comb \ram_rom_data_reg[29]~29 (
	.dataa(ram_block3a29),
	.datab(ram_block3a61),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[29]~29_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[29]~29 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[29]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N28
cycloneive_lcell_comb \ram_rom_data_reg[30]~30 (
	.dataa(ram_block3a62),
	.datab(ram_block3a30),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[30]~30_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[30]~30 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[30]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N28
cycloneive_lcell_comb \ram_rom_data_reg[31]~31 (
	.dataa(ram_block3a31),
	.datab(ram_block3a63),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[31]~31_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[31]~31 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[31]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N12
cycloneive_lcell_comb \process_0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(irf_reg_4_1),
	.datad(ir_in[0]),
	.cin(gnd),
	.combout(\process_0~0_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~0 .lut_mask = 16'hFFF0;
defparam \process_0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N14
cycloneive_lcell_comb \process_0~1 (
	.dataa(state_5),
	.datab(virtual_ir_scan_reg),
	.datac(node_ena_1),
	.datad(ir_in[3]),
	.cin(gnd),
	.combout(\process_0~1_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~1 .lut_mask = 16'h2000;
defparam \process_0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N26
cycloneive_lcell_comb \ir_loaded_address_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_1),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y34_N22
cycloneive_lcell_comb \ir_loaded_address_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_3),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N10
cycloneive_lcell_comb \bypass_reg_out~0 (
	.dataa(altera_internal_jtag),
	.datab(node_ena_1),
	.datac(\bypass_reg_out~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\bypass_reg_out~0_combout ),
	.cout());
// synopsys translate_off
defparam \bypass_reg_out~0 .lut_mask = 16'hB8B8;
defparam \bypass_reg_out~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N11
dffeas bypass_reg_out(
	.clk(raw_tck),
	.d(\bypass_reg_out~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\bypass_reg_out~q ),
	.prn(vcc));
// synopsys translate_off
defparam bypass_reg_out.is_wysiwyg = "true";
defparam bypass_reg_out.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N12
cycloneive_lcell_comb \tdo~0 (
	.dataa(irf_reg_1_1),
	.datab(ram_rom_data_reg_0),
	.datac(irf_reg_2_1),
	.datad(\bypass_reg_out~q ),
	.cin(gnd),
	.combout(\tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \tdo~0 .lut_mask = 16'hCDC8;
defparam \tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_rom_sr (
	WORD_SR_0,
	sdr,
	altera_internal_jtag,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	TCK,
	devpor,
	devclrn,
	devoe);
output 	WORD_SR_0;
input 	sdr;
input 	altera_internal_jtag;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	TCK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \word_counter[1]~9_combout ;
wire \WORD_SR~2_combout ;
wire \WORD_SR~7_combout ;
wire \WORD_SR~13_combout ;
wire \clear_signal~combout ;
wire \word_counter[0]~7_combout ;
wire \word_counter[0]~8 ;
wire \word_counter[1]~10 ;
wire \word_counter[2]~11_combout ;
wire \word_counter[0]~14_combout ;
wire \word_counter[2]~12 ;
wire \word_counter[3]~16 ;
wire \word_counter[4]~17_combout ;
wire \word_counter[3]~15_combout ;
wire \word_counter[0]~13_combout ;
wire \word_counter[0]~19_combout ;
wire \WORD_SR~14_combout ;
wire \WORD_SR~15_combout ;
wire \WORD_SR[3]~6_combout ;
wire \WORD_SR~10_combout ;
wire \WORD_SR~11_combout ;
wire \WORD_SR~12_combout ;
wire \WORD_SR~8_combout ;
wire \WORD_SR~9_combout ;
wire \WORD_SR~3_combout ;
wire \WORD_SR~4_combout ;
wire \WORD_SR~5_combout ;
wire [4:0] word_counter;
wire [3:0] WORD_SR;


// Location: FF_X43_Y34_N23
dffeas \word_counter[1] (
	.clk(TCK),
	.d(\word_counter[1]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[0]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[0]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[1]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[1] .is_wysiwyg = "true";
defparam \word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N22
cycloneive_lcell_comb \word_counter[1]~9 (
	.dataa(word_counter[1]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[0]~8 ),
	.combout(\word_counter[1]~9_combout ),
	.cout(\word_counter[1]~10 ));
// synopsys translate_off
defparam \word_counter[1]~9 .lut_mask = 16'h5A5F;
defparam \word_counter[1]~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X39_Y34_N12
cycloneive_lcell_comb \WORD_SR~2 (
	.dataa(word_counter[1]),
	.datab(word_counter[4]),
	.datac(word_counter[2]),
	.datad(word_counter[3]),
	.cin(gnd),
	.combout(\WORD_SR~2_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~2 .lut_mask = 16'h3005;
defparam \WORD_SR~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N12
cycloneive_lcell_comb \WORD_SR~7 (
	.dataa(state_4),
	.datab(word_counter[4]),
	.datac(word_counter[1]),
	.datad(word_counter[0]),
	.cin(gnd),
	.combout(\WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~7 .lut_mask = 16'h0051;
defparam \WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y34_N10
cycloneive_lcell_comb \WORD_SR~13 (
	.dataa(word_counter[1]),
	.datab(word_counter[4]),
	.datac(word_counter[2]),
	.datad(word_counter[3]),
	.cin(gnd),
	.combout(\WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~13 .lut_mask = 16'h2000;
defparam \WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N1
dffeas \WORD_SR[0] (
	.clk(TCK),
	.d(\WORD_SR~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[3]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR_0),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[0] .is_wysiwyg = "true";
defparam \WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N16
cycloneive_lcell_comb clear_signal(
	.dataa(gnd),
	.datab(state_8),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam clear_signal.lut_mask = 16'hCC00;
defparam clear_signal.sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N20
cycloneive_lcell_comb \word_counter[0]~7 (
	.dataa(gnd),
	.datab(word_counter[0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\word_counter[0]~7_combout ),
	.cout(\word_counter[0]~8 ));
// synopsys translate_off
defparam \word_counter[0]~7 .lut_mask = 16'h33CC;
defparam \word_counter[0]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N24
cycloneive_lcell_comb \word_counter[2]~11 (
	.dataa(gnd),
	.datab(word_counter[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[1]~10 ),
	.combout(\word_counter[2]~11_combout ),
	.cout(\word_counter[2]~12 ));
// synopsys translate_off
defparam \word_counter[2]~11 .lut_mask = 16'hC30C;
defparam \word_counter[2]~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N4
cycloneive_lcell_comb \word_counter[0]~14 (
	.dataa(state_4),
	.datab(\clear_signal~combout ),
	.datac(state_3),
	.datad(sdr),
	.cin(gnd),
	.combout(\word_counter[0]~14_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[0]~14 .lut_mask = 16'hDCCC;
defparam \word_counter[0]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N25
dffeas \word_counter[2] (
	.clk(TCK),
	.d(\word_counter[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[0]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[0]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[2]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[2] .is_wysiwyg = "true";
defparam \word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N26
cycloneive_lcell_comb \word_counter[3]~15 (
	.dataa(word_counter[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[2]~12 ),
	.combout(\word_counter[3]~15_combout ),
	.cout(\word_counter[3]~16 ));
// synopsys translate_off
defparam \word_counter[3]~15 .lut_mask = 16'h5A5F;
defparam \word_counter[3]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N28
cycloneive_lcell_comb \word_counter[4]~17 (
	.dataa(gnd),
	.datab(word_counter[4]),
	.datac(gnd),
	.datad(gnd),
	.cin(\word_counter[3]~16 ),
	.combout(\word_counter[4]~17_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[4]~17 .lut_mask = 16'hC3C3;
defparam \word_counter[4]~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X43_Y34_N29
dffeas \word_counter[4] (
	.clk(TCK),
	.d(\word_counter[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[0]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[0]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[4]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[4] .is_wysiwyg = "true";
defparam \word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y34_N27
dffeas \word_counter[3] (
	.clk(TCK),
	.d(\word_counter[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[0]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[0]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[3]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[3] .is_wysiwyg = "true";
defparam \word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N30
cycloneive_lcell_comb \word_counter[0]~13 (
	.dataa(word_counter[1]),
	.datab(word_counter[4]),
	.datac(word_counter[3]),
	.datad(word_counter[2]),
	.cin(gnd),
	.combout(\word_counter[0]~13_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[0]~13 .lut_mask = 16'hFBFF;
defparam \word_counter[0]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N2
cycloneive_lcell_comb \word_counter[0]~19 (
	.dataa(virtual_ir_scan_reg),
	.datab(state_8),
	.datac(\word_counter[0]~13_combout ),
	.datad(word_counter[0]),
	.cin(gnd),
	.combout(\word_counter[0]~19_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[0]~19 .lut_mask = 16'h888F;
defparam \word_counter[0]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N21
dffeas \word_counter[0] (
	.clk(TCK),
	.d(\word_counter[0]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[0]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[0]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[0]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[0] .is_wysiwyg = "true";
defparam \word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y34_N0
cycloneive_lcell_comb \WORD_SR~14 (
	.dataa(\WORD_SR~13_combout ),
	.datab(state_4),
	.datac(altera_internal_jtag),
	.datad(word_counter[0]),
	.cin(gnd),
	.combout(\WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~14 .lut_mask = 16'hC0E2;
defparam \WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N18
cycloneive_lcell_comb \WORD_SR~15 (
	.dataa(gnd),
	.datab(state_8),
	.datac(\WORD_SR~14_combout ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\WORD_SR~15_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~15 .lut_mask = 16'h30F0;
defparam \WORD_SR~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N10
cycloneive_lcell_comb \WORD_SR[3]~6 (
	.dataa(state_4),
	.datab(\clear_signal~combout ),
	.datac(state_3),
	.datad(sdr),
	.cin(gnd),
	.combout(\WORD_SR[3]~6_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR[3]~6 .lut_mask = 16'hFECC;
defparam \WORD_SR[3]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N19
dffeas \WORD_SR[3] (
	.clk(TCK),
	.d(\WORD_SR~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[3]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[3]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[3] .is_wysiwyg = "true";
defparam \WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y34_N22
cycloneive_lcell_comb \WORD_SR~10 (
	.dataa(word_counter[1]),
	.datab(word_counter[4]),
	.datac(word_counter[2]),
	.datad(word_counter[0]),
	.cin(gnd),
	.combout(\WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~10 .lut_mask = 16'hEC5C;
defparam \WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y34_N8
cycloneive_lcell_comb \WORD_SR~11 (
	.dataa(\WORD_SR~2_combout ),
	.datab(gnd),
	.datac(\WORD_SR~10_combout ),
	.datad(word_counter[0]),
	.cin(gnd),
	.combout(\WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~11 .lut_mask = 16'hF00A;
defparam \WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N8
cycloneive_lcell_comb \WORD_SR~12 (
	.dataa(state_4),
	.datab(WORD_SR[3]),
	.datac(\WORD_SR~11_combout ),
	.datad(\clear_signal~combout ),
	.cin(gnd),
	.combout(\WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~12 .lut_mask = 16'h00D8;
defparam \WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N9
dffeas \WORD_SR[2] (
	.clk(TCK),
	.d(\WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[3]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[2]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[2] .is_wysiwyg = "true";
defparam \WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N6
cycloneive_lcell_comb \WORD_SR~8 (
	.dataa(\WORD_SR~7_combout ),
	.datab(gnd),
	.datac(word_counter[3]),
	.datad(word_counter[2]),
	.cin(gnd),
	.combout(\WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~8 .lut_mask = 16'h000A;
defparam \WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N14
cycloneive_lcell_comb \WORD_SR~9 (
	.dataa(state_4),
	.datab(\clear_signal~combout ),
	.datac(WORD_SR[2]),
	.datad(\WORD_SR~8_combout ),
	.cin(gnd),
	.combout(\WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~9 .lut_mask = 16'h3320;
defparam \WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y34_N15
dffeas \WORD_SR[1] (
	.clk(TCK),
	.d(\WORD_SR~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[3]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[1]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[1] .is_wysiwyg = "true";
defparam \WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y34_N2
cycloneive_lcell_comb \WORD_SR~3 (
	.dataa(word_counter[1]),
	.datab(word_counter[4]),
	.datac(word_counter[2]),
	.datad(word_counter[0]),
	.cin(gnd),
	.combout(\WORD_SR~3_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~3 .lut_mask = 16'h88AC;
defparam \WORD_SR~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y34_N16
cycloneive_lcell_comb \WORD_SR~4 (
	.dataa(\WORD_SR~2_combout ),
	.datab(\WORD_SR~3_combout ),
	.datac(gnd),
	.datad(word_counter[0]),
	.cin(gnd),
	.combout(\WORD_SR~4_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~4 .lut_mask = 16'hCC88;
defparam \WORD_SR~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y34_N0
cycloneive_lcell_comb \WORD_SR~5 (
	.dataa(state_4),
	.datab(WORD_SR[1]),
	.datac(\WORD_SR~4_combout ),
	.datad(\clear_signal~combout ),
	.cin(gnd),
	.combout(\WORD_SR~5_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~5 .lut_mask = 16'h00D8;
defparam \WORD_SR~5 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule
