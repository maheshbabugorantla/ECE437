// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 64-Bit"
// VERSION "Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"

// DATE "09/18/2017 16:43:29"

// 
// Device: Altera EP4CE115F29C8 Package FBGA780
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module system (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	CLK,
	nRST,
	\syif.halt ,
	\syif.load ,
	\syif.addr ,
	\syif.store ,
	\syif.REN ,
	\syif.WEN ,
	\syif.tbCTRL );
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	CLK;
input 	nRST;
output 	\syif.halt ;
output 	[31:0] \syif.load ;
input 	[31:0] \syif.addr ;
input 	[31:0] \syif.store ;
input 	\syif.REN ;
input 	\syif.WEN ;
input 	\syif.tbCTRL ;

// Design Ports Information
// syif.halt	=>  Location: PIN_T3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[0]	=>  Location: PIN_H16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[1]	=>  Location: PIN_J12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[2]	=>  Location: PIN_AC15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[3]	=>  Location: PIN_R6,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[4]	=>  Location: PIN_U3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[5]	=>  Location: PIN_C13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[6]	=>  Location: PIN_AH17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[7]	=>  Location: PIN_D15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[8]	=>  Location: PIN_A12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[9]	=>  Location: PIN_B11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[10]	=>  Location: PIN_AD11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[11]	=>  Location: PIN_R3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[12]	=>  Location: PIN_AB13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[13]	=>  Location: PIN_AB16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[14]	=>  Location: PIN_AC11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[15]	=>  Location: PIN_B10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[16]	=>  Location: PIN_AB14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[17]	=>  Location: PIN_AF16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[18]	=>  Location: PIN_T22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[19]	=>  Location: PIN_D14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[20]	=>  Location: PIN_P25,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[21]	=>  Location: PIN_AA12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[22]	=>  Location: PIN_H15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[23]	=>  Location: PIN_C16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[24]	=>  Location: PIN_J16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[25]	=>  Location: PIN_C12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[26]	=>  Location: PIN_E15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[27]	=>  Location: PIN_R26,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[28]	=>  Location: PIN_AD14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[29]	=>  Location: PIN_H17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[30]	=>  Location: PIN_AE13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[31]	=>  Location: PIN_M24,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.tbCTRL	=>  Location: PIN_AG15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[1]	=>  Location: PIN_AH15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[0]	=>  Location: PIN_R7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[3]	=>  Location: PIN_G16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[2]	=>  Location: PIN_R4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[5]	=>  Location: PIN_AA13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[4]	=>  Location: PIN_C14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[7]	=>  Location: PIN_R2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[6]	=>  Location: PIN_P26,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[9]	=>  Location: PIN_J17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[8]	=>  Location: PIN_J15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[11]	=>  Location: PIN_R25,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[10]	=>  Location: PIN_B17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[13]	=>  Location: PIN_AE17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[12]	=>  Location: PIN_R1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[15]	=>  Location: PIN_F17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[14]	=>  Location: PIN_P21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[17]	=>  Location: PIN_R23,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[16]	=>  Location: PIN_AB15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[19]	=>  Location: PIN_R22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[18]	=>  Location: PIN_E17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[21]	=>  Location: PIN_A17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[20]	=>  Location: PIN_AE15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[23]	=>  Location: PIN_C15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[22]	=>  Location: PIN_AH12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[25]	=>  Location: PIN_AA16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[24]	=>  Location: PIN_AD15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[27]	=>  Location: PIN_AG18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[26]	=>  Location: PIN_R24,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[29]	=>  Location: PIN_F15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[28]	=>  Location: PIN_D16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[31]	=>  Location: PIN_G18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[30]	=>  Location: PIN_AG19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.WEN	=>  Location: PIN_AF17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.REN	=>  Location: PIN_R21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// nRST	=>  Location: PIN_Y2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// CLK	=>  Location: PIN_J1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[0]	=>  Location: PIN_G14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[1]	=>  Location: PIN_R5,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[2]	=>  Location: PIN_AD12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[3]	=>  Location: PIN_G15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[4]	=>  Location: PIN_A11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[5]	=>  Location: PIN_Y13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[6]	=>  Location: PIN_H14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[7]	=>  Location: PIN_F14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[8]	=>  Location: PIN_AG17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[9]	=>  Location: PIN_Y14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[10]	=>  Location: PIN_D13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[11]	=>  Location: PIN_AG12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[12]	=>  Location: PIN_AB12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[13]	=>  Location: PIN_AA14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[14]	=>  Location: PIN_Y12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[15]	=>  Location: PIN_AF14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[16]	=>  Location: PIN_J14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[17]	=>  Location: PIN_U4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[18]	=>  Location: PIN_J13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[19]	=>  Location: PIN_D12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[20]	=>  Location: PIN_AE16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[21]	=>  Location: PIN_AC12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[22]	=>  Location: PIN_AE14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[23]	=>  Location: PIN_R28,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[24]	=>  Location: PIN_AC14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[25]	=>  Location: PIN_Y15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[26]	=>  Location: PIN_R27,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[27]	=>  Location: PIN_AH19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[28]	=>  Location: PIN_AA15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[29]	=>  Location: PIN_AH18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[30]	=>  Location: PIN_E14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[31]	=>  Location: PIN_AF15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tms	=>  Location: PIN_P8,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tck	=>  Location: PIN_P5,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdi	=>  Location: PIN_P7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdo	=>  Location: PIN_P6,	 I/O Standard: 2.5 V,	 Current Strength: Default


wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ;
wire \CPU|DP|ru_dut|ruif.dmemREN~q ;
wire \CPU|DP|ru_dut|ruif.dmemWEN~q ;
wire \ramaddr~0_combout ;
wire \ramaddr~1_combout ;
wire \ramaddr~2_combout ;
wire \ramaddr~3_combout ;
wire \ramaddr~4_combout ;
wire \ramaddr~5_combout ;
wire \ramaddr~6_combout ;
wire \ramaddr~7_combout ;
wire \ramaddr~8_combout ;
wire \ramaddr~9_combout ;
wire \ramaddr~10_combout ;
wire \ramaddr~11_combout ;
wire \ramaddr~12_combout ;
wire \ramaddr~13_combout ;
wire \ramaddr~14_combout ;
wire \ramaddr~15_combout ;
wire \ramaddr~16_combout ;
wire \ramaddr~17_combout ;
wire \ramaddr~18_combout ;
wire \ramaddr~19_combout ;
wire \ramaddr~20_combout ;
wire \ramaddr~21_combout ;
wire \ramaddr~22_combout ;
wire \ramaddr~23_combout ;
wire \ramaddr~24_combout ;
wire \ramaddr~25_combout ;
wire \ramaddr~26_combout ;
wire \ramaddr~27_combout ;
wire \ramaddr~28_combout ;
wire \ramaddr~29_combout ;
wire \ramaddr~30_combout ;
wire \ramaddr~31_combout ;
wire \ramaddr~32_combout ;
wire \ramaddr~33_combout ;
wire \ramaddr~34_combout ;
wire \ramaddr~35_combout ;
wire \ramaddr~36_combout ;
wire \ramaddr~37_combout ;
wire \ramaddr~38_combout ;
wire \ramaddr~39_combout ;
wire \ramaddr~40_combout ;
wire \ramaddr~41_combout ;
wire \ramaddr~42_combout ;
wire \ramaddr~43_combout ;
wire \ramaddr~44_combout ;
wire \ramaddr~45_combout ;
wire \ramaddr~46_combout ;
wire \ramaddr~47_combout ;
wire \ramaddr~48_combout ;
wire \ramaddr~49_combout ;
wire \ramaddr~50_combout ;
wire \ramaddr~51_combout ;
wire \ramaddr~52_combout ;
wire \ramaddr~53_combout ;
wire \ramaddr~54_combout ;
wire \ramaddr~55_combout ;
wire \ramaddr~56_combout ;
wire \ramaddr~57_combout ;
wire \ramaddr~58_combout ;
wire \ramaddr~59_combout ;
wire \ramaddr~60_combout ;
wire \ramaddr~61_combout ;
wire \ramaddr~62_combout ;
wire \ramaddr~63_combout ;
wire \ramWEN~0_combout ;
wire \ramREN~0_combout ;
wire \RAM|always1~0_combout ;
wire \RAM|ramif.ramload[0]~12_combout ;
wire \RAM|ramif.ramload[1]~13_combout ;
wire \RAM|ramif.ramload[2]~14_combout ;
wire \RAM|ramif.ramload[3]~15_combout ;
wire \RAM|ramif.ramload[4]~16_combout ;
wire \RAM|ramif.ramload[5]~17_combout ;
wire \RAM|ramif.ramload[6]~18_combout ;
wire \RAM|ramif.ramload[7]~19_combout ;
wire \RAM|ramif.ramload[8]~20_combout ;
wire \RAM|ramif.ramload[9]~21_combout ;
wire \RAM|ramif.ramload[10]~22_combout ;
wire \RAM|ramif.ramload[11]~23_combout ;
wire \RAM|ramif.ramload[12]~24_combout ;
wire \RAM|ramif.ramload[13]~25_combout ;
wire \RAM|ramif.ramload[14]~26_combout ;
wire \RAM|ramif.ramload[15]~27_combout ;
wire \RAM|ramif.ramload[16]~28_combout ;
wire \RAM|ramif.ramload[17]~29_combout ;
wire \RAM|ramif.ramload[18]~30_combout ;
wire \RAM|ramif.ramload[19]~31_combout ;
wire \RAM|ramif.ramload[20]~32_combout ;
wire \RAM|ramif.ramload[21]~33_combout ;
wire \RAM|ramif.ramload[22]~34_combout ;
wire \RAM|ramif.ramload[23]~35_combout ;
wire \RAM|ramif.ramload[24]~36_combout ;
wire \RAM|ramif.ramload[25]~37_combout ;
wire \RAM|ramif.ramload[26]~38_combout ;
wire \RAM|ramif.ramload[27]~39_combout ;
wire \RAM|ramif.ramload[28]~40_combout ;
wire \RAM|ramif.ramload[29]~41_combout ;
wire \RAM|ramif.ramload[30]~42_combout ;
wire \RAM|ramif.ramload[31]~43_combout ;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ;
wire \CPUCLK~q ;
wire \CPU|DP|rf_dut|Mux63~9_combout ;
wire \CPU|DP|rf_dut|Mux63~19_combout ;
wire \CPU|DP|cu_dut|cuif.regT[4]~6_combout ;
wire \ramstore~0_combout ;
wire \ramstore~1_combout ;
wire \CPU|DP|rf_dut|Mux32~9_combout ;
wire \CPU|DP|rf_dut|Mux32~19_combout ;
wire \CPU|DP|rf_dut|Mux33~9_combout ;
wire \CPU|DP|rf_dut|Mux33~19_combout ;
wire \CPU|DP|rf_dut|Mux34~9_combout ;
wire \CPU|DP|rf_dut|Mux34~19_combout ;
wire \CPU|DP|rf_dut|Mux35~9_combout ;
wire \CPU|DP|rf_dut|Mux35~19_combout ;
wire \CPU|DP|rf_dut|Mux36~9_combout ;
wire \CPU|DP|rf_dut|Mux36~19_combout ;
wire \CPU|DP|rf_dut|Mux37~9_combout ;
wire \CPU|DP|rf_dut|Mux37~19_combout ;
wire \CPU|DP|rf_dut|Mux38~9_combout ;
wire \CPU|DP|rf_dut|Mux38~19_combout ;
wire \CPU|DP|rf_dut|Mux39~9_combout ;
wire \CPU|DP|rf_dut|Mux39~19_combout ;
wire \CPU|DP|rf_dut|Mux40~9_combout ;
wire \CPU|DP|rf_dut|Mux40~19_combout ;
wire \CPU|DP|rf_dut|Mux41~9_combout ;
wire \CPU|DP|rf_dut|Mux41~19_combout ;
wire \CPU|DP|rf_dut|Mux42~9_combout ;
wire \CPU|DP|rf_dut|Mux42~19_combout ;
wire \CPU|DP|rf_dut|Mux43~9_combout ;
wire \CPU|DP|rf_dut|Mux43~19_combout ;
wire \CPU|DP|rf_dut|Mux58~9_combout ;
wire \CPU|DP|rf_dut|Mux58~19_combout ;
wire \CPU|DP|rf_dut|Mux44~9_combout ;
wire \CPU|DP|rf_dut|Mux44~19_combout ;
wire \CPU|DP|rf_dut|Mux45~9_combout ;
wire \CPU|DP|rf_dut|Mux45~19_combout ;
wire \CPU|DP|rf_dut|Mux46~9_combout ;
wire \CPU|DP|rf_dut|Mux46~19_combout ;
wire \CPU|DP|rf_dut|Mux47~9_combout ;
wire \CPU|DP|rf_dut|Mux47~19_combout ;
wire \CPU|DP|rf_dut|Mux48~9_combout ;
wire \CPU|DP|rf_dut|Mux48~19_combout ;
wire \CPU|DP|rf_dut|Mux49~9_combout ;
wire \CPU|DP|rf_dut|Mux49~19_combout ;
wire \CPU|DP|rf_dut|Mux50~9_combout ;
wire \CPU|DP|rf_dut|Mux50~19_combout ;
wire \CPU|DP|rf_dut|Mux51~9_combout ;
wire \CPU|DP|rf_dut|Mux51~19_combout ;
wire \CPU|DP|rf_dut|Mux52~9_combout ;
wire \CPU|DP|rf_dut|Mux52~19_combout ;
wire \CPU|DP|rf_dut|Mux53~9_combout ;
wire \CPU|DP|rf_dut|Mux53~19_combout ;
wire \CPU|DP|rf_dut|Mux54~9_combout ;
wire \CPU|DP|rf_dut|Mux54~19_combout ;
wire \CPU|DP|rf_dut|Mux55~9_combout ;
wire \CPU|DP|rf_dut|Mux55~19_combout ;
wire \CPU|DP|rf_dut|Mux56~9_combout ;
wire \CPU|DP|rf_dut|Mux56~19_combout ;
wire \CPU|DP|rf_dut|Mux57~9_combout ;
wire \CPU|DP|rf_dut|Mux57~19_combout ;
wire \CPU|DP|rf_dut|Mux62~9_combout ;
wire \CPU|DP|rf_dut|Mux62~19_combout ;
wire \CPU|DP|rf_dut|Mux61~9_combout ;
wire \CPU|DP|rf_dut|Mux61~19_combout ;
wire \CPU|DP|rf_dut|Mux60~9_combout ;
wire \CPU|DP|rf_dut|Mux60~19_combout ;
wire \CPU|DP|rf_dut|Mux59~9_combout ;
wire \CPU|DP|rf_dut|Mux59~19_combout ;
wire \ramstore~2_combout ;
wire \ramstore~3_combout ;
wire \ramstore~4_combout ;
wire \ramstore~5_combout ;
wire \ramstore~6_combout ;
wire \ramstore~7_combout ;
wire \ramstore~8_combout ;
wire \ramstore~9_combout ;
wire \ramstore~10_combout ;
wire \ramstore~11_combout ;
wire \ramstore~12_combout ;
wire \ramstore~13_combout ;
wire \ramstore~14_combout ;
wire \ramstore~15_combout ;
wire \ramstore~16_combout ;
wire \ramstore~17_combout ;
wire \ramstore~18_combout ;
wire \ramstore~19_combout ;
wire \ramstore~20_combout ;
wire \ramstore~21_combout ;
wire \ramstore~22_combout ;
wire \ramstore~23_combout ;
wire \ramstore~24_combout ;
wire \ramstore~25_combout ;
wire \ramstore~26_combout ;
wire \ramstore~27_combout ;
wire \ramstore~28_combout ;
wire \ramstore~29_combout ;
wire \ramstore~30_combout ;
wire \ramstore~31_combout ;
wire \ramstore~32_combout ;
wire \ramstore~33_combout ;
wire \ramstore~34_combout ;
wire \ramstore~35_combout ;
wire \ramstore~36_combout ;
wire \ramstore~37_combout ;
wire \ramstore~38_combout ;
wire \ramstore~39_combout ;
wire \ramstore~40_combout ;
wire \ramstore~41_combout ;
wire \ramstore~42_combout ;
wire \ramstore~43_combout ;
wire \ramstore~44_combout ;
wire \ramstore~45_combout ;
wire \ramstore~46_combout ;
wire \ramstore~47_combout ;
wire \ramstore~48_combout ;
wire \ramstore~49_combout ;
wire \ramstore~50_combout ;
wire \ramstore~51_combout ;
wire \ramstore~52_combout ;
wire \ramstore~53_combout ;
wire \ramstore~54_combout ;
wire \ramstore~55_combout ;
wire \ramstore~56_combout ;
wire \ramstore~57_combout ;
wire \ramstore~58_combout ;
wire \ramstore~59_combout ;
wire \ramstore~60_combout ;
wire \ramstore~61_combout ;
wire \ramstore~62_combout ;
wire \ramstore~63_combout ;
wire \Equal0~0_combout ;
wire \CPUCLK~0_combout ;
wire \count[3]~0_combout ;
wire \count[2]~1_combout ;
wire \count[1]~2_combout ;
wire \count~3_combout ;
wire \RAM|ramif.ramload[26]~44_combout ;
wire \RAM|ramif.ramload[27]~45_combout ;
wire \RAM|ramif.ramload[28]~46_combout ;
wire \RAM|ramif.ramload[29]~47_combout ;
wire \RAM|ramif.ramload[30]~48_combout ;
wire \RAM|ramif.ramload[31]~49_combout ;
wire \ramaddr~29_wirecell_combout ;
wire \altera_internal_jtag~TCKUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ;
wire \syif.tbCTRL~input_o ;
wire \syif.addr[1]~input_o ;
wire \syif.addr[0]~input_o ;
wire \syif.addr[3]~input_o ;
wire \syif.addr[2]~input_o ;
wire \syif.addr[5]~input_o ;
wire \syif.addr[4]~input_o ;
wire \syif.addr[7]~input_o ;
wire \syif.addr[6]~input_o ;
wire \syif.addr[9]~input_o ;
wire \syif.addr[8]~input_o ;
wire \syif.addr[11]~input_o ;
wire \syif.addr[10]~input_o ;
wire \syif.addr[13]~input_o ;
wire \syif.addr[12]~input_o ;
wire \syif.addr[15]~input_o ;
wire \syif.addr[14]~input_o ;
wire \syif.addr[17]~input_o ;
wire \syif.addr[16]~input_o ;
wire \syif.addr[19]~input_o ;
wire \syif.addr[18]~input_o ;
wire \syif.addr[21]~input_o ;
wire \syif.addr[20]~input_o ;
wire \syif.addr[23]~input_o ;
wire \syif.addr[22]~input_o ;
wire \syif.addr[25]~input_o ;
wire \syif.addr[24]~input_o ;
wire \syif.addr[27]~input_o ;
wire \syif.addr[26]~input_o ;
wire \syif.addr[29]~input_o ;
wire \syif.addr[28]~input_o ;
wire \syif.addr[31]~input_o ;
wire \syif.addr[30]~input_o ;
wire \syif.WEN~input_o ;
wire \syif.REN~input_o ;
wire \nRST~input_o ;
wire \CLK~input_o ;
wire \syif.store[0]~input_o ;
wire \syif.store[1]~input_o ;
wire \syif.store[2]~input_o ;
wire \syif.store[3]~input_o ;
wire \syif.store[4]~input_o ;
wire \syif.store[5]~input_o ;
wire \syif.store[6]~input_o ;
wire \syif.store[7]~input_o ;
wire \syif.store[8]~input_o ;
wire \syif.store[9]~input_o ;
wire \syif.store[10]~input_o ;
wire \syif.store[11]~input_o ;
wire \syif.store[12]~input_o ;
wire \syif.store[13]~input_o ;
wire \syif.store[14]~input_o ;
wire \syif.store[15]~input_o ;
wire \syif.store[16]~input_o ;
wire \syif.store[17]~input_o ;
wire \syif.store[18]~input_o ;
wire \syif.store[19]~input_o ;
wire \syif.store[20]~input_o ;
wire \syif.store[21]~input_o ;
wire \syif.store[22]~input_o ;
wire \syif.store[23]~input_o ;
wire \syif.store[24]~input_o ;
wire \syif.store[25]~input_o ;
wire \syif.store[26]~input_o ;
wire \syif.store[27]~input_o ;
wire \syif.store[28]~input_o ;
wire \syif.store[29]~input_o ;
wire \syif.store[30]~input_o ;
wire \syif.store[31]~input_o ;
wire \altera_internal_jtag~TCKUTAPclkctrl_outclk ;
wire \CPUCLK~clkctrl_outclk ;
wire \nRST~inputclkctrl_outclk ;
wire \CLK~inputclkctrl_outclk ;
wire \CPU|DP|dpif.halt~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ;
wire \~QIC_CREATED_GND~I_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~14 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~8 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~12 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ;
wire \altera_internal_jtag~TDO ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg ;
wire [9:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg ;
wire [5:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt ;
wire [15:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR ;
wire [3:0] count;
wire [31:0] \CPU|DP|pc_dut|pcif.imemaddr ;
wire [31:0] \CPU|CM|daddr ;
wire [3:0] \RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg ;


ram RAM(
	.is_in_use_reg(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.ramaddr(\ramaddr~1_combout ),
	.ramaddr1(\ramaddr~3_combout ),
	.ramaddr2(\ramaddr~5_combout ),
	.ramaddr3(\ramaddr~7_combout ),
	.ramaddr4(\ramaddr~9_combout ),
	.ramaddr5(\ramaddr~11_combout ),
	.ramaddr6(\ramaddr~13_combout ),
	.ramaddr7(\ramaddr~15_combout ),
	.ramaddr8(\ramaddr~17_combout ),
	.ramaddr9(\ramaddr~19_combout ),
	.ramaddr10(\ramaddr~21_combout ),
	.ramaddr11(\ramaddr~23_combout ),
	.ramaddr12(\ramaddr~25_combout ),
	.ramaddr13(\ramaddr~27_combout ),
	.ramaddr14(\ramaddr~29_combout ),
	.ramaddr15(\ramaddr~31_combout ),
	.\ramif.ramaddr ({gnd,gnd,gnd,gnd,gnd,gnd,\ramaddr~49_combout ,gnd,gnd,gnd,\ramaddr~41_combout ,gnd,\ramaddr~37_combout ,gnd,\ramaddr~33_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.ramaddr16(\ramaddr~35_combout ),
	.ramaddr17(\ramaddr~39_combout ),
	.ramaddr18(\ramaddr~43_combout ),
	.ramaddr19(\ramaddr~45_combout ),
	.ramaddr20(\ramaddr~47_combout ),
	.ramaddr21(\ramaddr~51_combout ),
	.ramaddr22(\ramaddr~53_combout ),
	.ramaddr23(\ramaddr~55_combout ),
	.ramaddr24(\ramaddr~57_combout ),
	.ramaddr25(\ramaddr~59_combout ),
	.ramaddr26(\ramaddr~61_combout ),
	.ramaddr27(\ramaddr~63_combout ),
	.ramWEN(\ramWEN~0_combout ),
	.ramREN(\ramREN~0_combout ),
	.always1(\RAM|always1~0_combout ),
	.ramiframload_0(\RAM|ramif.ramload[0]~12_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~13_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~14_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~15_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~16_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~17_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~18_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~19_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~20_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~21_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~22_combout ),
	.ramiframload_11(\RAM|ramif.ramload[11]~23_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~24_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~25_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~26_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~27_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~28_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~29_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~30_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~31_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~32_combout ),
	.ramiframload_21(\RAM|ramif.ramload[21]~33_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~34_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~35_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~36_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~37_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~38_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~39_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~40_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~41_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~42_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~43_combout ),
	.ir_loaded_address_reg_0(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.ir_loaded_address_reg_1(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.ir_loaded_address_reg_2(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.ir_loaded_address_reg_3(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.tdo(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.ramstore(\ramstore~1_combout ),
	.ramstore1(\ramstore~3_combout ),
	.ramstore2(\ramstore~5_combout ),
	.ramstore3(\ramstore~7_combout ),
	.ramstore4(\ramstore~9_combout ),
	.ramstore5(\ramstore~11_combout ),
	.ramstore6(\ramstore~13_combout ),
	.ramstore7(\ramstore~15_combout ),
	.ramstore8(\ramstore~17_combout ),
	.ramstore9(\ramstore~19_combout ),
	.ramstore10(\ramstore~21_combout ),
	.ramstore11(\ramstore~23_combout ),
	.ramstore12(\ramstore~25_combout ),
	.ramstore13(\ramstore~27_combout ),
	.ramstore14(\ramstore~29_combout ),
	.ramstore15(\ramstore~31_combout ),
	.ramstore16(\ramstore~33_combout ),
	.ramstore17(\ramstore~35_combout ),
	.ramstore18(\ramstore~37_combout ),
	.ramstore19(\ramstore~39_combout ),
	.ramstore20(\ramstore~41_combout ),
	.ramstore21(\ramstore~43_combout ),
	.ramstore22(\ramstore~45_combout ),
	.ramstore23(\ramstore~47_combout ),
	.ramstore24(\ramstore~49_combout ),
	.ramstore25(\ramstore~51_combout ),
	.ramstore26(\ramstore~53_combout ),
	.ramstore27(\ramstore~55_combout ),
	.ramstore28(\ramstore~57_combout ),
	.ramstore29(\ramstore~59_combout ),
	.ramstore30(\ramstore~61_combout ),
	.ramstore31(\ramstore~63_combout ),
	.ramiframload_261(\RAM|ramif.ramload[26]~44_combout ),
	.ramiframload_271(\RAM|ramif.ramload[27]~45_combout ),
	.ramiframload_281(\RAM|ramif.ramload[28]~46_combout ),
	.ramiframload_291(\RAM|ramif.ramload[29]~47_combout ),
	.ramiframload_301(\RAM|ramif.ramload[30]~48_combout ),
	.ramiframload_311(\RAM|ramif.ramload[31]~49_combout ),
	.ramaddr28(\ramaddr~29_wirecell_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.irf_reg_0_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.irf_reg_1_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.irf_reg_2_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.irf_reg_3_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.irf_reg_4_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.node_ena_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.clr_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.virtual_ir_scan_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.state_5(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.state_8(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.nRST(\nRST~input_o ),
	.altera_internal_jtag1(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.nRST1(\nRST~inputclkctrl_outclk ),
	.CLK(\CLK~inputclkctrl_outclk ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

singlecycle CPU(
	.pcifimemaddr_29(\CPU|DP|pc_dut|pcif.imemaddr [29]),
	.pcifimemaddr_28(\CPU|DP|pc_dut|pcif.imemaddr [28]),
	.pcifimemaddr_31(\CPU|DP|pc_dut|pcif.imemaddr [31]),
	.pcifimemaddr_30(\CPU|DP|pc_dut|pcif.imemaddr [30]),
	.daddr_1(\CPU|CM|daddr [1]),
	.pcifimemaddr_1(\CPU|DP|pc_dut|pcif.imemaddr [1]),
	.ruifdmemREN(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.ruifdmemWEN(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.daddr_0(\CPU|CM|daddr [0]),
	.pcifimemaddr_0(\CPU|DP|pc_dut|pcif.imemaddr [0]),
	.daddr_3(\CPU|CM|daddr [3]),
	.pcifimemaddr_3(\CPU|DP|pc_dut|pcif.imemaddr [3]),
	.daddr_2(\CPU|CM|daddr [2]),
	.pcifimemaddr_2(\CPU|DP|pc_dut|pcif.imemaddr [2]),
	.daddr_5(\CPU|CM|daddr [5]),
	.pcifimemaddr_5(\CPU|DP|pc_dut|pcif.imemaddr [5]),
	.daddr_4(\CPU|CM|daddr [4]),
	.pcifimemaddr_4(\CPU|DP|pc_dut|pcif.imemaddr [4]),
	.daddr_7(\CPU|CM|daddr [7]),
	.pcifimemaddr_7(\CPU|DP|pc_dut|pcif.imemaddr [7]),
	.daddr_6(\CPU|CM|daddr [6]),
	.pcifimemaddr_6(\CPU|DP|pc_dut|pcif.imemaddr [6]),
	.daddr_9(\CPU|CM|daddr [9]),
	.pcifimemaddr_9(\CPU|DP|pc_dut|pcif.imemaddr [9]),
	.pcifimemaddr_8(\CPU|DP|pc_dut|pcif.imemaddr [8]),
	.daddr_8(\CPU|CM|daddr [8]),
	.daddr_11(\CPU|CM|daddr [11]),
	.pcifimemaddr_11(\CPU|DP|pc_dut|pcif.imemaddr [11]),
	.pcifimemaddr_10(\CPU|DP|pc_dut|pcif.imemaddr [10]),
	.daddr_10(\CPU|CM|daddr [10]),
	.daddr_13(\CPU|CM|daddr [13]),
	.pcifimemaddr_13(\CPU|DP|pc_dut|pcif.imemaddr [13]),
	.daddr_12(\CPU|CM|daddr [12]),
	.pcifimemaddr_12(\CPU|DP|pc_dut|pcif.imemaddr [12]),
	.daddr_15(\CPU|CM|daddr [15]),
	.pcifimemaddr_15(\CPU|DP|pc_dut|pcif.imemaddr [15]),
	.daddr_14(\CPU|CM|daddr [14]),
	.pcifimemaddr_14(\CPU|DP|pc_dut|pcif.imemaddr [14]),
	.daddr_17(\CPU|CM|daddr [17]),
	.pcifimemaddr_17(\CPU|DP|pc_dut|pcif.imemaddr [17]),
	.pcifimemaddr_16(\CPU|DP|pc_dut|pcif.imemaddr [16]),
	.daddr_16(\CPU|CM|daddr [16]),
	.daddr_19(\CPU|CM|daddr [19]),
	.pcifimemaddr_19(\CPU|DP|pc_dut|pcif.imemaddr [19]),
	.daddr_18(\CPU|CM|daddr [18]),
	.pcifimemaddr_18(\CPU|DP|pc_dut|pcif.imemaddr [18]),
	.daddr_21(\CPU|CM|daddr [21]),
	.pcifimemaddr_21(\CPU|DP|pc_dut|pcif.imemaddr [21]),
	.daddr_20(\CPU|CM|daddr [20]),
	.pcifimemaddr_20(\CPU|DP|pc_dut|pcif.imemaddr [20]),
	.daddr_23(\CPU|CM|daddr [23]),
	.pcifimemaddr_23(\CPU|DP|pc_dut|pcif.imemaddr [23]),
	.daddr_22(\CPU|CM|daddr [22]),
	.pcifimemaddr_22(\CPU|DP|pc_dut|pcif.imemaddr [22]),
	.daddr_25(\CPU|CM|daddr [25]),
	.pcifimemaddr_25(\CPU|DP|pc_dut|pcif.imemaddr [25]),
	.daddr_24(\CPU|CM|daddr [24]),
	.pcifimemaddr_24(\CPU|DP|pc_dut|pcif.imemaddr [24]),
	.daddr_27(\CPU|CM|daddr [27]),
	.pcifimemaddr_27(\CPU|DP|pc_dut|pcif.imemaddr [27]),
	.daddr_26(\CPU|CM|daddr [26]),
	.pcifimemaddr_26(\CPU|DP|pc_dut|pcif.imemaddr [26]),
	.daddr_29(\CPU|CM|daddr [29]),
	.daddr_28(\CPU|CM|daddr [28]),
	.daddr_31(\CPU|CM|daddr [31]),
	.daddr_30(\CPU|CM|daddr [30]),
	.always1(\RAM|always1~0_combout ),
	.ramiframload_0(\RAM|ramif.ramload[0]~12_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~13_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~14_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~15_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~16_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~17_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~18_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~19_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~20_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~21_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~22_combout ),
	.ramiframload_11(\RAM|ramif.ramload[11]~23_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~24_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~25_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~26_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~27_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~28_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~29_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~30_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~31_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~32_combout ),
	.ramiframload_21(\RAM|ramif.ramload[21]~33_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~34_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~35_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~36_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~37_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~38_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~39_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~40_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~41_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~42_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~43_combout ),
	.Mux63(\CPU|DP|rf_dut|Mux63~9_combout ),
	.Mux631(\CPU|DP|rf_dut|Mux63~19_combout ),
	.cuifregT_4(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.Mux32(\CPU|DP|rf_dut|Mux32~9_combout ),
	.Mux321(\CPU|DP|rf_dut|Mux32~19_combout ),
	.Mux33(\CPU|DP|rf_dut|Mux33~9_combout ),
	.Mux331(\CPU|DP|rf_dut|Mux33~19_combout ),
	.Mux34(\CPU|DP|rf_dut|Mux34~9_combout ),
	.Mux341(\CPU|DP|rf_dut|Mux34~19_combout ),
	.Mux35(\CPU|DP|rf_dut|Mux35~9_combout ),
	.Mux351(\CPU|DP|rf_dut|Mux35~19_combout ),
	.Mux36(\CPU|DP|rf_dut|Mux36~9_combout ),
	.Mux361(\CPU|DP|rf_dut|Mux36~19_combout ),
	.Mux37(\CPU|DP|rf_dut|Mux37~9_combout ),
	.Mux371(\CPU|DP|rf_dut|Mux37~19_combout ),
	.Mux38(\CPU|DP|rf_dut|Mux38~9_combout ),
	.Mux381(\CPU|DP|rf_dut|Mux38~19_combout ),
	.Mux39(\CPU|DP|rf_dut|Mux39~9_combout ),
	.Mux391(\CPU|DP|rf_dut|Mux39~19_combout ),
	.Mux40(\CPU|DP|rf_dut|Mux40~9_combout ),
	.Mux401(\CPU|DP|rf_dut|Mux40~19_combout ),
	.Mux41(\CPU|DP|rf_dut|Mux41~9_combout ),
	.Mux411(\CPU|DP|rf_dut|Mux41~19_combout ),
	.Mux42(\CPU|DP|rf_dut|Mux42~9_combout ),
	.Mux421(\CPU|DP|rf_dut|Mux42~19_combout ),
	.Mux43(\CPU|DP|rf_dut|Mux43~9_combout ),
	.Mux431(\CPU|DP|rf_dut|Mux43~19_combout ),
	.Mux58(\CPU|DP|rf_dut|Mux58~9_combout ),
	.Mux581(\CPU|DP|rf_dut|Mux58~19_combout ),
	.Mux44(\CPU|DP|rf_dut|Mux44~9_combout ),
	.Mux441(\CPU|DP|rf_dut|Mux44~19_combout ),
	.Mux45(\CPU|DP|rf_dut|Mux45~9_combout ),
	.Mux451(\CPU|DP|rf_dut|Mux45~19_combout ),
	.Mux46(\CPU|DP|rf_dut|Mux46~9_combout ),
	.Mux461(\CPU|DP|rf_dut|Mux46~19_combout ),
	.Mux47(\CPU|DP|rf_dut|Mux47~9_combout ),
	.Mux471(\CPU|DP|rf_dut|Mux47~19_combout ),
	.Mux48(\CPU|DP|rf_dut|Mux48~9_combout ),
	.Mux481(\CPU|DP|rf_dut|Mux48~19_combout ),
	.Mux49(\CPU|DP|rf_dut|Mux49~9_combout ),
	.Mux491(\CPU|DP|rf_dut|Mux49~19_combout ),
	.Mux50(\CPU|DP|rf_dut|Mux50~9_combout ),
	.Mux501(\CPU|DP|rf_dut|Mux50~19_combout ),
	.Mux51(\CPU|DP|rf_dut|Mux51~9_combout ),
	.Mux511(\CPU|DP|rf_dut|Mux51~19_combout ),
	.Mux52(\CPU|DP|rf_dut|Mux52~9_combout ),
	.Mux521(\CPU|DP|rf_dut|Mux52~19_combout ),
	.Mux53(\CPU|DP|rf_dut|Mux53~9_combout ),
	.Mux531(\CPU|DP|rf_dut|Mux53~19_combout ),
	.Mux54(\CPU|DP|rf_dut|Mux54~9_combout ),
	.Mux541(\CPU|DP|rf_dut|Mux54~19_combout ),
	.Mux55(\CPU|DP|rf_dut|Mux55~9_combout ),
	.Mux551(\CPU|DP|rf_dut|Mux55~19_combout ),
	.Mux56(\CPU|DP|rf_dut|Mux56~9_combout ),
	.Mux561(\CPU|DP|rf_dut|Mux56~19_combout ),
	.Mux57(\CPU|DP|rf_dut|Mux57~9_combout ),
	.Mux571(\CPU|DP|rf_dut|Mux57~19_combout ),
	.Mux62(\CPU|DP|rf_dut|Mux62~9_combout ),
	.Mux621(\CPU|DP|rf_dut|Mux62~19_combout ),
	.Mux61(\CPU|DP|rf_dut|Mux61~9_combout ),
	.Mux611(\CPU|DP|rf_dut|Mux61~19_combout ),
	.Mux60(\CPU|DP|rf_dut|Mux60~9_combout ),
	.Mux601(\CPU|DP|rf_dut|Mux60~19_combout ),
	.Mux59(\CPU|DP|rf_dut|Mux59~9_combout ),
	.Mux591(\CPU|DP|rf_dut|Mux59~19_combout ),
	.ramiframload_261(\RAM|ramif.ramload[26]~44_combout ),
	.ramiframload_271(\RAM|ramif.ramload[27]~45_combout ),
	.ramiframload_281(\RAM|ramif.ramload[28]~46_combout ),
	.ramiframload_291(\RAM|ramif.ramload[29]~47_combout ),
	.ramiframload_301(\RAM|ramif.ramload[30]~48_combout ),
	.ramiframload_311(\RAM|ramif.ramload[31]~49_combout ),
	.nRST(\nRST~input_o ),
	.CLK(\CPUCLK~clkctrl_outclk ),
	.nRST1(\nRST~inputclkctrl_outclk ),
	.dpifhalt(\CPU|DP|dpif.halt~q ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X55_Y36_N6
cycloneive_lcell_comb \ramaddr~0 (
// Equation(s):
// \ramaddr~0_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[1]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdmemREN) # (ruifdmemWEN))))

	.dataa(\syif.addr[1]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datad(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~0 .lut_mask = 16'hBBB8;
defparam \ramaddr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N20
cycloneive_lcell_comb \ramaddr~1 (
// Equation(s):
// \ramaddr~1_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~0_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~0_combout  & (daddr_1)) # (!\ramaddr~0_combout  & ((pcifimemaddr_1)))))

	.dataa(\CPU|CM|daddr [1]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|pc_dut|pcif.imemaddr [1]),
	.datad(\ramaddr~0_combout ),
	.cin(gnd),
	.combout(\ramaddr~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~1 .lut_mask = 16'hEE30;
defparam \ramaddr~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N0
cycloneive_lcell_comb \ramaddr~2 (
// Equation(s):
// \ramaddr~2_combout  = (ruifdmemREN & (daddr_0)) # (!ruifdmemREN & ((ruifdmemWEN & (daddr_0)) # (!ruifdmemWEN & ((pcifimemaddr_0)))))

	.dataa(\CPU|CM|daddr [0]),
	.datab(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datac(\CPU|DP|pc_dut|pcif.imemaddr [0]),
	.datad(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~2 .lut_mask = 16'hAAB8;
defparam \ramaddr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N2
cycloneive_lcell_comb \ramaddr~3 (
// Equation(s):
// \ramaddr~3_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[0]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~2_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[0]~input_o ),
	.datad(\ramaddr~2_combout ),
	.cin(gnd),
	.combout(\ramaddr~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~3 .lut_mask = 16'hF3C0;
defparam \ramaddr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N6
cycloneive_lcell_comb \ramaddr~4 (
// Equation(s):
// \ramaddr~4_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[3]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdmemREN) # (ruifdmemWEN))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[3]~input_o ),
	.datac(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datad(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~4 .lut_mask = 16'hDDD8;
defparam \ramaddr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N2
cycloneive_lcell_comb \ramaddr~5 (
// Equation(s):
// \ramaddr~5_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~4_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~4_combout  & ((daddr_3))) # (!\ramaddr~4_combout  & (pcifimemaddr_3))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|pc_dut|pcif.imemaddr [3]),
	.datac(\CPU|CM|daddr [3]),
	.datad(\ramaddr~4_combout ),
	.cin(gnd),
	.combout(\ramaddr~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~5 .lut_mask = 16'hFA44;
defparam \ramaddr~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N18
cycloneive_lcell_comb \ramaddr~6 (
// Equation(s):
// \ramaddr~6_combout  = (ruifdmemREN & (daddr_2)) # (!ruifdmemREN & ((ruifdmemWEN & (daddr_2)) # (!ruifdmemWEN & ((pcifimemaddr_2)))))

	.dataa(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datab(\CPU|CM|daddr [2]),
	.datac(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datad(\CPU|DP|pc_dut|pcif.imemaddr [2]),
	.cin(gnd),
	.combout(\ramaddr~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~6 .lut_mask = 16'hCDC8;
defparam \ramaddr~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N0
cycloneive_lcell_comb \ramaddr~7 (
// Equation(s):
// \ramaddr~7_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[2]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~6_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[2]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~6_combout ),
	.cin(gnd),
	.combout(\ramaddr~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~7 .lut_mask = 16'hDD88;
defparam \ramaddr~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N18
cycloneive_lcell_comb \ramaddr~8 (
// Equation(s):
// \ramaddr~8_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[5]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdmemWEN) # (ruifdmemREN))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[5]~input_o ),
	.datac(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datad(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~8 .lut_mask = 16'hDDD8;
defparam \ramaddr~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N6
cycloneive_lcell_comb \ramaddr~9 (
// Equation(s):
// \ramaddr~9_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~8_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~8_combout  & (daddr_5)) # (!\ramaddr~8_combout  & ((pcifimemaddr_5)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [5]),
	.datac(\CPU|DP|pc_dut|pcif.imemaddr [5]),
	.datad(\ramaddr~8_combout ),
	.cin(gnd),
	.combout(\ramaddr~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~9 .lut_mask = 16'hEE50;
defparam \ramaddr~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N2
cycloneive_lcell_comb \ramaddr~10 (
// Equation(s):
// \ramaddr~10_combout  = (ruifdmemWEN & (((daddr_4)))) # (!ruifdmemWEN & ((ruifdmemREN & ((daddr_4))) # (!ruifdmemREN & (pcifimemaddr_4))))

	.dataa(\CPU|DP|pc_dut|pcif.imemaddr [4]),
	.datab(\CPU|CM|daddr [4]),
	.datac(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datad(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~10 .lut_mask = 16'hCCCA;
defparam \ramaddr~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N16
cycloneive_lcell_comb \ramaddr~11 (
// Equation(s):
// \ramaddr~11_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[4]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~10_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[4]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~10_combout ),
	.cin(gnd),
	.combout(\ramaddr~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~11 .lut_mask = 16'hDD88;
defparam \ramaddr~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N16
cycloneive_lcell_comb \ramaddr~12 (
// Equation(s):
// \ramaddr~12_combout  = (ruifdmemWEN & (((daddr_7)))) # (!ruifdmemWEN & ((ruifdmemREN & ((daddr_7))) # (!ruifdmemREN & (pcifimemaddr_7))))

	.dataa(\CPU|DP|pc_dut|pcif.imemaddr [7]),
	.datab(\CPU|CM|daddr [7]),
	.datac(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datad(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~12 .lut_mask = 16'hCCCA;
defparam \ramaddr~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N28
cycloneive_lcell_comb \ramaddr~13 (
// Equation(s):
// \ramaddr~13_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[7]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~12_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[7]~input_o ),
	.datad(\ramaddr~12_combout ),
	.cin(gnd),
	.combout(\ramaddr~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~13 .lut_mask = 16'hF3C0;
defparam \ramaddr~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N0
cycloneive_lcell_comb \ramaddr~14 (
// Equation(s):
// \ramaddr~14_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[6]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdmemREN) # (ruifdmemWEN))))

	.dataa(\syif.addr[6]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datad(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~14 .lut_mask = 16'hBBB8;
defparam \ramaddr~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N14
cycloneive_lcell_comb \ramaddr~15 (
// Equation(s):
// \ramaddr~15_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~14_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~14_combout  & (daddr_6)) # (!\ramaddr~14_combout  & ((pcifimemaddr_6)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [6]),
	.datac(\CPU|DP|pc_dut|pcif.imemaddr [6]),
	.datad(\ramaddr~14_combout ),
	.cin(gnd),
	.combout(\ramaddr~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~15 .lut_mask = 16'hEE50;
defparam \ramaddr~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N6
cycloneive_lcell_comb \ramaddr~16 (
// Equation(s):
// \ramaddr~16_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[9]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdmemWEN) # (ruifdmemREN))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[9]~input_o ),
	.datac(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datad(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~16 .lut_mask = 16'hDDD8;
defparam \ramaddr~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N14
cycloneive_lcell_comb \ramaddr~17 (
// Equation(s):
// \ramaddr~17_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~16_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~16_combout  & (daddr_9)) # (!\ramaddr~16_combout  & ((pcifimemaddr_9)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [9]),
	.datac(\CPU|DP|pc_dut|pcif.imemaddr [9]),
	.datad(\ramaddr~16_combout ),
	.cin(gnd),
	.combout(\ramaddr~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~17 .lut_mask = 16'hEE50;
defparam \ramaddr~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N10
cycloneive_lcell_comb \ramaddr~18 (
// Equation(s):
// \ramaddr~18_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[8]~input_o )) # (!\syif.tbCTRL~input_o  & (((!ruifdmemWEN & !ruifdmemREN))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[8]~input_o ),
	.datac(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datad(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~18 .lut_mask = 16'h888D;
defparam \ramaddr~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N12
cycloneive_lcell_comb \ramaddr~19 (
// Equation(s):
// \ramaddr~19_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~18_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~18_combout  & (pcifimemaddr_8)) # (!\ramaddr~18_combout  & ((daddr_8)))))

	.dataa(\CPU|DP|pc_dut|pcif.imemaddr [8]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|CM|daddr [8]),
	.datad(\ramaddr~18_combout ),
	.cin(gnd),
	.combout(\ramaddr~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~19 .lut_mask = 16'hEE30;
defparam \ramaddr~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N6
cycloneive_lcell_comb \ramaddr~20 (
// Equation(s):
// \ramaddr~20_combout  = (ruifdmemREN & (daddr_11)) # (!ruifdmemREN & ((ruifdmemWEN & (daddr_11)) # (!ruifdmemWEN & ((pcifimemaddr_11)))))

	.dataa(\CPU|CM|daddr [11]),
	.datab(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datac(\CPU|DP|pc_dut|pcif.imemaddr [11]),
	.datad(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~20 .lut_mask = 16'hAAB8;
defparam \ramaddr~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N30
cycloneive_lcell_comb \ramaddr~21 (
// Equation(s):
// \ramaddr~21_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[11]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~20_combout )))

	.dataa(\syif.addr[11]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~20_combout ),
	.cin(gnd),
	.combout(\ramaddr~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~21 .lut_mask = 16'hAFA0;
defparam \ramaddr~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N14
cycloneive_lcell_comb \ramaddr~22 (
// Equation(s):
// \ramaddr~22_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[10]~input_o )) # (!\syif.tbCTRL~input_o  & (((!ruifdmemREN & !ruifdmemWEN))))

	.dataa(\syif.addr[10]~input_o ),
	.datab(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~22 .lut_mask = 16'hA0A3;
defparam \ramaddr~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N28
cycloneive_lcell_comb \ramaddr~23 (
// Equation(s):
// \ramaddr~23_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~22_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~22_combout  & (pcifimemaddr_10)) # (!\ramaddr~22_combout  & ((daddr_10)))))

	.dataa(\CPU|DP|pc_dut|pcif.imemaddr [10]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramaddr~22_combout ),
	.datad(\CPU|CM|daddr [10]),
	.cin(gnd),
	.combout(\ramaddr~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~23 .lut_mask = 16'hE3E0;
defparam \ramaddr~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N16
cycloneive_lcell_comb \ramaddr~24 (
// Equation(s):
// \ramaddr~24_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[13]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdmemWEN) # (ruifdmemREN))))

	.dataa(\syif.addr[13]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datad(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~24 .lut_mask = 16'hBBB8;
defparam \ramaddr~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N22
cycloneive_lcell_comb \ramaddr~25 (
// Equation(s):
// \ramaddr~25_combout  = (\syif.tbCTRL~input_o  & (\ramaddr~24_combout )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~24_combout  & (daddr_13)) # (!\ramaddr~24_combout  & ((pcifimemaddr_13)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\ramaddr~24_combout ),
	.datac(\CPU|CM|daddr [13]),
	.datad(\CPU|DP|pc_dut|pcif.imemaddr [13]),
	.cin(gnd),
	.combout(\ramaddr~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~25 .lut_mask = 16'hD9C8;
defparam \ramaddr~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N0
cycloneive_lcell_comb \ramaddr~26 (
// Equation(s):
// \ramaddr~26_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[12]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdmemWEN) # (ruifdmemREN))))

	.dataa(\syif.addr[12]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datad(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~26 .lut_mask = 16'hBBB8;
defparam \ramaddr~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N10
cycloneive_lcell_comb \ramaddr~27 (
// Equation(s):
// \ramaddr~27_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~26_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~26_combout  & (daddr_12)) # (!\ramaddr~26_combout  & ((pcifimemaddr_12)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [12]),
	.datac(\CPU|DP|pc_dut|pcif.imemaddr [12]),
	.datad(\ramaddr~26_combout ),
	.cin(gnd),
	.combout(\ramaddr~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~27 .lut_mask = 16'hEE50;
defparam \ramaddr~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N28
cycloneive_lcell_comb \ramaddr~28 (
// Equation(s):
// \ramaddr~28_combout  = (ruifdmemREN & (((daddr_15)))) # (!ruifdmemREN & ((ruifdmemWEN & ((daddr_15))) # (!ruifdmemWEN & (pcifimemaddr_15))))

	.dataa(\CPU|DP|pc_dut|pcif.imemaddr [15]),
	.datab(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datac(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datad(\CPU|CM|daddr [15]),
	.cin(gnd),
	.combout(\ramaddr~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~28 .lut_mask = 16'hFE02;
defparam \ramaddr~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N2
cycloneive_lcell_comb \ramaddr~29 (
// Equation(s):
// \ramaddr~29_combout  = (\syif.tbCTRL~input_o  & (!\syif.addr[15]~input_o )) # (!\syif.tbCTRL~input_o  & ((!\ramaddr~28_combout )))

	.dataa(\syif.addr[15]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~28_combout ),
	.cin(gnd),
	.combout(\ramaddr~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~29 .lut_mask = 16'h4477;
defparam \ramaddr~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N18
cycloneive_lcell_comb \ramaddr~30 (
// Equation(s):
// \ramaddr~30_combout  = (ruifdmemWEN & (((daddr_14)))) # (!ruifdmemWEN & ((ruifdmemREN & ((daddr_14))) # (!ruifdmemREN & (pcifimemaddr_14))))

	.dataa(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datab(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datac(\CPU|DP|pc_dut|pcif.imemaddr [14]),
	.datad(\CPU|CM|daddr [14]),
	.cin(gnd),
	.combout(\ramaddr~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~30 .lut_mask = 16'hFE10;
defparam \ramaddr~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N12
cycloneive_lcell_comb \ramaddr~31 (
// Equation(s):
// \ramaddr~31_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[14]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~30_combout )))

	.dataa(\syif.addr[14]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~30_combout ),
	.cin(gnd),
	.combout(\ramaddr~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~31 .lut_mask = 16'hBB88;
defparam \ramaddr~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N0
cycloneive_lcell_comb \ramaddr~32 (
// Equation(s):
// \ramaddr~32_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[17]~input_o )))) # (!\syif.tbCTRL~input_o  & ((ruifdmemREN) # ((ruifdmemWEN))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datac(\syif.addr[17]~input_o ),
	.datad(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~32_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~32 .lut_mask = 16'hF5E4;
defparam \ramaddr~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N10
cycloneive_lcell_comb \ramaddr~33 (
// Equation(s):
// \ramaddr~33_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~32_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~32_combout  & (daddr_17)) # (!\ramaddr~32_combout  & ((pcifimemaddr_17)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [17]),
	.datac(\CPU|DP|pc_dut|pcif.imemaddr [17]),
	.datad(\ramaddr~32_combout ),
	.cin(gnd),
	.combout(\ramaddr~33_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~33 .lut_mask = 16'hEE50;
defparam \ramaddr~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N6
cycloneive_lcell_comb \ramaddr~34 (
// Equation(s):
// \ramaddr~34_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[16]~input_o )))) # (!\syif.tbCTRL~input_o  & (!ruifdmemREN & ((!ruifdmemWEN))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datac(\syif.addr[16]~input_o ),
	.datad(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~34_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~34 .lut_mask = 16'hA0B1;
defparam \ramaddr~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N8
cycloneive_lcell_comb \ramaddr~35 (
// Equation(s):
// \ramaddr~35_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~34_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~34_combout  & (pcifimemaddr_16)) # (!\ramaddr~34_combout  & ((daddr_16)))))

	.dataa(\CPU|DP|pc_dut|pcif.imemaddr [16]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|CM|daddr [16]),
	.datad(\ramaddr~34_combout ),
	.cin(gnd),
	.combout(\ramaddr~35_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~35 .lut_mask = 16'hEE30;
defparam \ramaddr~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N6
cycloneive_lcell_comb \ramaddr~36 (
// Equation(s):
// \ramaddr~36_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[19]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdmemWEN) # (ruifdmemREN))))

	.dataa(\syif.addr[19]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datad(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~36_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~36 .lut_mask = 16'hBBB8;
defparam \ramaddr~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N28
cycloneive_lcell_comb \ramaddr~37 (
// Equation(s):
// \ramaddr~37_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~36_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~36_combout  & (daddr_19)) # (!\ramaddr~36_combout  & ((pcifimemaddr_19)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [19]),
	.datac(\CPU|DP|pc_dut|pcif.imemaddr [19]),
	.datad(\ramaddr~36_combout ),
	.cin(gnd),
	.combout(\ramaddr~37_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~37 .lut_mask = 16'hEE50;
defparam \ramaddr~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N18
cycloneive_lcell_comb \ramaddr~38 (
// Equation(s):
// \ramaddr~38_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[18]~input_o )))) # (!\syif.tbCTRL~input_o  & ((ruifdmemREN) # ((ruifdmemWEN))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datac(\syif.addr[18]~input_o ),
	.datad(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~38_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~38 .lut_mask = 16'hF5E4;
defparam \ramaddr~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N20
cycloneive_lcell_comb \ramaddr~39 (
// Equation(s):
// \ramaddr~39_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~38_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~38_combout  & ((daddr_18))) # (!\ramaddr~38_combout  & (pcifimemaddr_18))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|pc_dut|pcif.imemaddr [18]),
	.datac(\CPU|CM|daddr [18]),
	.datad(\ramaddr~38_combout ),
	.cin(gnd),
	.combout(\ramaddr~39_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~39 .lut_mask = 16'hFA44;
defparam \ramaddr~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N20
cycloneive_lcell_comb \ramaddr~40 (
// Equation(s):
// \ramaddr~40_combout  = (ruifdmemREN & (daddr_21)) # (!ruifdmemREN & ((ruifdmemWEN & (daddr_21)) # (!ruifdmemWEN & ((pcifimemaddr_21)))))

	.dataa(\CPU|CM|daddr [21]),
	.datab(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datac(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datad(\CPU|DP|pc_dut|pcif.imemaddr [21]),
	.cin(gnd),
	.combout(\ramaddr~40_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~40 .lut_mask = 16'hABA8;
defparam \ramaddr~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N16
cycloneive_lcell_comb \ramaddr~41 (
// Equation(s):
// \ramaddr~41_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[21]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~40_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[21]~input_o ),
	.datad(\ramaddr~40_combout ),
	.cin(gnd),
	.combout(\ramaddr~41_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~41 .lut_mask = 16'hF5A0;
defparam \ramaddr~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N2
cycloneive_lcell_comb \ramaddr~42 (
// Equation(s):
// \ramaddr~42_combout  = (ruifdmemREN & (daddr_20)) # (!ruifdmemREN & ((ruifdmemWEN & (daddr_20)) # (!ruifdmemWEN & ((pcifimemaddr_20)))))

	.dataa(\CPU|CM|daddr [20]),
	.datab(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datac(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datad(\CPU|DP|pc_dut|pcif.imemaddr [20]),
	.cin(gnd),
	.combout(\ramaddr~42_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~42 .lut_mask = 16'hABA8;
defparam \ramaddr~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N24
cycloneive_lcell_comb \ramaddr~43 (
// Equation(s):
// \ramaddr~43_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[20]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~42_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[20]~input_o ),
	.datad(\ramaddr~42_combout ),
	.cin(gnd),
	.combout(\ramaddr~43_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~43 .lut_mask = 16'hF5A0;
defparam \ramaddr~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N16
cycloneive_lcell_comb \ramaddr~44 (
// Equation(s):
// \ramaddr~44_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[23]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdmemWEN) # (ruifdmemREN))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[23]~input_o ),
	.datac(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datad(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~44_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~44 .lut_mask = 16'hDDD8;
defparam \ramaddr~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N30
cycloneive_lcell_comb \ramaddr~45 (
// Equation(s):
// \ramaddr~45_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~44_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~44_combout  & (daddr_23)) # (!\ramaddr~44_combout  & ((pcifimemaddr_23)))))

	.dataa(\CPU|CM|daddr [23]),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|pc_dut|pcif.imemaddr [23]),
	.datad(\ramaddr~44_combout ),
	.cin(gnd),
	.combout(\ramaddr~45_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~45 .lut_mask = 16'hEE30;
defparam \ramaddr~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N2
cycloneive_lcell_comb \ramaddr~46 (
// Equation(s):
// \ramaddr~46_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[22]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdmemWEN) # (ruifdmemREN))))

	.dataa(\syif.addr[22]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datad(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~46_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~46 .lut_mask = 16'hBBB8;
defparam \ramaddr~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N0
cycloneive_lcell_comb \ramaddr~47 (
// Equation(s):
// \ramaddr~47_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~46_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~46_combout  & ((daddr_22))) # (!\ramaddr~46_combout  & (pcifimemaddr_22))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|pc_dut|pcif.imemaddr [22]),
	.datac(\CPU|CM|daddr [22]),
	.datad(\ramaddr~46_combout ),
	.cin(gnd),
	.combout(\ramaddr~47_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~47 .lut_mask = 16'hFA44;
defparam \ramaddr~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N24
cycloneive_lcell_comb \ramaddr~48 (
// Equation(s):
// \ramaddr~48_combout  = (ruifdmemREN & (daddr_25)) # (!ruifdmemREN & ((ruifdmemWEN & (daddr_25)) # (!ruifdmemWEN & ((pcifimemaddr_25)))))

	.dataa(\CPU|CM|daddr [25]),
	.datab(\CPU|DP|pc_dut|pcif.imemaddr [25]),
	.datac(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datad(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~48_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~48 .lut_mask = 16'hAAAC;
defparam \ramaddr~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N12
cycloneive_lcell_comb \ramaddr~49 (
// Equation(s):
// \ramaddr~49_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[25]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~48_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[25]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~48_combout ),
	.cin(gnd),
	.combout(\ramaddr~49_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~49 .lut_mask = 16'hDD88;
defparam \ramaddr~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N20
cycloneive_lcell_comb \ramaddr~50 (
// Equation(s):
// \ramaddr~50_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[24]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdmemREN) # (ruifdmemWEN))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[24]~input_o ),
	.datac(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datad(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~50_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~50 .lut_mask = 16'hDDD8;
defparam \ramaddr~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N22
cycloneive_lcell_comb \ramaddr~51 (
// Equation(s):
// \ramaddr~51_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~50_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~50_combout  & (daddr_24)) # (!\ramaddr~50_combout  & ((pcifimemaddr_24)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [24]),
	.datac(\CPU|DP|pc_dut|pcif.imemaddr [24]),
	.datad(\ramaddr~50_combout ),
	.cin(gnd),
	.combout(\ramaddr~51_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~51 .lut_mask = 16'hEE50;
defparam \ramaddr~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N26
cycloneive_lcell_comb \ramaddr~52 (
// Equation(s):
// \ramaddr~52_combout  = (\syif.tbCTRL~input_o  & (((\syif.addr[27]~input_o )))) # (!\syif.tbCTRL~input_o  & ((ruifdmemREN) # ((ruifdmemWEN))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datac(\syif.addr[27]~input_o ),
	.datad(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~52_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~52 .lut_mask = 16'hF5E4;
defparam \ramaddr~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N24
cycloneive_lcell_comb \ramaddr~53 (
// Equation(s):
// \ramaddr~53_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~52_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~52_combout  & (daddr_27)) # (!\ramaddr~52_combout  & ((pcifimemaddr_27)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [27]),
	.datac(\ramaddr~52_combout ),
	.datad(\CPU|DP|pc_dut|pcif.imemaddr [27]),
	.cin(gnd),
	.combout(\ramaddr~53_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~53 .lut_mask = 16'hE5E0;
defparam \ramaddr~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N2
cycloneive_lcell_comb \ramaddr~54 (
// Equation(s):
// \ramaddr~54_combout  = (ruifdmemREN & (daddr_26)) # (!ruifdmemREN & ((ruifdmemWEN & (daddr_26)) # (!ruifdmemWEN & ((pcifimemaddr_26)))))

	.dataa(\CPU|CM|daddr [26]),
	.datab(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datac(\CPU|DP|pc_dut|pcif.imemaddr [26]),
	.datad(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~54_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~54 .lut_mask = 16'hAAB8;
defparam \ramaddr~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N16
cycloneive_lcell_comb \ramaddr~55 (
// Equation(s):
// \ramaddr~55_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[26]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~54_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[26]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~54_combout ),
	.cin(gnd),
	.combout(\ramaddr~55_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~55 .lut_mask = 16'hDD88;
defparam \ramaddr~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N22
cycloneive_lcell_comb \ramaddr~56 (
// Equation(s):
// \ramaddr~56_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[29]~input_o )) # (!\syif.tbCTRL~input_o  & (((ruifdmemWEN) # (ruifdmemREN))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[29]~input_o ),
	.datac(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datad(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~56_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~56 .lut_mask = 16'hDDD8;
defparam \ramaddr~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N8
cycloneive_lcell_comb \ramaddr~57 (
// Equation(s):
// \ramaddr~57_combout  = (\syif.tbCTRL~input_o  & (((\ramaddr~56_combout )))) # (!\syif.tbCTRL~input_o  & ((\ramaddr~56_combout  & (daddr_29)) # (!\ramaddr~56_combout  & ((pcifimemaddr_29)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|CM|daddr [29]),
	.datac(\ramaddr~56_combout ),
	.datad(\CPU|DP|pc_dut|pcif.imemaddr [29]),
	.cin(gnd),
	.combout(\ramaddr~57_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~57 .lut_mask = 16'hE5E0;
defparam \ramaddr~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N16
cycloneive_lcell_comb \ramaddr~58 (
// Equation(s):
// \ramaddr~58_combout  = (ruifdmemWEN & (daddr_28)) # (!ruifdmemWEN & ((ruifdmemREN & (daddr_28)) # (!ruifdmemREN & ((pcifimemaddr_28)))))

	.dataa(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datab(\CPU|CM|daddr [28]),
	.datac(\CPU|DP|pc_dut|pcif.imemaddr [28]),
	.datad(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.cin(gnd),
	.combout(\ramaddr~58_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~58 .lut_mask = 16'hCCD8;
defparam \ramaddr~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N2
cycloneive_lcell_comb \ramaddr~59 (
// Equation(s):
// \ramaddr~59_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[28]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~58_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[28]~input_o ),
	.datad(\ramaddr~58_combout ),
	.cin(gnd),
	.combout(\ramaddr~59_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~59 .lut_mask = 16'hF5A0;
defparam \ramaddr~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N16
cycloneive_lcell_comb \ramaddr~60 (
// Equation(s):
// \ramaddr~60_combout  = (ruifdmemREN & (daddr_31)) # (!ruifdmemREN & ((ruifdmemWEN & (daddr_31)) # (!ruifdmemWEN & ((pcifimemaddr_31)))))

	.dataa(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datab(\CPU|CM|daddr [31]),
	.datac(\CPU|DP|pc_dut|pcif.imemaddr [31]),
	.datad(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~60_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~60 .lut_mask = 16'hCCD8;
defparam \ramaddr~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N10
cycloneive_lcell_comb \ramaddr~61 (
// Equation(s):
// \ramaddr~61_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[31]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~60_combout )))

	.dataa(\syif.addr[31]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~60_combout ),
	.cin(gnd),
	.combout(\ramaddr~61_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~61 .lut_mask = 16'hBB88;
defparam \ramaddr~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N24
cycloneive_lcell_comb \ramaddr~62 (
// Equation(s):
// \ramaddr~62_combout  = (ruifdmemREN & (daddr_30)) # (!ruifdmemREN & ((ruifdmemWEN & (daddr_30)) # (!ruifdmemWEN & ((pcifimemaddr_30)))))

	.dataa(\CPU|DP|ru_dut|ruif.dmemREN~q ),
	.datab(\CPU|CM|daddr [30]),
	.datac(\CPU|DP|pc_dut|pcif.imemaddr [30]),
	.datad(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.cin(gnd),
	.combout(\ramaddr~62_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~62 .lut_mask = 16'hCCD8;
defparam \ramaddr~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N18
cycloneive_lcell_comb \ramaddr~63 (
// Equation(s):
// \ramaddr~63_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[30]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~62_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[30]~input_o ),
	.datad(\ramaddr~62_combout ),
	.cin(gnd),
	.combout(\ramaddr~63_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~63 .lut_mask = 16'hF3C0;
defparam \ramaddr~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N0
cycloneive_lcell_comb \ramWEN~0 (
// Equation(s):
// \ramWEN~0_combout  = (\syif.tbCTRL~input_o  & (!\syif.WEN~input_o )) # (!\syif.tbCTRL~input_o  & ((!ruifdmemWEN)))

	.dataa(gnd),
	.datab(\syif.WEN~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.cin(gnd),
	.combout(\ramWEN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramWEN~0 .lut_mask = 16'h303F;
defparam \ramWEN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N4
cycloneive_lcell_comb \ramREN~0 (
// Equation(s):
// \ramREN~0_combout  = (\syif.tbCTRL~input_o  & ((!\syif.REN~input_o ))) # (!\syif.tbCTRL~input_o  & (ruifdmemWEN))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|ru_dut|ruif.dmemWEN~q ),
	.datac(\syif.REN~input_o ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramREN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramREN~0 .lut_mask = 16'h4E4E;
defparam \ramREN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X114_Y37_N17
dffeas CPUCLK(
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\CPUCLK~0_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\CPUCLK~q ),
	.prn(vcc));
// synopsys translate_off
defparam CPUCLK.is_wysiwyg = "true";
defparam CPUCLK.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N24
cycloneive_lcell_comb \ramstore~0 (
// Equation(s):
// \ramstore~0_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux63)) # (!cuifregT_4 & ((Mux631)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|rf_dut|Mux63~9_combout ),
	.datac(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datad(\CPU|DP|rf_dut|Mux63~19_combout ),
	.cin(gnd),
	.combout(\ramstore~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~0 .lut_mask = 16'h4540;
defparam \ramstore~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N26
cycloneive_lcell_comb \ramstore~1 (
// Equation(s):
// \ramstore~1_combout  = (\ramstore~0_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[0]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[0]~input_o ),
	.datac(gnd),
	.datad(\ramstore~0_combout ),
	.cin(gnd),
	.combout(\ramstore~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~1 .lut_mask = 16'hFF88;
defparam \ramstore~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N24
cycloneive_lcell_comb \ramstore~2 (
// Equation(s):
// \ramstore~2_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux621)) # (!cuifregT_4 & ((Mux62)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datac(\CPU|DP|rf_dut|Mux62~19_combout ),
	.datad(\CPU|DP|rf_dut|Mux62~9_combout ),
	.cin(gnd),
	.combout(\ramstore~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~2 .lut_mask = 16'h5140;
defparam \ramstore~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N14
cycloneive_lcell_comb \ramstore~3 (
// Equation(s):
// \ramstore~3_combout  = (\ramstore~2_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[1]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[1]~input_o ),
	.datad(\ramstore~2_combout ),
	.cin(gnd),
	.combout(\ramstore~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~3 .lut_mask = 16'hFFC0;
defparam \ramstore~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N6
cycloneive_lcell_comb \ramstore~4 (
// Equation(s):
// \ramstore~4_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux61)) # (!cuifregT_4 & ((Mux611)))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf_dut|Mux61~9_combout ),
	.datad(\CPU|DP|rf_dut|Mux61~19_combout ),
	.cin(gnd),
	.combout(\ramstore~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~4 .lut_mask = 16'h3120;
defparam \ramstore~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N28
cycloneive_lcell_comb \ramstore~5 (
// Equation(s):
// \ramstore~5_combout  = (\ramstore~4_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[2]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[2]~input_o ),
	.datad(\ramstore~4_combout ),
	.cin(gnd),
	.combout(\ramstore~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~5 .lut_mask = 16'hFFC0;
defparam \ramstore~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N6
cycloneive_lcell_comb \ramstore~6 (
// Equation(s):
// \ramstore~6_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux60)) # (!cuifregT_4 & ((Mux601)))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\CPU|DP|rf_dut|Mux60~9_combout ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rf_dut|Mux60~19_combout ),
	.cin(gnd),
	.combout(\ramstore~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~6 .lut_mask = 16'h0D08;
defparam \ramstore~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N28
cycloneive_lcell_comb \ramstore~7 (
// Equation(s):
// \ramstore~7_combout  = (\ramstore~6_combout ) # ((\syif.store[3]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[3]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~6_combout ),
	.cin(gnd),
	.combout(\ramstore~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~7 .lut_mask = 16'hFFA0;
defparam \ramstore~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N18
cycloneive_lcell_comb \ramstore~8 (
// Equation(s):
// \ramstore~8_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux59)) # (!cuifregT_4 & ((Mux591)))))

	.dataa(\CPU|DP|rf_dut|Mux59~9_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datad(\CPU|DP|rf_dut|Mux59~19_combout ),
	.cin(gnd),
	.combout(\ramstore~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~8 .lut_mask = 16'h2320;
defparam \ramstore~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N12
cycloneive_lcell_comb \ramstore~9 (
// Equation(s):
// \ramstore~9_combout  = (\ramstore~8_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[4]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[4]~input_o ),
	.datad(\ramstore~8_combout ),
	.cin(gnd),
	.combout(\ramstore~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~9 .lut_mask = 16'hFFA0;
defparam \ramstore~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N6
cycloneive_lcell_comb \ramstore~10 (
// Equation(s):
// \ramstore~10_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux581)) # (!cuifregT_4 & ((Mux58)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datac(\CPU|DP|rf_dut|Mux58~19_combout ),
	.datad(\CPU|DP|rf_dut|Mux58~9_combout ),
	.cin(gnd),
	.combout(\ramstore~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~10 .lut_mask = 16'h5140;
defparam \ramstore~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N16
cycloneive_lcell_comb \ramstore~11 (
// Equation(s):
// \ramstore~11_combout  = (\ramstore~10_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[5]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[5]~input_o ),
	.datac(gnd),
	.datad(\ramstore~10_combout ),
	.cin(gnd),
	.combout(\ramstore~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~11 .lut_mask = 16'hFF88;
defparam \ramstore~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N12
cycloneive_lcell_comb \ramstore~12 (
// Equation(s):
// \ramstore~12_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & ((Mux571))) # (!cuifregT_4 & (Mux57))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf_dut|Mux57~9_combout ),
	.datad(\CPU|DP|rf_dut|Mux57~19_combout ),
	.cin(gnd),
	.combout(\ramstore~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~12 .lut_mask = 16'h3210;
defparam \ramstore~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N22
cycloneive_lcell_comb \ramstore~13 (
// Equation(s):
// \ramstore~13_combout  = (\ramstore~12_combout ) # ((\syif.store[6]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(\syif.store[6]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~12_combout ),
	.cin(gnd),
	.combout(\ramstore~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~13 .lut_mask = 16'hFFC0;
defparam \ramstore~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N12
cycloneive_lcell_comb \ramstore~14 (
// Equation(s):
// \ramstore~14_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux561)) # (!cuifregT_4 & ((Mux56)))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf_dut|Mux56~19_combout ),
	.datad(\CPU|DP|rf_dut|Mux56~9_combout ),
	.cin(gnd),
	.combout(\ramstore~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~14 .lut_mask = 16'h3120;
defparam \ramstore~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N22
cycloneive_lcell_comb \ramstore~15 (
// Equation(s):
// \ramstore~15_combout  = (\ramstore~14_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[7]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[7]~input_o ),
	.datad(\ramstore~14_combout ),
	.cin(gnd),
	.combout(\ramstore~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~15 .lut_mask = 16'hFFC0;
defparam \ramstore~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N28
cycloneive_lcell_comb \ramstore~16 (
// Equation(s):
// \ramstore~16_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux551)) # (!cuifregT_4 & ((Mux55)))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\CPU|DP|rf_dut|Mux55~19_combout ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rf_dut|Mux55~9_combout ),
	.cin(gnd),
	.combout(\ramstore~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~16 .lut_mask = 16'h0D08;
defparam \ramstore~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N22
cycloneive_lcell_comb \ramstore~17 (
// Equation(s):
// \ramstore~17_combout  = (\ramstore~16_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[8]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[8]~input_o ),
	.datac(gnd),
	.datad(\ramstore~16_combout ),
	.cin(gnd),
	.combout(\ramstore~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~17 .lut_mask = 16'hFF88;
defparam \ramstore~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N28
cycloneive_lcell_comb \ramstore~18 (
// Equation(s):
// \ramstore~18_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux541)) # (!cuifregT_4 & ((Mux54)))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\CPU|DP|rf_dut|Mux54~19_combout ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rf_dut|Mux54~9_combout ),
	.cin(gnd),
	.combout(\ramstore~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~18 .lut_mask = 16'h0D08;
defparam \ramstore~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N14
cycloneive_lcell_comb \ramstore~19 (
// Equation(s):
// \ramstore~19_combout  = (\ramstore~18_combout ) # ((\syif.store[9]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[9]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~18_combout ),
	.cin(gnd),
	.combout(\ramstore~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~19 .lut_mask = 16'hFFA0;
defparam \ramstore~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N20
cycloneive_lcell_comb \ramstore~20 (
// Equation(s):
// \ramstore~20_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux531)) # (!cuifregT_4 & ((Mux53)))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf_dut|Mux53~19_combout ),
	.datad(\CPU|DP|rf_dut|Mux53~9_combout ),
	.cin(gnd),
	.combout(\ramstore~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~20 .lut_mask = 16'h3120;
defparam \ramstore~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N30
cycloneive_lcell_comb \ramstore~21 (
// Equation(s):
// \ramstore~21_combout  = (\ramstore~20_combout ) # ((\syif.store[10]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(\syif.store[10]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~20_combout ),
	.cin(gnd),
	.combout(\ramstore~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~21 .lut_mask = 16'hFFC0;
defparam \ramstore~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N16
cycloneive_lcell_comb \ramstore~22 (
// Equation(s):
// \ramstore~22_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & ((Mux521))) # (!cuifregT_4 & (Mux52))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf_dut|Mux52~9_combout ),
	.datad(\CPU|DP|rf_dut|Mux52~19_combout ),
	.cin(gnd),
	.combout(\ramstore~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~22 .lut_mask = 16'h3210;
defparam \ramstore~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N26
cycloneive_lcell_comb \ramstore~23 (
// Equation(s):
// \ramstore~23_combout  = (\ramstore~22_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[11]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[11]~input_o ),
	.datad(\ramstore~22_combout ),
	.cin(gnd),
	.combout(\ramstore~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~23 .lut_mask = 16'hFFC0;
defparam \ramstore~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N30
cycloneive_lcell_comb \ramstore~24 (
// Equation(s):
// \ramstore~24_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux511)) # (!cuifregT_4 & ((Mux51)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datac(\CPU|DP|rf_dut|Mux51~19_combout ),
	.datad(\CPU|DP|rf_dut|Mux51~9_combout ),
	.cin(gnd),
	.combout(\ramstore~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~24 .lut_mask = 16'h5140;
defparam \ramstore~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N28
cycloneive_lcell_comb \ramstore~25 (
// Equation(s):
// \ramstore~25_combout  = (\ramstore~24_combout ) # ((\syif.store[12]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\ramstore~24_combout ),
	.datab(\syif.store[12]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramstore~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~25 .lut_mask = 16'hEAEA;
defparam \ramstore~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N12
cycloneive_lcell_comb \ramstore~26 (
// Equation(s):
// \ramstore~26_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux501)) # (!cuifregT_4 & ((Mux50)))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\CPU|DP|rf_dut|Mux50~19_combout ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rf_dut|Mux50~9_combout ),
	.cin(gnd),
	.combout(\ramstore~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~26 .lut_mask = 16'h0D08;
defparam \ramstore~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N18
cycloneive_lcell_comb \ramstore~27 (
// Equation(s):
// \ramstore~27_combout  = (\ramstore~26_combout ) # ((\syif.store[13]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(\syif.store[13]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~26_combout ),
	.cin(gnd),
	.combout(\ramstore~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~27 .lut_mask = 16'hFFC0;
defparam \ramstore~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N12
cycloneive_lcell_comb \ramstore~28 (
// Equation(s):
// \ramstore~28_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux491)) # (!cuifregT_4 & ((Mux49)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datac(\CPU|DP|rf_dut|Mux49~19_combout ),
	.datad(\CPU|DP|rf_dut|Mux49~9_combout ),
	.cin(gnd),
	.combout(\ramstore~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~28 .lut_mask = 16'h5140;
defparam \ramstore~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N6
cycloneive_lcell_comb \ramstore~29 (
// Equation(s):
// \ramstore~29_combout  = (\ramstore~28_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[14]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[14]~input_o ),
	.datad(\ramstore~28_combout ),
	.cin(gnd),
	.combout(\ramstore~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~29 .lut_mask = 16'hFFA0;
defparam \ramstore~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N12
cycloneive_lcell_comb \ramstore~30 (
// Equation(s):
// \ramstore~30_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & ((Mux481))) # (!cuifregT_4 & (Mux48))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\CPU|DP|rf_dut|Mux48~9_combout ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rf_dut|Mux48~19_combout ),
	.cin(gnd),
	.combout(\ramstore~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~30 .lut_mask = 16'h0E04;
defparam \ramstore~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N30
cycloneive_lcell_comb \ramstore~31 (
// Equation(s):
// \ramstore~31_combout  = (\ramstore~30_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[15]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[15]~input_o ),
	.datad(\ramstore~30_combout ),
	.cin(gnd),
	.combout(\ramstore~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~31 .lut_mask = 16'hFFA0;
defparam \ramstore~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N16
cycloneive_lcell_comb \ramstore~32 (
// Equation(s):
// \ramstore~32_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & ((Mux47))) # (!cuifregT_4 & (Mux471))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\CPU|DP|rf_dut|Mux47~19_combout ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rf_dut|Mux47~9_combout ),
	.cin(gnd),
	.combout(\ramstore~32_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~32 .lut_mask = 16'h0E04;
defparam \ramstore~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N18
cycloneive_lcell_comb \ramstore~33 (
// Equation(s):
// \ramstore~33_combout  = (\ramstore~32_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[16]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[16]~input_o ),
	.datad(\ramstore~32_combout ),
	.cin(gnd),
	.combout(\ramstore~33_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~33 .lut_mask = 16'hFFC0;
defparam \ramstore~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N10
cycloneive_lcell_comb \ramstore~34 (
// Equation(s):
// \ramstore~34_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux461)) # (!cuifregT_4 & ((Mux46)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datac(\CPU|DP|rf_dut|Mux46~19_combout ),
	.datad(\CPU|DP|rf_dut|Mux46~9_combout ),
	.cin(gnd),
	.combout(\ramstore~34_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~34 .lut_mask = 16'h5140;
defparam \ramstore~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N28
cycloneive_lcell_comb \ramstore~35 (
// Equation(s):
// \ramstore~35_combout  = (\ramstore~34_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[17]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[17]~input_o ),
	.datad(\ramstore~34_combout ),
	.cin(gnd),
	.combout(\ramstore~35_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~35 .lut_mask = 16'hFFC0;
defparam \ramstore~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N2
cycloneive_lcell_comb \ramstore~36 (
// Equation(s):
// \ramstore~36_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & ((Mux451))) # (!cuifregT_4 & (Mux45))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\CPU|DP|rf_dut|Mux45~9_combout ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rf_dut|Mux45~19_combout ),
	.cin(gnd),
	.combout(\ramstore~36_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~36 .lut_mask = 16'h0E04;
defparam \ramstore~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N8
cycloneive_lcell_comb \ramstore~37 (
// Equation(s):
// \ramstore~37_combout  = (\ramstore~36_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[18]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[18]~input_o ),
	.datad(\ramstore~36_combout ),
	.cin(gnd),
	.combout(\ramstore~37_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~37 .lut_mask = 16'hFFC0;
defparam \ramstore~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N22
cycloneive_lcell_comb \ramstore~38 (
// Equation(s):
// \ramstore~38_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & ((Mux441))) # (!cuifregT_4 & (Mux44))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datac(\CPU|DP|rf_dut|Mux44~9_combout ),
	.datad(\CPU|DP|rf_dut|Mux44~19_combout ),
	.cin(gnd),
	.combout(\ramstore~38_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~38 .lut_mask = 16'h5410;
defparam \ramstore~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N22
cycloneive_lcell_comb \ramstore~39 (
// Equation(s):
// \ramstore~39_combout  = (\ramstore~38_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[19]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[19]~input_o ),
	.datad(\ramstore~38_combout ),
	.cin(gnd),
	.combout(\ramstore~39_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~39 .lut_mask = 16'hFFA0;
defparam \ramstore~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N20
cycloneive_lcell_comb \ramstore~40 (
// Equation(s):
// \ramstore~40_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux431)) # (!cuifregT_4 & ((Mux43)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datac(\CPU|DP|rf_dut|Mux43~19_combout ),
	.datad(\CPU|DP|rf_dut|Mux43~9_combout ),
	.cin(gnd),
	.combout(\ramstore~40_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~40 .lut_mask = 16'h5140;
defparam \ramstore~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N6
cycloneive_lcell_comb \ramstore~41 (
// Equation(s):
// \ramstore~41_combout  = (\ramstore~40_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[20]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[20]~input_o ),
	.datac(gnd),
	.datad(\ramstore~40_combout ),
	.cin(gnd),
	.combout(\ramstore~41_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~41 .lut_mask = 16'hFF88;
defparam \ramstore~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N20
cycloneive_lcell_comb \ramstore~42 (
// Equation(s):
// \ramstore~42_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & ((Mux421))) # (!cuifregT_4 & (Mux42))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datac(\CPU|DP|rf_dut|Mux42~9_combout ),
	.datad(\CPU|DP|rf_dut|Mux42~19_combout ),
	.cin(gnd),
	.combout(\ramstore~42_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~42 .lut_mask = 16'h5410;
defparam \ramstore~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N6
cycloneive_lcell_comb \ramstore~43 (
// Equation(s):
// \ramstore~43_combout  = (\ramstore~42_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[21]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[21]~input_o ),
	.datad(\ramstore~42_combout ),
	.cin(gnd),
	.combout(\ramstore~43_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~43 .lut_mask = 16'hFFA0;
defparam \ramstore~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N24
cycloneive_lcell_comb \ramstore~44 (
// Equation(s):
// \ramstore~44_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux411)) # (!cuifregT_4 & ((Mux41)))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf_dut|Mux41~19_combout ),
	.datad(\CPU|DP|rf_dut|Mux41~9_combout ),
	.cin(gnd),
	.combout(\ramstore~44_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~44 .lut_mask = 16'h3120;
defparam \ramstore~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N26
cycloneive_lcell_comb \ramstore~45 (
// Equation(s):
// \ramstore~45_combout  = (\ramstore~44_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[22]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[22]~input_o ),
	.datad(\ramstore~44_combout ),
	.cin(gnd),
	.combout(\ramstore~45_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~45 .lut_mask = 16'hFFC0;
defparam \ramstore~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N28
cycloneive_lcell_comb \ramstore~46 (
// Equation(s):
// \ramstore~46_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & ((Mux401))) # (!cuifregT_4 & (Mux40))))

	.dataa(\CPU|DP|rf_dut|Mux40~9_combout ),
	.datab(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|rf_dut|Mux40~19_combout ),
	.cin(gnd),
	.combout(\ramstore~46_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~46 .lut_mask = 16'h0E02;
defparam \ramstore~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N30
cycloneive_lcell_comb \ramstore~47 (
// Equation(s):
// \ramstore~47_combout  = (\ramstore~46_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[23]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[23]~input_o ),
	.datad(\ramstore~46_combout ),
	.cin(gnd),
	.combout(\ramstore~47_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~47 .lut_mask = 16'hFFC0;
defparam \ramstore~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N30
cycloneive_lcell_comb \ramstore~48 (
// Equation(s):
// \ramstore~48_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & ((Mux39))) # (!cuifregT_4 & (Mux391))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf_dut|Mux39~19_combout ),
	.datad(\CPU|DP|rf_dut|Mux39~9_combout ),
	.cin(gnd),
	.combout(\ramstore~48_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~48 .lut_mask = 16'h3210;
defparam \ramstore~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N28
cycloneive_lcell_comb \ramstore~49 (
// Equation(s):
// \ramstore~49_combout  = (\ramstore~48_combout ) # ((\syif.store[24]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[24]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramstore~48_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramstore~49_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~49 .lut_mask = 16'hF8F8;
defparam \ramstore~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N10
cycloneive_lcell_comb \ramstore~50 (
// Equation(s):
// \ramstore~50_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux381)) # (!cuifregT_4 & ((Mux38)))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf_dut|Mux38~19_combout ),
	.datad(\CPU|DP|rf_dut|Mux38~9_combout ),
	.cin(gnd),
	.combout(\ramstore~50_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~50 .lut_mask = 16'h3120;
defparam \ramstore~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N12
cycloneive_lcell_comb \ramstore~51 (
// Equation(s):
// \ramstore~51_combout  = (\ramstore~50_combout ) # ((\syif.store[25]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(\syif.store[25]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~50_combout ),
	.cin(gnd),
	.combout(\ramstore~51_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~51 .lut_mask = 16'hFFC0;
defparam \ramstore~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N2
cycloneive_lcell_comb \ramstore~52 (
// Equation(s):
// \ramstore~52_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & ((Mux371))) # (!cuifregT_4 & (Mux37))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf_dut|Mux37~9_combout ),
	.datad(\CPU|DP|rf_dut|Mux37~19_combout ),
	.cin(gnd),
	.combout(\ramstore~52_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~52 .lut_mask = 16'h3210;
defparam \ramstore~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N28
cycloneive_lcell_comb \ramstore~53 (
// Equation(s):
// \ramstore~53_combout  = (\ramstore~52_combout ) # ((\syif.store[26]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(\syif.store[26]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramstore~52_combout ),
	.cin(gnd),
	.combout(\ramstore~53_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~53 .lut_mask = 16'hFF88;
defparam \ramstore~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N30
cycloneive_lcell_comb \ramstore~54 (
// Equation(s):
// \ramstore~54_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux361)) # (!cuifregT_4 & ((Mux36)))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf_dut|Mux36~19_combout ),
	.datad(\CPU|DP|rf_dut|Mux36~9_combout ),
	.cin(gnd),
	.combout(\ramstore~54_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~54 .lut_mask = 16'h3120;
defparam \ramstore~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N0
cycloneive_lcell_comb \ramstore~55 (
// Equation(s):
// \ramstore~55_combout  = (\ramstore~54_combout ) # ((\syif.store[27]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(\syif.store[27]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramstore~54_combout ),
	.cin(gnd),
	.combout(\ramstore~55_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~55 .lut_mask = 16'hFFC0;
defparam \ramstore~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N28
cycloneive_lcell_comb \ramstore~56 (
// Equation(s):
// \ramstore~56_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux351)) # (!cuifregT_4 & ((Mux35)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datac(\CPU|DP|rf_dut|Mux35~19_combout ),
	.datad(\CPU|DP|rf_dut|Mux35~9_combout ),
	.cin(gnd),
	.combout(\ramstore~56_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~56 .lut_mask = 16'h5140;
defparam \ramstore~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N18
cycloneive_lcell_comb \ramstore~57 (
// Equation(s):
// \ramstore~57_combout  = (\ramstore~56_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[28]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.store[28]~input_o ),
	.datac(gnd),
	.datad(\ramstore~56_combout ),
	.cin(gnd),
	.combout(\ramstore~57_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~57 .lut_mask = 16'hFF88;
defparam \ramstore~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N10
cycloneive_lcell_comb \ramstore~58 (
// Equation(s):
// \ramstore~58_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux34)) # (!cuifregT_4 & ((Mux341)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datac(\CPU|DP|rf_dut|Mux34~9_combout ),
	.datad(\CPU|DP|rf_dut|Mux34~19_combout ),
	.cin(gnd),
	.combout(\ramstore~58_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~58 .lut_mask = 16'h5140;
defparam \ramstore~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N10
cycloneive_lcell_comb \ramstore~59 (
// Equation(s):
// \ramstore~59_combout  = (\ramstore~58_combout ) # ((\syif.store[29]~input_o  & \syif.tbCTRL~input_o ))

	.dataa(gnd),
	.datab(\syif.store[29]~input_o ),
	.datac(\ramstore~58_combout ),
	.datad(\syif.tbCTRL~input_o ),
	.cin(gnd),
	.combout(\ramstore~59_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~59 .lut_mask = 16'hFCF0;
defparam \ramstore~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N16
cycloneive_lcell_comb \ramstore~60 (
// Equation(s):
// \ramstore~60_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & ((Mux331))) # (!cuifregT_4 & (Mux33))))

	.dataa(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|rf_dut|Mux33~9_combout ),
	.datad(\CPU|DP|rf_dut|Mux33~19_combout ),
	.cin(gnd),
	.combout(\ramstore~60_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~60 .lut_mask = 16'h3210;
defparam \ramstore~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N6
cycloneive_lcell_comb \ramstore~61 (
// Equation(s):
// \ramstore~61_combout  = (\ramstore~60_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[30]~input_o ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[30]~input_o ),
	.datad(\ramstore~60_combout ),
	.cin(gnd),
	.combout(\ramstore~61_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~61 .lut_mask = 16'hFFC0;
defparam \ramstore~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N20
cycloneive_lcell_comb \ramstore~62 (
// Equation(s):
// \ramstore~62_combout  = (!\syif.tbCTRL~input_o  & ((cuifregT_4 & (Mux32)) # (!cuifregT_4 & ((Mux321)))))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\CPU|DP|cu_dut|cuif.regT[4]~6_combout ),
	.datac(\CPU|DP|rf_dut|Mux32~9_combout ),
	.datad(\CPU|DP|rf_dut|Mux32~19_combout ),
	.cin(gnd),
	.combout(\ramstore~62_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~62 .lut_mask = 16'h5140;
defparam \ramstore~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N14
cycloneive_lcell_comb \ramstore~63 (
// Equation(s):
// \ramstore~63_combout  = (\ramstore~62_combout ) # ((\syif.tbCTRL~input_o  & \syif.store[31]~input_o ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.store[31]~input_o ),
	.datad(\ramstore~62_combout ),
	.cin(gnd),
	.combout(\ramstore~63_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~63 .lut_mask = 16'hFFA0;
defparam \ramstore~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X114_Y36_N1
dffeas \count[3] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[3]~0_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[3]),
	.prn(vcc));
// synopsys translate_off
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X114_Y36_N23
dffeas \count[2] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[2]~1_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[2]),
	.prn(vcc));
// synopsys translate_off
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X114_Y36_N29
dffeas \count[1] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[1]~2_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[1]),
	.prn(vcc));
// synopsys translate_off
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X114_Y36_N27
dffeas \count[0] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[0]),
	.prn(vcc));
// synopsys translate_off
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X114_Y36_N12
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (!count[0] & (!count[1] & (!count[2] & !count[3])))

	.dataa(count[0]),
	.datab(count[1]),
	.datac(count[2]),
	.datad(count[3]),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h0001;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X114_Y37_N16
cycloneive_lcell_comb \CPUCLK~0 (
// Equation(s):
// \CPUCLK~0_combout  = \CPUCLK~q  $ (\Equal0~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\CPUCLK~q ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\CPUCLK~0_combout ),
	.cout());
// synopsys translate_off
defparam \CPUCLK~0 .lut_mask = 16'h0FF0;
defparam \CPUCLK~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X114_Y36_N0
cycloneive_lcell_comb \count[3]~0 (
// Equation(s):
// \count[3]~0_combout  = count[3] $ (((count[2] & (count[0] & count[1]))))

	.dataa(count[2]),
	.datab(count[0]),
	.datac(count[3]),
	.datad(count[1]),
	.cin(gnd),
	.combout(\count[3]~0_combout ),
	.cout());
// synopsys translate_off
defparam \count[3]~0 .lut_mask = 16'h78F0;
defparam \count[3]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X114_Y36_N22
cycloneive_lcell_comb \count[2]~1 (
// Equation(s):
// \count[2]~1_combout  = count[2] $ (((count[0] & count[1])))

	.dataa(count[0]),
	.datab(gnd),
	.datac(count[2]),
	.datad(count[1]),
	.cin(gnd),
	.combout(\count[2]~1_combout ),
	.cout());
// synopsys translate_off
defparam \count[2]~1 .lut_mask = 16'h5AF0;
defparam \count[2]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X114_Y36_N28
cycloneive_lcell_comb \count[1]~2 (
// Equation(s):
// \count[1]~2_combout  = count[0] $ (count[1])

	.dataa(count[0]),
	.datab(gnd),
	.datac(count[1]),
	.datad(gnd),
	.cin(gnd),
	.combout(\count[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \count[1]~2 .lut_mask = 16'h5A5A;
defparam \count[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X114_Y36_N26
cycloneive_lcell_comb \count~3 (
// Equation(s):
// \count~3_combout  = (!count[0] & ((count[2]) # ((count[1]) # (count[3]))))

	.dataa(count[2]),
	.datab(count[1]),
	.datac(count[0]),
	.datad(count[3]),
	.cin(gnd),
	.combout(\count~3_combout ),
	.cout());
// synopsys translate_off
defparam \count~3 .lut_mask = 16'h0F0E;
defparam \count~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N18
cycloneive_lcell_comb \ramaddr~29_wirecell (
// Equation(s):
// \ramaddr~29_wirecell_combout  = !\ramaddr~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\ramaddr~29_combout ),
	.cin(gnd),
	.combout(\ramaddr~29_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~29_wirecell .lut_mask = 16'h00FF;
defparam \ramaddr~29_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: JTAG_X1_Y37_N0
cycloneive_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

// Location: FF_X35_Y31_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X36_Y31_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y30_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y30_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y30_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y30_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y30_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X38_Y31_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .power_up = "low";
// synopsys translate_on

// Location: FF_X35_Y31_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X35_Y31_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X35_Y31_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y30_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .lut_mask = 16'hEE50;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y30_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .lut_mask = 16'hCC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y31_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .lut_mask = 16'hDF80;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y31_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .lut_mask = 16'h002A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y31_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y31_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .lut_mask = 16'hD8C8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y31_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .lut_mask = 16'h88B8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y31_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X35_Y31_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X35_Y31_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X32_Y31_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4 .lut_mask = 16'h550A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X32_Y31_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6 .lut_mask = 16'h022A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X32_Y31_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~6_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~4_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7 .lut_mask = 16'hF444;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y30_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .lut_mask = 16'hFC0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X35_Y31_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X35_Y31_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .lut_mask = 16'hFFAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y30_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .lut_mask = 16'h44C2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X32_Y31_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .lut_mask = 16'h0500;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X35_Y31_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X35_Y31_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .lut_mask = 16'h5500;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y31_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X33_Y31_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X35_Y31_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X35_Y31_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .lut_mask = 16'hFAFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X33_Y31_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X35_Y31_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y31_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N8
cycloneive_io_ibuf \syif.tbCTRL~input (
	.i(\syif.tbCTRL ),
	.ibar(gnd),
	.o(\syif.tbCTRL~input_o ));
// synopsys translate_off
defparam \syif.tbCTRL~input .bus_hold = "false";
defparam \syif.tbCTRL~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N1
cycloneive_io_ibuf \syif.addr[1]~input (
	.i(\syif.addr [1]),
	.ibar(gnd),
	.o(\syif.addr[1]~input_o ));
// synopsys translate_off
defparam \syif.addr[1]~input .bus_hold = "false";
defparam \syif.addr[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y35_N15
cycloneive_io_ibuf \syif.addr[0]~input (
	.i(\syif.addr [0]),
	.ibar(gnd),
	.o(\syif.addr[0]~input_o ));
// synopsys translate_off
defparam \syif.addr[0]~input .bus_hold = "false";
defparam \syif.addr[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N1
cycloneive_io_ibuf \syif.addr[3]~input (
	.i(\syif.addr [3]),
	.ibar(gnd),
	.o(\syif.addr[3]~input_o ));
// synopsys translate_off
defparam \syif.addr[3]~input .bus_hold = "false";
defparam \syif.addr[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y33_N15
cycloneive_io_ibuf \syif.addr[2]~input (
	.i(\syif.addr [2]),
	.ibar(gnd),
	.o(\syif.addr[2]~input_o ));
// synopsys translate_off
defparam \syif.addr[2]~input .bus_hold = "false";
defparam \syif.addr[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N1
cycloneive_io_ibuf \syif.addr[5]~input (
	.i(\syif.addr [5]),
	.ibar(gnd),
	.o(\syif.addr[5]~input_o ));
// synopsys translate_off
defparam \syif.addr[5]~input .bus_hold = "false";
defparam \syif.addr[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N1
cycloneive_io_ibuf \syif.addr[4]~input (
	.i(\syif.addr [4]),
	.ibar(gnd),
	.o(\syif.addr[4]~input_o ));
// synopsys translate_off
defparam \syif.addr[4]~input .bus_hold = "false";
defparam \syif.addr[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y35_N1
cycloneive_io_ibuf \syif.addr[7]~input (
	.i(\syif.addr [7]),
	.ibar(gnd),
	.o(\syif.addr[7]~input_o ));
// synopsys translate_off
defparam \syif.addr[7]~input .bus_hold = "false";
defparam \syif.addr[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y40_N1
cycloneive_io_ibuf \syif.addr[6]~input (
	.i(\syif.addr [6]),
	.ibar(gnd),
	.o(\syif.addr[6]~input_o ));
// synopsys translate_off
defparam \syif.addr[6]~input .bus_hold = "false";
defparam \syif.addr[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y73_N1
cycloneive_io_ibuf \syif.addr[9]~input (
	.i(\syif.addr [9]),
	.ibar(gnd),
	.o(\syif.addr[9]~input_o ));
// synopsys translate_off
defparam \syif.addr[9]~input .bus_hold = "false";
defparam \syif.addr[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N22
cycloneive_io_ibuf \syif.addr[8]~input (
	.i(\syif.addr [8]),
	.ibar(gnd),
	.o(\syif.addr[8]~input_o ));
// synopsys translate_off
defparam \syif.addr[8]~input .bus_hold = "false";
defparam \syif.addr[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y33_N1
cycloneive_io_ibuf \syif.addr[11]~input (
	.i(\syif.addr [11]),
	.ibar(gnd),
	.o(\syif.addr[11]~input_o ));
// synopsys translate_off
defparam \syif.addr[11]~input .bus_hold = "false";
defparam \syif.addr[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N8
cycloneive_io_ibuf \syif.addr[10]~input (
	.i(\syif.addr [10]),
	.ibar(gnd),
	.o(\syif.addr[10]~input_o ));
// synopsys translate_off
defparam \syif.addr[10]~input .bus_hold = "false";
defparam \syif.addr[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N8
cycloneive_io_ibuf \syif.addr[13]~input (
	.i(\syif.addr [13]),
	.ibar(gnd),
	.o(\syif.addr[13]~input_o ));
// synopsys translate_off
defparam \syif.addr[13]~input .bus_hold = "false";
defparam \syif.addr[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y35_N8
cycloneive_io_ibuf \syif.addr[12]~input (
	.i(\syif.addr [12]),
	.ibar(gnd),
	.o(\syif.addr[12]~input_o ));
// synopsys translate_off
defparam \syif.addr[12]~input .bus_hold = "false";
defparam \syif.addr[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N15
cycloneive_io_ibuf \syif.addr[15]~input (
	.i(\syif.addr [15]),
	.ibar(gnd),
	.o(\syif.addr[15]~input_o ));
// synopsys translate_off
defparam \syif.addr[15]~input .bus_hold = "false";
defparam \syif.addr[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y36_N1
cycloneive_io_ibuf \syif.addr[14]~input (
	.i(\syif.addr [14]),
	.ibar(gnd),
	.o(\syif.addr[14]~input_o ));
// synopsys translate_off
defparam \syif.addr[14]~input .bus_hold = "false";
defparam \syif.addr[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y35_N15
cycloneive_io_ibuf \syif.addr[17]~input (
	.i(\syif.addr [17]),
	.ibar(gnd),
	.o(\syif.addr[17]~input_o ));
// synopsys translate_off
defparam \syif.addr[17]~input .bus_hold = "false";
defparam \syif.addr[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N15
cycloneive_io_ibuf \syif.addr[16]~input (
	.i(\syif.addr [16]),
	.ibar(gnd),
	.o(\syif.addr[16]~input_o ));
// synopsys translate_off
defparam \syif.addr[16]~input .bus_hold = "false";
defparam \syif.addr[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y36_N15
cycloneive_io_ibuf \syif.addr[19]~input (
	.i(\syif.addr [19]),
	.ibar(gnd),
	.o(\syif.addr[19]~input_o ));
// synopsys translate_off
defparam \syif.addr[19]~input .bus_hold = "false";
defparam \syif.addr[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y73_N22
cycloneive_io_ibuf \syif.addr[18]~input (
	.i(\syif.addr [18]),
	.ibar(gnd),
	.o(\syif.addr[18]~input_o ));
// synopsys translate_off
defparam \syif.addr[18]~input .bus_hold = "false";
defparam \syif.addr[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N1
cycloneive_io_ibuf \syif.addr[21]~input (
	.i(\syif.addr [21]),
	.ibar(gnd),
	.o(\syif.addr[21]~input_o ));
// synopsys translate_off
defparam \syif.addr[21]~input .bus_hold = "false";
defparam \syif.addr[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y0_N8
cycloneive_io_ibuf \syif.addr[20]~input (
	.i(\syif.addr [20]),
	.ibar(gnd),
	.o(\syif.addr[20]~input_o ));
// synopsys translate_off
defparam \syif.addr[20]~input .bus_hold = "false";
defparam \syif.addr[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N15
cycloneive_io_ibuf \syif.addr[23]~input (
	.i(\syif.addr [23]),
	.ibar(gnd),
	.o(\syif.addr[23]~input_o ));
// synopsys translate_off
defparam \syif.addr[23]~input .bus_hold = "false";
defparam \syif.addr[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N1
cycloneive_io_ibuf \syif.addr[22]~input (
	.i(\syif.addr [22]),
	.ibar(gnd),
	.o(\syif.addr[22]~input_o ));
// synopsys translate_off
defparam \syif.addr[22]~input .bus_hold = "false";
defparam \syif.addr[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N8
cycloneive_io_ibuf \syif.addr[25]~input (
	.i(\syif.addr [25]),
	.ibar(gnd),
	.o(\syif.addr[25]~input_o ));
// synopsys translate_off
defparam \syif.addr[25]~input .bus_hold = "false";
defparam \syif.addr[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y0_N15
cycloneive_io_ibuf \syif.addr[24]~input (
	.i(\syif.addr [24]),
	.ibar(gnd),
	.o(\syif.addr[24]~input_o ));
// synopsys translate_off
defparam \syif.addr[24]~input .bus_hold = "false";
defparam \syif.addr[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N8
cycloneive_io_ibuf \syif.addr[27]~input (
	.i(\syif.addr [27]),
	.ibar(gnd),
	.o(\syif.addr[27]~input_o ));
// synopsys translate_off
defparam \syif.addr[27]~input .bus_hold = "false";
defparam \syif.addr[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y35_N22
cycloneive_io_ibuf \syif.addr[26]~input (
	.i(\syif.addr [26]),
	.ibar(gnd),
	.o(\syif.addr[26]~input_o ));
// synopsys translate_off
defparam \syif.addr[26]~input .bus_hold = "false";
defparam \syif.addr[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N1
cycloneive_io_ibuf \syif.addr[29]~input (
	.i(\syif.addr [29]),
	.ibar(gnd),
	.o(\syif.addr[29]~input_o ));
// synopsys translate_off
defparam \syif.addr[29]~input .bus_hold = "false";
defparam \syif.addr[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y73_N22
cycloneive_io_ibuf \syif.addr[28]~input (
	.i(\syif.addr [28]),
	.ibar(gnd),
	.o(\syif.addr[28]~input_o ));
// synopsys translate_off
defparam \syif.addr[28]~input .bus_hold = "false";
defparam \syif.addr[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y73_N22
cycloneive_io_ibuf \syif.addr[31]~input (
	.i(\syif.addr [31]),
	.ibar(gnd),
	.o(\syif.addr[31]~input_o ));
// synopsys translate_off
defparam \syif.addr[31]~input .bus_hold = "false";
defparam \syif.addr[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y0_N8
cycloneive_io_ibuf \syif.addr[30]~input (
	.i(\syif.addr [30]),
	.ibar(gnd),
	.o(\syif.addr[30]~input_o ));
// synopsys translate_off
defparam \syif.addr[30]~input .bus_hold = "false";
defparam \syif.addr[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N1
cycloneive_io_ibuf \syif.WEN~input (
	.i(\syif.WEN ),
	.ibar(gnd),
	.o(\syif.WEN~input_o ));
// synopsys translate_off
defparam \syif.WEN~input .bus_hold = "false";
defparam \syif.WEN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y36_N8
cycloneive_io_ibuf \syif.REN~input (
	.i(\syif.REN ),
	.ibar(gnd),
	.o(\syif.REN~input_o ));
// synopsys translate_off
defparam \syif.REN~input .bus_hold = "false";
defparam \syif.REN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N15
cycloneive_io_ibuf \nRST~input (
	.i(nRST),
	.ibar(gnd),
	.o(\nRST~input_o ));
// synopsys translate_off
defparam \nRST~input .bus_hold = "false";
defparam \nRST~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N8
cycloneive_io_ibuf \CLK~input (
	.i(CLK),
	.ibar(gnd),
	.o(\CLK~input_o ));
// synopsys translate_off
defparam \CLK~input .bus_hold = "false";
defparam \CLK~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X47_Y73_N15
cycloneive_io_ibuf \syif.store[0]~input (
	.i(\syif.store [0]),
	.ibar(gnd),
	.o(\syif.store[0]~input_o ));
// synopsys translate_off
defparam \syif.store[0]~input .bus_hold = "false";
defparam \syif.store[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y32_N22
cycloneive_io_ibuf \syif.store[1]~input (
	.i(\syif.store [1]),
	.ibar(gnd),
	.o(\syif.store[1]~input_o ));
// synopsys translate_off
defparam \syif.store[1]~input .bus_hold = "false";
defparam \syif.store[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X47_Y0_N1
cycloneive_io_ibuf \syif.store[2]~input (
	.i(\syif.store [2]),
	.ibar(gnd),
	.o(\syif.store[2]~input_o ));
// synopsys translate_off
defparam \syif.store[2]~input .bus_hold = "false";
defparam \syif.store[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y73_N8
cycloneive_io_ibuf \syif.store[3]~input (
	.i(\syif.store [3]),
	.ibar(gnd),
	.o(\syif.store[3]~input_o ));
// synopsys translate_off
defparam \syif.store[3]~input .bus_hold = "false";
defparam \syif.store[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y73_N1
cycloneive_io_ibuf \syif.store[4]~input (
	.i(\syif.store [4]),
	.ibar(gnd),
	.o(\syif.store[4]~input_o ));
// synopsys translate_off
defparam \syif.store[4]~input .bus_hold = "false";
defparam \syif.store[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N8
cycloneive_io_ibuf \syif.store[5]~input (
	.i(\syif.store [5]),
	.ibar(gnd),
	.o(\syif.store[5]~input_o ));
// synopsys translate_off
defparam \syif.store[5]~input .bus_hold = "false";
defparam \syif.store[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y73_N15
cycloneive_io_ibuf \syif.store[6]~input (
	.i(\syif.store [6]),
	.ibar(gnd),
	.o(\syif.store[6]~input_o ));
// synopsys translate_off
defparam \syif.store[6]~input .bus_hold = "false";
defparam \syif.store[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y73_N1
cycloneive_io_ibuf \syif.store[7]~input (
	.i(\syif.store [7]),
	.ibar(gnd),
	.o(\syif.store[7]~input_o ));
// synopsys translate_off
defparam \syif.store[7]~input .bus_hold = "false";
defparam \syif.store[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y0_N22
cycloneive_io_ibuf \syif.store[8]~input (
	.i(\syif.store [8]),
	.ibar(gnd),
	.o(\syif.store[8]~input_o ));
// synopsys translate_off
defparam \syif.store[8]~input .bus_hold = "false";
defparam \syif.store[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X56_Y0_N8
cycloneive_io_ibuf \syif.store[9]~input (
	.i(\syif.store [9]),
	.ibar(gnd),
	.o(\syif.store[9]~input_o ));
// synopsys translate_off
defparam \syif.store[9]~input .bus_hold = "false";
defparam \syif.store[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y73_N8
cycloneive_io_ibuf \syif.store[10]~input (
	.i(\syif.store [10]),
	.ibar(gnd),
	.o(\syif.store[10]~input_o ));
// synopsys translate_off
defparam \syif.store[10]~input .bus_hold = "false";
defparam \syif.store[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N8
cycloneive_io_ibuf \syif.store[11]~input (
	.i(\syif.store [11]),
	.ibar(gnd),
	.o(\syif.store[11]~input_o ));
// synopsys translate_off
defparam \syif.store[11]~input .bus_hold = "false";
defparam \syif.store[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y0_N15
cycloneive_io_ibuf \syif.store[12]~input (
	.i(\syif.store [12]),
	.ibar(gnd),
	.o(\syif.store[12]~input_o ));
// synopsys translate_off
defparam \syif.store[12]~input .bus_hold = "false";
defparam \syif.store[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N22
cycloneive_io_ibuf \syif.store[13]~input (
	.i(\syif.store [13]),
	.ibar(gnd),
	.o(\syif.store[13]~input_o ));
// synopsys translate_off
defparam \syif.store[13]~input .bus_hold = "false";
defparam \syif.store[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N22
cycloneive_io_ibuf \syif.store[14]~input (
	.i(\syif.store [14]),
	.ibar(gnd),
	.o(\syif.store[14]~input_o ));
// synopsys translate_off
defparam \syif.store[14]~input .bus_hold = "false";
defparam \syif.store[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N15
cycloneive_io_ibuf \syif.store[15]~input (
	.i(\syif.store [15]),
	.ibar(gnd),
	.o(\syif.store[15]~input_o ));
// synopsys translate_off
defparam \syif.store[15]~input .bus_hold = "false";
defparam \syif.store[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y73_N22
cycloneive_io_ibuf \syif.store[16]~input (
	.i(\syif.store [16]),
	.ibar(gnd),
	.o(\syif.store[16]~input_o ));
// synopsys translate_off
defparam \syif.store[16]~input .bus_hold = "false";
defparam \syif.store[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y34_N15
cycloneive_io_ibuf \syif.store[17]~input (
	.i(\syif.store [17]),
	.ibar(gnd),
	.o(\syif.store[17]~input_o ));
// synopsys translate_off
defparam \syif.store[17]~input .bus_hold = "false";
defparam \syif.store[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y73_N1
cycloneive_io_ibuf \syif.store[18]~input (
	.i(\syif.store [18]),
	.ibar(gnd),
	.o(\syif.store[18]~input_o ));
// synopsys translate_off
defparam \syif.store[18]~input .bus_hold = "false";
defparam \syif.store[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N22
cycloneive_io_ibuf \syif.store[19]~input (
	.i(\syif.store [19]),
	.ibar(gnd),
	.o(\syif.store[19]~input_o ));
// synopsys translate_off
defparam \syif.store[19]~input .bus_hold = "false";
defparam \syif.store[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N22
cycloneive_io_ibuf \syif.store[20]~input (
	.i(\syif.store [20]),
	.ibar(gnd),
	.o(\syif.store[20]~input_o ));
// synopsys translate_off
defparam \syif.store[20]~input .bus_hold = "false";
defparam \syif.store[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y0_N22
cycloneive_io_ibuf \syif.store[21]~input (
	.i(\syif.store [21]),
	.ibar(gnd),
	.o(\syif.store[21]~input_o ));
// synopsys translate_off
defparam \syif.store[21]~input .bus_hold = "false";
defparam \syif.store[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N22
cycloneive_io_ibuf \syif.store[22]~input (
	.i(\syif.store [22]),
	.ibar(gnd),
	.o(\syif.store[22]~input_o ));
// synopsys translate_off
defparam \syif.store[22]~input .bus_hold = "false";
defparam \syif.store[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y34_N22
cycloneive_io_ibuf \syif.store[23]~input (
	.i(\syif.store [23]),
	.ibar(gnd),
	.o(\syif.store[23]~input_o ));
// synopsys translate_off
defparam \syif.store[23]~input .bus_hold = "false";
defparam \syif.store[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X56_Y0_N22
cycloneive_io_ibuf \syif.store[24]~input (
	.i(\syif.store [24]),
	.ibar(gnd),
	.o(\syif.store[24]~input_o ));
// synopsys translate_off
defparam \syif.store[24]~input .bus_hold = "false";
defparam \syif.store[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X56_Y0_N1
cycloneive_io_ibuf \syif.store[25]~input (
	.i(\syif.store [25]),
	.ibar(gnd),
	.o(\syif.store[25]~input_o ));
// synopsys translate_off
defparam \syif.store[25]~input .bus_hold = "false";
defparam \syif.store[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y34_N15
cycloneive_io_ibuf \syif.store[26]~input (
	.i(\syif.store [26]),
	.ibar(gnd),
	.o(\syif.store[26]~input_o ));
// synopsys translate_off
defparam \syif.store[26]~input .bus_hold = "false";
defparam \syif.store[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y0_N1
cycloneive_io_ibuf \syif.store[27]~input (
	.i(\syif.store [27]),
	.ibar(gnd),
	.o(\syif.store[27]~input_o ));
// synopsys translate_off
defparam \syif.store[27]~input .bus_hold = "false";
defparam \syif.store[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N22
cycloneive_io_ibuf \syif.store[28]~input (
	.i(\syif.store [28]),
	.ibar(gnd),
	.o(\syif.store[28]~input_o ));
// synopsys translate_off
defparam \syif.store[28]~input .bus_hold = "false";
defparam \syif.store[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N1
cycloneive_io_ibuf \syif.store[29]~input (
	.i(\syif.store [29]),
	.ibar(gnd),
	.o(\syif.store[29]~input_o ));
// synopsys translate_off
defparam \syif.store[29]~input .bus_hold = "false";
defparam \syif.store[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y73_N8
cycloneive_io_ibuf \syif.store[30]~input (
	.i(\syif.store [30]),
	.ibar(gnd),
	.o(\syif.store[30]~input_o ));
// synopsys translate_off
defparam \syif.store[30]~input .bus_hold = "false";
defparam \syif.store[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y0_N1
cycloneive_io_ibuf \syif.store[31]~input (
	.i(\syif.store [31]),
	.ibar(gnd),
	.o(\syif.store[31]~input_o ));
// synopsys translate_off
defparam \syif.store[31]~input .bus_hold = "false";
defparam \syif.store[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: CLKCTRL_G0
cycloneive_clkctrl \altera_internal_jtag~TCKUTAPclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\altera_internal_jtag~TCKUTAP }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ));
// synopsys translate_off
defparam \altera_internal_jtag~TCKUTAPclkctrl .clock_type = "global clock";
defparam \altera_internal_jtag~TCKUTAPclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G5
cycloneive_clkctrl \CPUCLK~clkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CPUCLK~q }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CPUCLK~clkctrl_outclk ));
// synopsys translate_off
defparam \CPUCLK~clkctrl .clock_type = "global clock";
defparam \CPUCLK~clkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G1
cycloneive_clkctrl \nRST~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\nRST~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\nRST~inputclkctrl_outclk ));
// synopsys translate_off
defparam \nRST~inputclkctrl .clock_type = "global clock";
defparam \nRST~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G2
cycloneive_clkctrl \CLK~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CLK~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CLK~inputclkctrl_outclk ));
// synopsys translate_off
defparam \CLK~inputclkctrl .clock_type = "global clock";
defparam \CLK~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: LCCOMB_X40_Y30_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y30_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y30_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X33_Y31_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder .lut_mask = 16'hF0F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X33_Y31_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOOBUF_X0_Y32_N16
cycloneive_io_obuf \syif.halt~output (
	.i(\CPU|DP|dpif.halt~q ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.halt ),
	.obar());
// synopsys translate_off
defparam \syif.halt~output .bus_hold = "false";
defparam \syif.halt~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y73_N23
cycloneive_io_obuf \syif.load[0]~output (
	.i(\RAM|ramif.ramload[0]~12_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [0]),
	.obar());
// synopsys translate_off
defparam \syif.load[0]~output .bus_hold = "false";
defparam \syif.load[0]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X40_Y73_N9
cycloneive_io_obuf \syif.load[1]~output (
	.i(\RAM|ramif.ramload[1]~13_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [1]),
	.obar());
// synopsys translate_off
defparam \syif.load[1]~output .bus_hold = "false";
defparam \syif.load[1]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N23
cycloneive_io_obuf \syif.load[2]~output (
	.i(\RAM|ramif.ramload[2]~14_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [2]),
	.obar());
// synopsys translate_off
defparam \syif.load[2]~output .bus_hold = "false";
defparam \syif.load[2]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y34_N2
cycloneive_io_obuf \syif.load[3]~output (
	.i(\RAM|ramif.ramload[3]~15_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [3]),
	.obar());
// synopsys translate_off
defparam \syif.load[3]~output .bus_hold = "false";
defparam \syif.load[3]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y34_N9
cycloneive_io_obuf \syif.load[4]~output (
	.i(\RAM|ramif.ramload[4]~16_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [4]),
	.obar());
// synopsys translate_off
defparam \syif.load[4]~output .bus_hold = "false";
defparam \syif.load[4]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y73_N2
cycloneive_io_obuf \syif.load[5]~output (
	.i(\RAM|ramif.ramload[5]~17_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [5]),
	.obar());
// synopsys translate_off
defparam \syif.load[5]~output .bus_hold = "false";
defparam \syif.load[5]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y0_N16
cycloneive_io_obuf \syif.load[6]~output (
	.i(\RAM|ramif.ramload[6]~18_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [6]),
	.obar());
// synopsys translate_off
defparam \syif.load[6]~output .bus_hold = "false";
defparam \syif.load[6]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X58_Y73_N23
cycloneive_io_obuf \syif.load[7]~output (
	.i(\RAM|ramif.ramload[7]~19_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [7]),
	.obar());
// synopsys translate_off
defparam \syif.load[7]~output .bus_hold = "false";
defparam \syif.load[7]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X47_Y73_N2
cycloneive_io_obuf \syif.load[8]~output (
	.i(\RAM|ramif.ramload[8]~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [8]),
	.obar());
// synopsys translate_off
defparam \syif.load[8]~output .bus_hold = "false";
defparam \syif.load[8]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X42_Y73_N9
cycloneive_io_obuf \syif.load[9]~output (
	.i(\RAM|ramif.ramload[9]~21_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [9]),
	.obar());
// synopsys translate_off
defparam \syif.load[9]~output .bus_hold = "false";
defparam \syif.load[9]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X49_Y0_N2
cycloneive_io_obuf \syif.load[10]~output (
	.i(\RAM|ramif.ramload[10]~22_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [10]),
	.obar());
// synopsys translate_off
defparam \syif.load[10]~output .bus_hold = "false";
defparam \syif.load[10]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y34_N23
cycloneive_io_obuf \syif.load[11]~output (
	.i(\RAM|ramif.ramload[11]~23_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [11]),
	.obar());
// synopsys translate_off
defparam \syif.load[11]~output .bus_hold = "false";
defparam \syif.load[11]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X47_Y0_N9
cycloneive_io_obuf \syif.load[12]~output (
	.i(\RAM|ramif.ramload[12]~24_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [12]),
	.obar());
// synopsys translate_off
defparam \syif.load[12]~output .bus_hold = "false";
defparam \syif.load[12]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N2
cycloneive_io_obuf \syif.load[13]~output (
	.i(\RAM|ramif.ramload[13]~25_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [13]),
	.obar());
// synopsys translate_off
defparam \syif.load[13]~output .bus_hold = "false";
defparam \syif.load[13]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X49_Y0_N9
cycloneive_io_obuf \syif.load[14]~output (
	.i(\RAM|ramif.ramload[14]~26_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [14]),
	.obar());
// synopsys translate_off
defparam \syif.load[14]~output .bus_hold = "false";
defparam \syif.load[14]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X38_Y73_N9
cycloneive_io_obuf \syif.load[15]~output (
	.i(\RAM|ramif.ramload[15]~27_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [15]),
	.obar());
// synopsys translate_off
defparam \syif.load[15]~output .bus_hold = "false";
defparam \syif.load[15]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y0_N16
cycloneive_io_obuf \syif.load[16]~output (
	.i(\RAM|ramif.ramload[16]~28_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [16]),
	.obar());
// synopsys translate_off
defparam \syif.load[16]~output .bus_hold = "false";
defparam \syif.load[16]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N16
cycloneive_io_obuf \syif.load[17]~output (
	.i(\RAM|ramif.ramload[17]~29_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [17]),
	.obar());
// synopsys translate_off
defparam \syif.load[17]~output .bus_hold = "false";
defparam \syif.load[17]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y32_N9
cycloneive_io_obuf \syif.load[18]~output (
	.i(\RAM|ramif.ramload[18]~30_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [18]),
	.obar());
// synopsys translate_off
defparam \syif.load[18]~output .bus_hold = "false";
defparam \syif.load[18]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y73_N9
cycloneive_io_obuf \syif.load[19]~output (
	.i(\RAM|ramif.ramload[19]~31_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [19]),
	.obar());
// synopsys translate_off
defparam \syif.load[19]~output .bus_hold = "false";
defparam \syif.load[19]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y41_N9
cycloneive_io_obuf \syif.load[20]~output (
	.i(\RAM|ramif.ramload[20]~32_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [20]),
	.obar());
// synopsys translate_off
defparam \syif.load[20]~output .bus_hold = "false";
defparam \syif.load[20]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y0_N16
cycloneive_io_obuf \syif.load[21]~output (
	.i(\RAM|ramif.ramload[21]~33_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [21]),
	.obar());
// synopsys translate_off
defparam \syif.load[21]~output .bus_hold = "false";
defparam \syif.load[21]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N16
cycloneive_io_obuf \syif.load[22]~output (
	.i(\RAM|ramif.ramload[22]~34_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [22]),
	.obar());
// synopsys translate_off
defparam \syif.load[22]~output .bus_hold = "false";
defparam \syif.load[22]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y73_N16
cycloneive_io_obuf \syif.load[23]~output (
	.i(\RAM|ramif.ramload[23]~35_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [23]),
	.obar());
// synopsys translate_off
defparam \syif.load[23]~output .bus_hold = "false";
defparam \syif.load[23]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y73_N16
cycloneive_io_obuf \syif.load[24]~output (
	.i(\RAM|ramif.ramload[24]~36_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [24]),
	.obar());
// synopsys translate_off
defparam \syif.load[24]~output .bus_hold = "false";
defparam \syif.load[24]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y73_N16
cycloneive_io_obuf \syif.load[25]~output (
	.i(\RAM|ramif.ramload[25]~37_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [25]),
	.obar());
// synopsys translate_off
defparam \syif.load[25]~output .bus_hold = "false";
defparam \syif.load[25]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X58_Y73_N9
cycloneive_io_obuf \syif.load[26]~output (
	.i(\RAM|ramif.ramload[26]~44_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [26]),
	.obar());
// synopsys translate_off
defparam \syif.load[26]~output .bus_hold = "false";
defparam \syif.load[26]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y33_N9
cycloneive_io_obuf \syif.load[27]~output (
	.i(\RAM|ramif.ramload[27]~45_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [27]),
	.obar());
// synopsys translate_off
defparam \syif.load[27]~output .bus_hold = "false";
defparam \syif.load[27]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N16
cycloneive_io_obuf \syif.load[28]~output (
	.i(\RAM|ramif.ramload[28]~46_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [28]),
	.obar());
// synopsys translate_off
defparam \syif.load[28]~output .bus_hold = "false";
defparam \syif.load[28]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X67_Y73_N9
cycloneive_io_obuf \syif.load[29]~output (
	.i(\RAM|ramif.ramload[29]~47_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [29]),
	.obar());
// synopsys translate_off
defparam \syif.load[29]~output .bus_hold = "false";
defparam \syif.load[29]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X42_Y0_N23
cycloneive_io_obuf \syif.load[30]~output (
	.i(\RAM|ramif.ramload[30]~48_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [30]),
	.obar());
// synopsys translate_off
defparam \syif.load[30]~output .bus_hold = "false";
defparam \syif.load[30]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y41_N2
cycloneive_io_obuf \syif.load[31]~output (
	.i(\RAM|ramif.ramload[31]~49_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [31]),
	.obar());
// synopsys translate_off
defparam \syif.load[31]~output .bus_hold = "false";
defparam \syif.load[31]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y37_N1
cycloneive_io_obuf \altera_reserved_tdo~output (
	.i(\altera_internal_jtag~TDO ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(altera_reserved_tdo),
	.obar());
// synopsys translate_off
defparam \altera_reserved_tdo~output .bus_hold = "false";
defparam \altera_reserved_tdo~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOIBUF_X0_Y38_N1
cycloneive_io_ibuf \altera_reserved_tms~input (
	.i(altera_reserved_tms),
	.ibar(gnd),
	.o(\altera_reserved_tms~input_o ));
// synopsys translate_off
defparam \altera_reserved_tms~input .bus_hold = "false";
defparam \altera_reserved_tms~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y39_N1
cycloneive_io_ibuf \altera_reserved_tck~input (
	.i(altera_reserved_tck),
	.ibar(gnd),
	.o(\altera_reserved_tck~input_o ));
// synopsys translate_off
defparam \altera_reserved_tck~input .bus_hold = "false";
defparam \altera_reserved_tck~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y40_N1
cycloneive_io_ibuf \altera_reserved_tdi~input (
	.i(altera_reserved_tdi),
	.ibar(gnd),
	.o(\altera_reserved_tdi~input_o ));
// synopsys translate_off
defparam \altera_reserved_tdi~input .bus_hold = "false";
defparam \altera_reserved_tdi~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X35_Y31_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .lut_mask = 16'hFEFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X35_Y31_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y31_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .lut_mask = 16'hAA88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y31_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X35_Y31_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X35_Y31_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X35_Y31_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X35_Y31_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X35_Y31_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .lut_mask = 16'hF0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X35_Y31_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y31_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X36_Y31_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y31_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .lut_mask = 16'h5AF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X36_Y31_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y31_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y31_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X36_Y31_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y31_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .lut_mask = 16'h5575;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X36_Y31_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X35_Y31_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X35_Y31_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y31_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .lut_mask = 16'hF0E0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y31_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y31_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y31_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y30_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .lut_mask = 16'h3000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y31_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X35_Y31_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .lut_mask = 16'hA0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X35_Y31_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X35_Y31_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .lut_mask = 16'hFFFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X35_Y31_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X39_Y31_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X39_Y31_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y31_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y31_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y31_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y31_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y31_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y31_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y31_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y31_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y31_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y31_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y31_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .lut_mask = 16'h0F0F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y31_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y31_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .lut_mask = 16'h0010;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y31_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .lut_mask = 16'h0001;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y31_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y31_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X39_Y31_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .lut_mask = 16'h0040;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X35_Y31_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .lut_mask = 16'hC8C8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X35_Y31_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X35_Y31_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hF0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y31_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y31_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .lut_mask = 16'hE000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y30_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 .lut_mask = 16'h44F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y31_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .lut_mask = 16'hFC30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y31_N4
cycloneive_lcell_comb \~QIC_CREATED_GND~I (
// Equation(s):
// \~QIC_CREATED_GND~I_combout  = GND

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~QIC_CREATED_GND~I_combout ),
	.cout());
// synopsys translate_off
defparam \~QIC_CREATED_GND~I .lut_mask = 16'h0000;
defparam \~QIC_CREATED_GND~I .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y31_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.asdata(\~QIC_CREATED_GND~I_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y30_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 .lut_mask = 16'hF078;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X36_Y30_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y30_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .lut_mask = 16'h2000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X38_Y30_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y30_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y30_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 .lut_mask = 16'h44F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y30_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X38_Y31_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X38_Y31_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .power_up = "low";
// synopsys translate_on

// Location: FF_X36_Y30_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y30_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y31_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.datac(gnd),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .lut_mask = 16'hEE44;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y30_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .lut_mask = 16'hFC30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y30_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .lut_mask = 16'hB800;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y30_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y30_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .lut_mask = 16'hCFC0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y31_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y30_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .lut_mask = 16'hF3C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y30_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y30_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .lut_mask = 16'hFC30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y30_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y30_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .lut_mask = 16'hFC30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X40_Y30_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y31_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .lut_mask = 16'hCCF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X36_Y31_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X34_Y30_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h55AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X34_Y30_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .lut_mask = 16'h3C3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X34_Y30_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .lut_mask = 16'hC30C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X34_Y30_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h5A5F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X33_Y31_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y31_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .lut_mask = 16'h4000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X39_Y31_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X34_Y31_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .lut_mask = 16'hDCCC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X34_Y30_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X34_Y30_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X33_Y30_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .lut_mask = 16'hFFFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X34_Y30_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .lut_mask = 16'hC3C3;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X34_Y30_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X34_Y30_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .lut_mask = 16'hBA30;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X34_Y30_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X34_Y30_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X34_Y30_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .lut_mask = 16'hF0F1;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X34_Y30_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .lut_mask = 16'h0100;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X34_Y30_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .lut_mask = 16'h0054;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X34_Y30_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .lut_mask = 16'h3320;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X34_Y31_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .lut_mask = 16'hFCEC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X34_Y30_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X34_Y30_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .lut_mask = 16'hCECC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X34_Y30_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X34_Y30_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .lut_mask = 16'hBA10;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X34_Y30_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .lut_mask = 16'h50F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X34_Y30_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X34_Y30_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .lut_mask = 16'h8801;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X34_Y30_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .lut_mask = 16'h0100;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X34_Y30_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .lut_mask = 16'hFF08;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X34_Y30_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y30_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .lut_mask = 16'hCBC8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y30_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 (
	.dataa(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .lut_mask = 16'hB8B8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y30_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .lut_mask = 16'hEE04;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y30_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .lut_mask = 16'hFAAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y31_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y30_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .lut_mask = 16'h4000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y31_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .lut_mask = 16'h00A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X36_Y31_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y31_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder .lut_mask = 16'hF0F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X36_Y31_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y31_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X36_Y31_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y31_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X36_Y31_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X33_Y31_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder .lut_mask = 16'hF0F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y31_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .lut_mask = 16'h0040;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X33_Y31_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X31_Y31_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 .lut_mask = 16'h33CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X32_Y31_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .lut_mask = 16'h0055;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X31_Y31_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~12 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~14 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13 .lut_mask = 16'hC303;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X31_Y31_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~14 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 .lut_mask = 16'h3C3C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X34_Y31_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 .lut_mask = 16'hECA0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X31_Y31_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X32_Y31_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5 .lut_mask = 16'h000F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X31_Y31_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~8 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7 .lut_mask = 16'hA505;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X31_Y31_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X32_Y31_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 .lut_mask = 16'hAAEA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X31_Y31_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X31_Y31_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~8 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~12 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11 .lut_mask = 16'h5AAF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X31_Y31_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X32_Y31_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 .lut_mask = 16'hAA00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X32_Y31_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~9 .lut_mask = 16'h8000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X33_Y31_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~7_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .lut_mask = 16'hCCAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X32_Y31_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X31_Y31_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~9_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~10_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X32_Y31_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12 .lut_mask = 16'h3075;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X32_Y31_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~12_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 .lut_mask = 16'hF5A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X32_Y31_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 .lut_mask = 16'h70F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X33_Y31_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~13_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .lut_mask = 16'hAACC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X32_Y31_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 .lut_mask = 16'h0802;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X32_Y31_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~5_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 .lut_mask = 16'hDCED;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X33_Y31_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .lut_mask = 16'hAACC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X32_Y31_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 .lut_mask = 16'h3BCE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X32_Y31_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .lut_mask = 16'h8F80;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X33_Y31_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .lut_mask = 16'hAACC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X33_Y31_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .lut_mask = 16'h33FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X33_Y31_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .lut_mask = 16'hFC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X33_Y31_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X33_Y31_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X33_Y31_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X33_Y31_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y30_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .lut_mask = 16'h1D3D;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X35_Y31_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .lut_mask = 16'hFAFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X36_Y30_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo (
	.clk(!\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X36_Y30_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y9_N0
cycloneive_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X36_Y31_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X39_Y31_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module ram (
	is_in_use_reg,
	ramaddr,
	ramaddr1,
	ramaddr2,
	ramaddr3,
	ramaddr4,
	ramaddr5,
	ramaddr6,
	ramaddr7,
	ramaddr8,
	ramaddr9,
	ramaddr10,
	ramaddr11,
	ramaddr12,
	ramaddr13,
	ramaddr14,
	ramaddr15,
	\ramif.ramaddr ,
	ramaddr16,
	ramaddr17,
	ramaddr18,
	ramaddr19,
	ramaddr20,
	ramaddr21,
	ramaddr22,
	ramaddr23,
	ramaddr24,
	ramaddr25,
	ramaddr26,
	ramaddr27,
	ramWEN,
	ramREN,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	ramstore,
	ramstore1,
	ramstore2,
	ramstore3,
	ramstore4,
	ramstore5,
	ramstore6,
	ramstore7,
	ramstore8,
	ramstore9,
	ramstore10,
	ramstore11,
	ramstore12,
	ramstore13,
	ramstore14,
	ramstore15,
	ramstore16,
	ramstore17,
	ramstore18,
	ramstore19,
	ramstore20,
	ramstore21,
	ramstore22,
	ramstore23,
	ramstore24,
	ramstore25,
	ramstore26,
	ramstore27,
	ramstore28,
	ramstore29,
	ramstore30,
	ramstore31,
	ramiframload_261,
	ramiframload_271,
	ramiframload_281,
	ramiframload_291,
	ramiframload_301,
	ramiframload_311,
	ramaddr28,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	nRST,
	altera_internal_jtag1,
	nRST1,
	CLK,
	devpor,
	devclrn,
	devoe);
output 	is_in_use_reg;
input 	ramaddr;
input 	ramaddr1;
input 	ramaddr2;
input 	ramaddr3;
input 	ramaddr4;
input 	ramaddr5;
input 	ramaddr6;
input 	ramaddr7;
input 	ramaddr8;
input 	ramaddr9;
input 	ramaddr10;
input 	ramaddr11;
input 	ramaddr12;
input 	ramaddr13;
input 	ramaddr14;
input 	ramaddr15;
input 	[31:0] \ramif.ramaddr ;
input 	ramaddr16;
input 	ramaddr17;
input 	ramaddr18;
input 	ramaddr19;
input 	ramaddr20;
input 	ramaddr21;
input 	ramaddr22;
input 	ramaddr23;
input 	ramaddr24;
input 	ramaddr25;
input 	ramaddr26;
input 	ramaddr27;
input 	ramWEN;
input 	ramREN;
output 	always1;
output 	ramiframload_0;
output 	ramiframload_1;
output 	ramiframload_2;
output 	ramiframload_3;
output 	ramiframload_4;
output 	ramiframload_5;
output 	ramiframload_6;
output 	ramiframload_7;
output 	ramiframload_8;
output 	ramiframload_9;
output 	ramiframload_10;
output 	ramiframload_11;
output 	ramiframload_12;
output 	ramiframload_13;
output 	ramiframload_14;
output 	ramiframload_15;
output 	ramiframload_16;
output 	ramiframload_17;
output 	ramiframload_18;
output 	ramiframload_19;
output 	ramiframload_20;
output 	ramiframload_21;
output 	ramiframload_22;
output 	ramiframload_23;
output 	ramiframload_24;
output 	ramiframload_25;
output 	ramiframload_26;
output 	ramiframload_27;
output 	ramiframload_28;
output 	ramiframload_29;
output 	ramiframload_30;
output 	ramiframload_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	ramstore;
input 	ramstore1;
input 	ramstore2;
input 	ramstore3;
input 	ramstore4;
input 	ramstore5;
input 	ramstore6;
input 	ramstore7;
input 	ramstore8;
input 	ramstore9;
input 	ramstore10;
input 	ramstore11;
input 	ramstore12;
input 	ramstore13;
input 	ramstore14;
input 	ramstore15;
input 	ramstore16;
input 	ramstore17;
input 	ramstore18;
input 	ramstore19;
input 	ramstore20;
input 	ramstore21;
input 	ramstore22;
input 	ramstore23;
input 	ramstore24;
input 	ramstore25;
input 	ramstore26;
input 	ramstore27;
input 	ramstore28;
input 	ramstore29;
input 	ramstore30;
input 	ramstore31;
output 	ramiframload_261;
output 	ramiframload_271;
output 	ramiframload_281;
output 	ramiframload_291;
output 	ramiframload_301;
output 	ramiframload_311;
input 	ramaddr28;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	nRST;
input 	altera_internal_jtag1;
input 	nRST1;
input 	CLK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ;
wire \always0~1_combout ;
wire \always0~6_combout ;
wire \always0~11_combout ;
wire \always0~16_combout ;
wire \always0~22_combout ;
wire \addr[27]~feeder_combout ;
wire \always0~5_combout ;
wire \always0~7_combout ;
wire \always0~8_combout ;
wire \always0~9_combout ;
wire \always0~0_combout ;
wire \always0~2_combout ;
wire \always0~3_combout ;
wire \always0~4_combout ;
wire \always0~10_combout ;
wire \always0~19_combout ;
wire \always0~18_combout ;
wire \always0~17_combout ;
wire \always0~20_combout ;
wire \always0~12_combout ;
wire \always0~14_combout ;
wire \always0~13_combout ;
wire \always0~15_combout ;
wire \always0~21_combout ;
wire \always0~23_combout ;
wire \count[0]~3_combout ;
wire \count[1]~2_combout ;
wire \Add0~1_combout ;
wire \count[2]~1_combout ;
wire \Add0~0_combout ;
wire \count[3]~0_combout ;
wire \LessThan1~0_combout ;
wire [1:0] en;
wire [3:0] count;
wire [31:0] addr;
wire [0:0] \altsyncram_component|auto_generated|altsyncram1|address_reg_a ;


altsyncram_1 altsyncram_component(
	.ram_block3a32(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.ram_block3a0(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.ram_block3a33(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.ram_block3a1(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.ram_block3a34(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.ram_block3a2(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.ram_block3a35(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.ram_block3a3(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.ram_block3a36(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.ram_block3a4(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.ram_block3a37(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.ram_block3a5(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.ram_block3a38(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.ram_block3a6(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.ram_block3a39(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.ram_block3a7(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.ram_block3a40(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.ram_block3a8(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.ram_block3a41(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.ram_block3a9(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.ram_block3a42(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.ram_block3a10(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.ram_block3a43(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.ram_block3a11(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.ram_block3a44(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.ram_block3a12(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.ram_block3a45(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.ram_block3a13(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.ram_block3a46(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.ram_block3a14(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.ram_block3a47(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.ram_block3a15(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.ram_block3a48(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.ram_block3a16(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.ram_block3a49(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.ram_block3a17(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.ram_block3a50(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.ram_block3a18(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.ram_block3a51(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.ram_block3a19(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.ram_block3a52(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.ram_block3a20(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.ram_block3a53(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.ram_block3a21(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.ram_block3a54(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.ram_block3a22(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.ram_block3a55(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.ram_block3a23(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.ram_block3a56(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.ram_block3a24(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.ram_block3a57(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.ram_block3a25(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.ram_block3a58(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.ram_block3a26(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.ram_block3a59(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.ram_block3a27(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.ram_block3a60(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.ram_block3a28(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.ram_block3a61(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.ram_block3a29(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.ram_block3a62(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.ram_block3a30(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.ram_block3a63(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.ram_block3a31(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.address_a({gnd,ramaddr15,ramaddr12,ramaddr13,ramaddr10,ramaddr11,ramaddr8,ramaddr9,ramaddr6,ramaddr7,ramaddr4,ramaddr5,ramaddr2,ramaddr3}),
	.ramaddr(ramaddr14),
	.ramWEN(ramWEN),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.data_a({ramstore31,ramstore30,ramstore29,ramstore28,ramstore27,ramstore26,ramstore25,ramstore24,ramstore23,ramstore22,ramstore21,ramstore20,ramstore19,ramstore18,ramstore17,ramstore16,ramstore15,ramstore14,ramstore13,ramstore12,ramstore11,ramstore10,ramstore9,ramstore8,ramstore7,ramstore6,
ramstore5,ramstore4,ramstore3,ramstore2,ramstore1,ramstore}),
	.ramaddr1(ramaddr28),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(CLK),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: FF_X55_Y36_N19
dffeas \addr[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[1]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[1] .is_wysiwyg = "true";
defparam \addr[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N17
dffeas \addr[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr3),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[2]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[2] .is_wysiwyg = "true";
defparam \addr[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N3
dffeas \addr[3] (
	.clk(CLK),
	.d(ramaddr2),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[3]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[3] .is_wysiwyg = "true";
defparam \addr[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N16
cycloneive_lcell_comb \always0~1 (
// Equation(s):
// \always0~1_combout  = (addr[3] & (\ramaddr~5_combout  & (addr[2] $ (!\ramaddr~7_combout )))) # (!addr[3] & (!\ramaddr~5_combout  & (addr[2] $ (!\ramaddr~7_combout ))))

	.dataa(addr[3]),
	.datab(ramaddr2),
	.datac(addr[2]),
	.datad(ramaddr3),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
// synopsys translate_off
defparam \always0~1 .lut_mask = 16'h9009;
defparam \always0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N7
dffeas \addr[5] (
	.clk(CLK),
	.d(ramaddr4),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[5]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[5] .is_wysiwyg = "true";
defparam \addr[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N17
dffeas \addr[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr11),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[10]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[10] .is_wysiwyg = "true";
defparam \addr[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N31
dffeas \addr[11] (
	.clk(CLK),
	.d(ramaddr10),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[11]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[11] .is_wysiwyg = "true";
defparam \addr[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N16
cycloneive_lcell_comb \always0~6 (
// Equation(s):
// \always0~6_combout  = (\ramaddr~21_combout  & (addr[11] & (\ramaddr~23_combout  $ (!addr[10])))) # (!\ramaddr~21_combout  & (!addr[11] & (\ramaddr~23_combout  $ (!addr[10]))))

	.dataa(ramaddr10),
	.datab(ramaddr11),
	.datac(addr[10]),
	.datad(addr[11]),
	.cin(gnd),
	.combout(\always0~6_combout ),
	.cout());
// synopsys translate_off
defparam \always0~6 .lut_mask = 16'h8241;
defparam \always0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N27
dffeas \addr[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr28),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[15]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[15] .is_wysiwyg = "true";
defparam \addr[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N13
dffeas \addr[16] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr16),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[16]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[16] .is_wysiwyg = "true";
defparam \addr[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N11
dffeas \addr[17] (
	.clk(CLK),
	.d(\ramif.ramaddr [17]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[17]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[17] .is_wysiwyg = "true";
defparam \addr[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N12
cycloneive_lcell_comb \always0~11 (
// Equation(s):
// \always0~11_combout  = (addr[17] & (\ramaddr~33_combout  & (\ramaddr~35_combout  $ (!addr[16])))) # (!addr[17] & (!\ramaddr~33_combout  & (\ramaddr~35_combout  $ (!addr[16]))))

	.dataa(addr[17]),
	.datab(ramaddr16),
	.datac(addr[16]),
	.datad(\ramif.ramaddr [17]),
	.cin(gnd),
	.combout(\always0~11_combout ),
	.cout());
// synopsys translate_off
defparam \always0~11 .lut_mask = 16'h8241;
defparam \always0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N29
dffeas \addr[19] (
	.clk(CLK),
	.d(\ramif.ramaddr [19]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[19]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[19] .is_wysiwyg = "true";
defparam \addr[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N17
dffeas \addr[21] (
	.clk(CLK),
	.d(\ramif.ramaddr [21]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[21]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[21] .is_wysiwyg = "true";
defparam \addr[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N11
dffeas \addr[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr21),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[24]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[24] .is_wysiwyg = "true";
defparam \addr[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N13
dffeas \addr[25] (
	.clk(CLK),
	.d(\ramif.ramaddr [25]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[25]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[25] .is_wysiwyg = "true";
defparam \addr[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N10
cycloneive_lcell_comb \always0~16 (
// Equation(s):
// \always0~16_combout  = (\ramaddr~51_combout  & (addr[24] & (addr[25] $ (!\ramaddr~49_combout )))) # (!\ramaddr~51_combout  & (!addr[24] & (addr[25] $ (!\ramaddr~49_combout ))))

	.dataa(ramaddr21),
	.datab(addr[25]),
	.datac(addr[24]),
	.datad(\ramif.ramaddr [25]),
	.cin(gnd),
	.combout(\always0~16_combout ),
	.cout());
// synopsys translate_off
defparam \always0~16 .lut_mask = 16'h8421;
defparam \always0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N5
dffeas \addr[27] (
	.clk(CLK),
	.d(\addr[27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[27]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[27] .is_wysiwyg = "true";
defparam \addr[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N7
dffeas \addr[29] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr24),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[29]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[29] .is_wysiwyg = "true";
defparam \addr[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y37_N7
dffeas \addr[31] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr26),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[31]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[31] .is_wysiwyg = "true";
defparam \addr[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N3
dffeas \en[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramREN),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[1]),
	.prn(vcc));
// synopsys translate_off
defparam \en[1] .is_wysiwyg = "true";
defparam \en[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N31
dffeas \en[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramWEN),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[0]),
	.prn(vcc));
// synopsys translate_off
defparam \en[0] .is_wysiwyg = "true";
defparam \en[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N30
cycloneive_lcell_comb \always0~22 (
// Equation(s):
// \always0~22_combout  = (\ramWEN~0_combout  & ((en[1] $ (\ramREN~0_combout )) # (!en[0]))) # (!\ramWEN~0_combout  & ((en[0]) # (en[1] $ (\ramREN~0_combout ))))

	.dataa(ramWEN),
	.datab(en[1]),
	.datac(en[0]),
	.datad(ramREN),
	.cin(gnd),
	.combout(\always0~22_combout ),
	.cout());
// synopsys translate_off
defparam \always0~22 .lut_mask = 16'h7BDE;
defparam \always0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N4
cycloneive_lcell_comb \addr[27]~feeder (
// Equation(s):
// \addr[27]~feeder_combout  = \ramaddr~53_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr22),
	.cin(gnd),
	.combout(\addr[27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[27]~feeder .lut_mask = 16'hFF00;
defparam \addr[27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N16
cycloneive_lcell_comb \always1~0 (
// Equation(s):
// always1 = ((\LessThan1~0_combout  & (\always0~21_combout  & \always0~10_combout ))) # (!\nRST~input_o )

	.dataa(\LessThan1~0_combout ),
	.datab(nRST),
	.datac(\always0~21_combout ),
	.datad(\always0~10_combout ),
	.cin(gnd),
	.combout(always1),
	.cout());
// synopsys translate_off
defparam \always1~0 .lut_mask = 16'hB333;
defparam \always1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N12
cycloneive_lcell_comb \ramif.ramload[0]~12 (
// Equation(s):
// ramiframload_0 = ((address_reg_a_0 & ((ram_block3a321))) # (!address_reg_a_0 & (ram_block3a01))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_0),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[0]~12 .lut_mask = 16'hE4FF;
defparam \ramif.ramload[0]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N8
cycloneive_lcell_comb \ramif.ramload[1]~13 (
// Equation(s):
// ramiframload_1 = (always1 & ((address_reg_a_0 & ((ram_block3a331))) # (!address_reg_a_0 & (ram_block3a110))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_1),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[1]~13 .lut_mask = 16'hE200;
defparam \ramif.ramload[1]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N12
cycloneive_lcell_comb \ramif.ramload[2]~14 (
// Equation(s):
// ramiframload_2 = (always1 & ((address_reg_a_0 & ((ram_block3a341))) # (!address_reg_a_0 & (ram_block3a210))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_2),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[2]~14 .lut_mask = 16'hE200;
defparam \ramif.ramload[2]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N6
cycloneive_lcell_comb \ramif.ramload[3]~15 (
// Equation(s):
// ramiframload_3 = (always1 & ((address_reg_a_0 & ((ram_block3a351))) # (!address_reg_a_0 & (ram_block3a310))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_3),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[3]~15 .lut_mask = 16'hE200;
defparam \ramif.ramload[3]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N4
cycloneive_lcell_comb \ramif.ramload[4]~16 (
// Equation(s):
// ramiframload_4 = ((address_reg_a_0 & ((ram_block3a361))) # (!address_reg_a_0 & (ram_block3a410))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.cin(gnd),
	.combout(ramiframload_4),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[4]~16 .lut_mask = 16'hFD75;
defparam \ramif.ramload[4]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N12
cycloneive_lcell_comb \ramif.ramload[5]~17 (
// Equation(s):
// ramiframload_5 = (always1 & ((address_reg_a_0 & (ram_block3a371)) # (!address_reg_a_0 & ((ram_block3a510)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_5),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[5]~17 .lut_mask = 16'hD800;
defparam \ramif.ramload[5]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N26
cycloneive_lcell_comb \ramif.ramload[6]~18 (
// Equation(s):
// ramiframload_6 = ((address_reg_a_0 & ((ram_block3a381))) # (!address_reg_a_0 & (ram_block3a64))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.cin(gnd),
	.combout(ramiframload_6),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[6]~18 .lut_mask = 16'hFD75;
defparam \ramif.ramload[6]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N28
cycloneive_lcell_comb \ramif.ramload[7]~19 (
// Equation(s):
// ramiframload_7 = ((address_reg_a_0 & (ram_block3a391)) # (!address_reg_a_0 & ((ram_block3a71)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.cin(gnd),
	.combout(ramiframload_7),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[7]~19 .lut_mask = 16'hF7D5;
defparam \ramif.ramload[7]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N22
cycloneive_lcell_comb \ramif.ramload[8]~20 (
// Equation(s):
// ramiframload_8 = (always1 & ((address_reg_a_0 & (ram_block3a401)) # (!address_reg_a_0 & ((ram_block3a81)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_8),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[8]~20 .lut_mask = 16'hB800;
defparam \ramif.ramload[8]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N28
cycloneive_lcell_comb \ramif.ramload[9]~21 (
// Equation(s):
// ramiframload_9 = ((address_reg_a_0 & ((ram_block3a412))) # (!address_reg_a_0 & (ram_block3a91))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.cin(gnd),
	.combout(ramiframload_9),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[9]~21 .lut_mask = 16'hFB73;
defparam \ramif.ramload[9]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N22
cycloneive_lcell_comb \ramif.ramload[10]~22 (
// Equation(s):
// ramiframload_10 = (always1 & ((address_reg_a_0 & ((ram_block3a421))) # (!address_reg_a_0 & (ram_block3a101))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.cin(gnd),
	.combout(ramiframload_10),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[10]~22 .lut_mask = 16'hC808;
defparam \ramif.ramload[10]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N4
cycloneive_lcell_comb \ramif.ramload[11]~23 (
// Equation(s):
// ramiframload_11 = ((address_reg_a_0 & ((ram_block3a431))) # (!address_reg_a_0 & (ram_block3a112))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_11),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[11]~23 .lut_mask = 16'hE4FF;
defparam \ramif.ramload[11]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N12
cycloneive_lcell_comb \ramif.ramload[12]~24 (
// Equation(s):
// ramiframload_12 = ((address_reg_a_0 & ((ram_block3a441))) # (!address_reg_a_0 & (ram_block3a121))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_12),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[12]~24 .lut_mask = 16'hE2FF;
defparam \ramif.ramload[12]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N26
cycloneive_lcell_comb \ramif.ramload[13]~25 (
// Equation(s):
// ramiframload_13 = ((address_reg_a_0 & ((ram_block3a451))) # (!address_reg_a_0 & (ram_block3a131))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_13),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[13]~25 .lut_mask = 16'hCAFF;
defparam \ramif.ramload[13]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N12
cycloneive_lcell_comb \ramif.ramload[14]~26 (
// Equation(s):
// ramiframload_14 = (always1 & ((address_reg_a_0 & ((ram_block3a461))) # (!address_reg_a_0 & (ram_block3a141))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.cin(gnd),
	.combout(ramiframload_14),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[14]~26 .lut_mask = 16'hC840;
defparam \ramif.ramload[14]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N2
cycloneive_lcell_comb \ramif.ramload[15]~27 (
// Equation(s):
// ramiframload_15 = ((address_reg_a_0 & ((ram_block3a471))) # (!address_reg_a_0 & (ram_block3a151))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.cin(gnd),
	.combout(ramiframload_15),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[15]~27 .lut_mask = 16'hFB3B;
defparam \ramif.ramload[15]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N10
cycloneive_lcell_comb \ramif.ramload[16]~28 (
// Equation(s):
// ramiframload_16 = ((address_reg_a_0 & ((ram_block3a481))) # (!address_reg_a_0 & (ram_block3a161))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_16),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[16]~28 .lut_mask = 16'hE4FF;
defparam \ramif.ramload[16]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N18
cycloneive_lcell_comb \ramif.ramload[17]~29 (
// Equation(s):
// ramiframload_17 = (always1 & ((address_reg_a_0 & (ram_block3a491)) # (!address_reg_a_0 & ((ram_block3a171)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_17),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[17]~29 .lut_mask = 16'hB800;
defparam \ramif.ramload[17]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N0
cycloneive_lcell_comb \ramif.ramload[18]~30 (
// Equation(s):
// ramiframload_18 = (always1 & ((address_reg_a_0 & (ram_block3a501)) # (!address_reg_a_0 & ((ram_block3a181)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_18),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[18]~30 .lut_mask = 16'hAC00;
defparam \ramif.ramload[18]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N24
cycloneive_lcell_comb \ramif.ramload[19]~31 (
// Equation(s):
// ramiframload_19 = (always1 & ((address_reg_a_0 & ((ram_block3a512))) # (!address_reg_a_0 & (ram_block3a191))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_19),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[19]~31 .lut_mask = 16'hE400;
defparam \ramif.ramload[19]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N18
cycloneive_lcell_comb \ramif.ramload[20]~32 (
// Equation(s):
// ramiframload_20 = ((address_reg_a_0 & ((ram_block3a521))) # (!address_reg_a_0 & (ram_block3a201))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_20),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[20]~32 .lut_mask = 16'hE2FF;
defparam \ramif.ramload[20]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N20
cycloneive_lcell_comb \ramif.ramload[21]~33 (
// Equation(s):
// ramiframload_21 = (always1 & ((address_reg_a_0 & (ram_block3a531)) # (!address_reg_a_0 & ((ram_block3a212)))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.cin(gnd),
	.combout(ramiframload_21),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[21]~33 .lut_mask = 16'hA280;
defparam \ramif.ramload[21]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N2
cycloneive_lcell_comb \ramif.ramload[22]~34 (
// Equation(s):
// ramiframload_22 = ((address_reg_a_0 & ((ram_block3a541))) # (!address_reg_a_0 & (ram_block3a221))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_22),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[22]~34 .lut_mask = 16'hE2FF;
defparam \ramif.ramload[22]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N30
cycloneive_lcell_comb \ramif.ramload[23]~35 (
// Equation(s):
// ramiframload_23 = ((address_reg_a_0 & ((ram_block3a551))) # (!address_reg_a_0 & (ram_block3a231))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.cin(gnd),
	.combout(ramiframload_23),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[23]~35 .lut_mask = 16'hFD75;
defparam \ramif.ramload[23]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N0
cycloneive_lcell_comb \ramif.ramload[24]~36 (
// Equation(s):
// ramiframload_24 = (always1 & ((address_reg_a_0 & ((ram_block3a561))) # (!address_reg_a_0 & (ram_block3a241))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.cin(gnd),
	.combout(ramiframload_24),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[24]~36 .lut_mask = 16'hE020;
defparam \ramif.ramload[24]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N28
cycloneive_lcell_comb \ramif.ramload[25]~37 (
// Equation(s):
// ramiframload_25 = ((address_reg_a_0 & (ram_block3a571)) # (!address_reg_a_0 & ((ram_block3a251)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.cin(gnd),
	.combout(ramiframload_25),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[25]~37 .lut_mask = 16'hF7D5;
defparam \ramif.ramload[25]~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N22
cycloneive_lcell_comb \ramif.ramload[26]~38 (
// Equation(s):
// ramiframload_26 = (address_reg_a_0 & ((ram_block3a581))) # (!address_reg_a_0 & (ram_block3a261))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(gnd),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.cin(gnd),
	.combout(ramiframload_26),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[26]~38 .lut_mask = 16'hEE22;
defparam \ramif.ramload[26]~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N24
cycloneive_lcell_comb \ramif.ramload[27]~39 (
// Equation(s):
// ramiframload_27 = (address_reg_a_0 & (ram_block3a591)) # (!address_reg_a_0 & ((ram_block3a271)))

	.dataa(gnd),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.cin(gnd),
	.combout(ramiframload_27),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[27]~39 .lut_mask = 16'hF3C0;
defparam \ramif.ramload[27]~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N6
cycloneive_lcell_comb \ramif.ramload[28]~40 (
// Equation(s):
// ramiframload_28 = (address_reg_a_0 & ((ram_block3a601))) # (!address_reg_a_0 & (ram_block3a281))

	.dataa(gnd),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.cin(gnd),
	.combout(ramiframload_28),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[28]~40 .lut_mask = 16'hFC30;
defparam \ramif.ramload[28]~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N4
cycloneive_lcell_comb \ramif.ramload[29]~41 (
// Equation(s):
// ramiframload_29 = (address_reg_a_0 & (ram_block3a611)) # (!address_reg_a_0 & ((ram_block3a291)))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(gnd),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.cin(gnd),
	.combout(ramiframload_29),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[29]~41 .lut_mask = 16'hF5A0;
defparam \ramif.ramload[29]~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N6
cycloneive_lcell_comb \ramif.ramload[30]~42 (
// Equation(s):
// ramiframload_30 = (address_reg_a_0 & (ram_block3a621)) # (!address_reg_a_0 & ((ram_block3a301)))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(gnd),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.cin(gnd),
	.combout(ramiframload_30),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[30]~42 .lut_mask = 16'hF5A0;
defparam \ramif.ramload[30]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N8
cycloneive_lcell_comb \ramif.ramload[31]~43 (
// Equation(s):
// ramiframload_31 = (address_reg_a_0 & ((ram_block3a631))) # (!address_reg_a_0 & (ram_block3a312))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(gnd),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.cin(gnd),
	.combout(ramiframload_31),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[31]~43 .lut_mask = 16'hFA50;
defparam \ramif.ramload[31]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N30
cycloneive_lcell_comb \ramif.ramload[26]~44 (
// Equation(s):
// ramiframload_261 = (always1 & ((address_reg_a_0 & ((ram_block3a581))) # (!address_reg_a_0 & (ram_block3a261))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.cin(gnd),
	.combout(ramiframload_261),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[26]~44 .lut_mask = 16'hE020;
defparam \ramif.ramload[26]~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N6
cycloneive_lcell_comb \ramif.ramload[27]~45 (
// Equation(s):
// ramiframload_271 = ((address_reg_a_0 & ((ram_block3a591))) # (!address_reg_a_0 & (ram_block3a271))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_271),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[27]~45 .lut_mask = 16'hE4FF;
defparam \ramif.ramload[27]~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N8
cycloneive_lcell_comb \ramif.ramload[28]~46 (
// Equation(s):
// ramiframload_281 = ((address_reg_a_0 & (ram_block3a601)) # (!address_reg_a_0 & ((ram_block3a281)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.cin(gnd),
	.combout(ramiframload_281),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[28]~46 .lut_mask = 16'hBFB3;
defparam \ramif.ramload[28]~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N2
cycloneive_lcell_comb \ramif.ramload[29]~47 (
// Equation(s):
// ramiframload_291 = ((address_reg_a_0 & ((ram_block3a611))) # (!address_reg_a_0 & (ram_block3a291))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.cin(gnd),
	.combout(ramiframload_291),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[29]~47 .lut_mask = 16'hEF2F;
defparam \ramif.ramload[29]~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N16
cycloneive_lcell_comb \ramif.ramload[30]~48 (
// Equation(s):
// ramiframload_301 = (always1 & ((address_reg_a_0 & (ram_block3a621)) # (!address_reg_a_0 & ((ram_block3a301)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.cin(gnd),
	.combout(ramiframload_301),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[30]~48 .lut_mask = 16'hC480;
defparam \ramif.ramload[30]~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N6
cycloneive_lcell_comb \ramif.ramload[31]~49 (
// Equation(s):
// ramiframload_311 = ((address_reg_a_0 & ((ram_block3a631))) # (!address_reg_a_0 & (ram_block3a312))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_311),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[31]~49 .lut_mask = 16'hE4FF;
defparam \ramif.ramload[31]~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N15
dffeas \addr[9] (
	.clk(CLK),
	.d(ramaddr8),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[9]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[9] .is_wysiwyg = "true";
defparam \addr[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N1
dffeas \addr[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr9),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[8]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[8] .is_wysiwyg = "true";
defparam \addr[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N0
cycloneive_lcell_comb \always0~5 (
// Equation(s):
// \always0~5_combout  = (\ramaddr~19_combout  & (addr[8] & (addr[9] $ (!\ramaddr~17_combout )))) # (!\ramaddr~19_combout  & (!addr[8] & (addr[9] $ (!\ramaddr~17_combout ))))

	.dataa(ramaddr9),
	.datab(addr[9]),
	.datac(addr[8]),
	.datad(ramaddr8),
	.cin(gnd),
	.combout(\always0~5_combout ),
	.cout());
// synopsys translate_off
defparam \always0~5 .lut_mask = 16'h8421;
defparam \always0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N19
dffeas \addr[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr12),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[13]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[13] .is_wysiwyg = "true";
defparam \addr[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N9
dffeas \addr[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr13),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[12]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[12] .is_wysiwyg = "true";
defparam \addr[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N8
cycloneive_lcell_comb \always0~7 (
// Equation(s):
// \always0~7_combout  = (\ramaddr~25_combout  & (addr[13] & (addr[12] $ (!\ramaddr~27_combout )))) # (!\ramaddr~25_combout  & (!addr[13] & (addr[12] $ (!\ramaddr~27_combout ))))

	.dataa(ramaddr12),
	.datab(addr[13]),
	.datac(addr[12]),
	.datad(ramaddr13),
	.cin(gnd),
	.combout(\always0~7_combout ),
	.cout());
// synopsys translate_off
defparam \always0~7 .lut_mask = 16'h9009;
defparam \always0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y36_N13
dffeas \addr[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr15),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[14]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[14] .is_wysiwyg = "true";
defparam \addr[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N12
cycloneive_lcell_comb \always0~8 (
// Equation(s):
// \always0~8_combout  = (addr[15] & (!\ramaddr~29_combout  & (\ramaddr~31_combout  $ (!addr[14])))) # (!addr[15] & (\ramaddr~29_combout  & (\ramaddr~31_combout  $ (!addr[14]))))

	.dataa(addr[15]),
	.datab(ramaddr15),
	.datac(addr[14]),
	.datad(ramaddr14),
	.cin(gnd),
	.combout(\always0~8_combout ),
	.cout());
// synopsys translate_off
defparam \always0~8 .lut_mask = 16'h4182;
defparam \always0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N20
cycloneive_lcell_comb \always0~9 (
// Equation(s):
// \always0~9_combout  = (\always0~7_combout  & \always0~8_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\always0~7_combout ),
	.datad(\always0~8_combout ),
	.cin(gnd),
	.combout(\always0~9_combout ),
	.cout());
// synopsys translate_off
defparam \always0~9 .lut_mask = 16'hF000;
defparam \always0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y36_N29
dffeas \addr[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr1),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[0]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[0] .is_wysiwyg = "true";
defparam \addr[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N28
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// \always0~0_combout  = (addr[1] & (\ramaddr~1_combout  & (addr[0] $ (!\ramaddr~3_combout )))) # (!addr[1] & (!\ramaddr~1_combout  & (addr[0] $ (!\ramaddr~3_combout ))))

	.dataa(addr[1]),
	.datab(ramaddr),
	.datac(addr[0]),
	.datad(ramaddr1),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'h9009;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y38_N5
dffeas \addr[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr5),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[4]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[4] .is_wysiwyg = "true";
defparam \addr[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N4
cycloneive_lcell_comb \always0~2 (
// Equation(s):
// \always0~2_combout  = (addr[5] & (\ramaddr~9_combout  & (\ramaddr~11_combout  $ (!addr[4])))) # (!addr[5] & (!\ramaddr~9_combout  & (\ramaddr~11_combout  $ (!addr[4]))))

	.dataa(addr[5]),
	.datab(ramaddr5),
	.datac(addr[4]),
	.datad(ramaddr4),
	.cin(gnd),
	.combout(\always0~2_combout ),
	.cout());
// synopsys translate_off
defparam \always0~2 .lut_mask = 16'h8241;
defparam \always0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y35_N29
dffeas \addr[7] (
	.clk(CLK),
	.d(ramaddr6),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[7]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[7] .is_wysiwyg = "true";
defparam \addr[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N7
dffeas \addr[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr7),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[6]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[6] .is_wysiwyg = "true";
defparam \addr[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N6
cycloneive_lcell_comb \always0~3 (
// Equation(s):
// \always0~3_combout  = (\ramaddr~15_combout  & (addr[6] & (addr[7] $ (!\ramaddr~13_combout )))) # (!\ramaddr~15_combout  & (!addr[6] & (addr[7] $ (!\ramaddr~13_combout ))))

	.dataa(ramaddr7),
	.datab(addr[7]),
	.datac(addr[6]),
	.datad(ramaddr6),
	.cin(gnd),
	.combout(\always0~3_combout ),
	.cout());
// synopsys translate_off
defparam \always0~3 .lut_mask = 16'h8421;
defparam \always0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N26
cycloneive_lcell_comb \always0~4 (
// Equation(s):
// \always0~4_combout  = (\always0~1_combout  & (\always0~0_combout  & (\always0~2_combout  & \always0~3_combout )))

	.dataa(\always0~1_combout ),
	.datab(\always0~0_combout ),
	.datac(\always0~2_combout ),
	.datad(\always0~3_combout ),
	.cin(gnd),
	.combout(\always0~4_combout ),
	.cout());
// synopsys translate_off
defparam \always0~4 .lut_mask = 16'h8000;
defparam \always0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N20
cycloneive_lcell_comb \always0~10 (
// Equation(s):
// \always0~10_combout  = (\always0~6_combout  & (\always0~5_combout  & (\always0~9_combout  & \always0~4_combout )))

	.dataa(\always0~6_combout ),
	.datab(\always0~5_combout ),
	.datac(\always0~9_combout ),
	.datad(\always0~4_combout ),
	.cin(gnd),
	.combout(\always0~10_combout ),
	.cout());
// synopsys translate_off
defparam \always0~10 .lut_mask = 16'h8000;
defparam \always0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N13
dffeas \addr[30] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr27),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[30]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[30] .is_wysiwyg = "true";
defparam \addr[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N12
cycloneive_lcell_comb \always0~19 (
// Equation(s):
// \always0~19_combout  = (addr[31] & (\ramaddr~61_combout  & (\ramaddr~63_combout  $ (!addr[30])))) # (!addr[31] & (!\ramaddr~61_combout  & (\ramaddr~63_combout  $ (!addr[30]))))

	.dataa(addr[31]),
	.datab(ramaddr27),
	.datac(addr[30]),
	.datad(ramaddr26),
	.cin(gnd),
	.combout(\always0~19_combout ),
	.cout());
// synopsys translate_off
defparam \always0~19 .lut_mask = 16'h8241;
defparam \always0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y34_N1
dffeas \addr[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr25),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[28]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[28] .is_wysiwyg = "true";
defparam \addr[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N0
cycloneive_lcell_comb \always0~18 (
// Equation(s):
// \always0~18_combout  = (addr[29] & (\ramaddr~57_combout  & (addr[28] $ (!\ramaddr~59_combout )))) # (!addr[29] & (!\ramaddr~57_combout  & (addr[28] $ (!\ramaddr~59_combout ))))

	.dataa(addr[29]),
	.datab(ramaddr24),
	.datac(addr[28]),
	.datad(ramaddr25),
	.cin(gnd),
	.combout(\always0~18_combout ),
	.cout());
// synopsys translate_off
defparam \always0~18 .lut_mask = 16'h9009;
defparam \always0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N31
dffeas \addr[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr23),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[26]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[26] .is_wysiwyg = "true";
defparam \addr[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N30
cycloneive_lcell_comb \always0~17 (
// Equation(s):
// \always0~17_combout  = (addr[27] & (\ramaddr~53_combout  & (addr[26] $ (!\ramaddr~55_combout )))) # (!addr[27] & (!\ramaddr~53_combout  & (addr[26] $ (!\ramaddr~55_combout ))))

	.dataa(addr[27]),
	.datab(ramaddr22),
	.datac(addr[26]),
	.datad(ramaddr23),
	.cin(gnd),
	.combout(\always0~17_combout ),
	.cout());
// synopsys translate_off
defparam \always0~17 .lut_mask = 16'h9009;
defparam \always0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N4
cycloneive_lcell_comb \always0~20 (
// Equation(s):
// \always0~20_combout  = (\always0~16_combout  & (\always0~19_combout  & (\always0~18_combout  & \always0~17_combout )))

	.dataa(\always0~16_combout ),
	.datab(\always0~19_combout ),
	.datac(\always0~18_combout ),
	.datad(\always0~17_combout ),
	.cin(gnd),
	.combout(\always0~20_combout ),
	.cout());
// synopsys translate_off
defparam \always0~20 .lut_mask = 16'h8000;
defparam \always0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y38_N23
dffeas \addr[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr17),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[18]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[18] .is_wysiwyg = "true";
defparam \addr[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N22
cycloneive_lcell_comb \always0~12 (
// Equation(s):
// \always0~12_combout  = (addr[19] & (\ramaddr~37_combout  & (addr[18] $ (!\ramaddr~39_combout )))) # (!addr[19] & (!\ramaddr~37_combout  & (addr[18] $ (!\ramaddr~39_combout ))))

	.dataa(addr[19]),
	.datab(\ramif.ramaddr [19]),
	.datac(addr[18]),
	.datad(ramaddr17),
	.cin(gnd),
	.combout(\always0~12_combout ),
	.cout());
// synopsys translate_off
defparam \always0~12 .lut_mask = 16'h9009;
defparam \always0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y39_N9
dffeas \addr[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr19),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[23]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[23] .is_wysiwyg = "true";
defparam \addr[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N19
dffeas \addr[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr20),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[22]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[22] .is_wysiwyg = "true";
defparam \addr[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N18
cycloneive_lcell_comb \always0~14 (
// Equation(s):
// \always0~14_combout  = (\ramaddr~45_combout  & (addr[23] & (addr[22] $ (!\ramaddr~47_combout )))) # (!\ramaddr~45_combout  & (!addr[23] & (addr[22] $ (!\ramaddr~47_combout ))))

	.dataa(ramaddr19),
	.datab(addr[23]),
	.datac(addr[22]),
	.datad(ramaddr20),
	.cin(gnd),
	.combout(\always0~14_combout ),
	.cout());
// synopsys translate_off
defparam \always0~14 .lut_mask = 16'h9009;
defparam \always0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y38_N19
dffeas \addr[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr18),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[20]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[20] .is_wysiwyg = "true";
defparam \addr[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N18
cycloneive_lcell_comb \always0~13 (
// Equation(s):
// \always0~13_combout  = (addr[21] & (\ramaddr~41_combout  & (addr[20] $ (!\ramaddr~43_combout )))) # (!addr[21] & (!\ramaddr~41_combout  & (addr[20] $ (!\ramaddr~43_combout ))))

	.dataa(addr[21]),
	.datab(\ramif.ramaddr [21]),
	.datac(addr[20]),
	.datad(ramaddr18),
	.cin(gnd),
	.combout(\always0~13_combout ),
	.cout());
// synopsys translate_off
defparam \always0~13 .lut_mask = 16'h9009;
defparam \always0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N30
cycloneive_lcell_comb \always0~15 (
// Equation(s):
// \always0~15_combout  = (\always0~11_combout  & (\always0~12_combout  & (\always0~14_combout  & \always0~13_combout )))

	.dataa(\always0~11_combout ),
	.datab(\always0~12_combout ),
	.datac(\always0~14_combout ),
	.datad(\always0~13_combout ),
	.cin(gnd),
	.combout(\always0~15_combout ),
	.cout());
// synopsys translate_off
defparam \always0~15 .lut_mask = 16'h8000;
defparam \always0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N14
cycloneive_lcell_comb \always0~21 (
// Equation(s):
// \always0~21_combout  = (\always0~20_combout  & (\always0~15_combout  & ((!\ramWEN~0_combout ) # (!\ramREN~0_combout ))))

	.dataa(ramREN),
	.datab(ramWEN),
	.datac(\always0~20_combout ),
	.datad(\always0~15_combout ),
	.cin(gnd),
	.combout(\always0~21_combout ),
	.cout());
// synopsys translate_off
defparam \always0~21 .lut_mask = 16'h7000;
defparam \always0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N26
cycloneive_lcell_comb \always0~23 (
// Equation(s):
// \always0~23_combout  = (\always0~22_combout ) # ((!\always0~21_combout ) # (!\always0~10_combout ))

	.dataa(\always0~22_combout ),
	.datab(\always0~10_combout ),
	.datac(gnd),
	.datad(\always0~21_combout ),
	.cin(gnd),
	.combout(\always0~23_combout ),
	.cout());
// synopsys translate_off
defparam \always0~23 .lut_mask = 16'hBBFF;
defparam \always0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N28
cycloneive_lcell_comb \count[0]~3 (
// Equation(s):
// \count[0]~3_combout  = (!\always0~23_combout  & (\LessThan1~0_combout  $ (!count[0])))

	.dataa(\LessThan1~0_combout ),
	.datab(gnd),
	.datac(count[0]),
	.datad(\always0~23_combout ),
	.cin(gnd),
	.combout(\count[0]~3_combout ),
	.cout());
// synopsys translate_off
defparam \count[0]~3 .lut_mask = 16'h00A5;
defparam \count[0]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N29
dffeas \count[0] (
	.clk(CLK),
	.d(\count[0]~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[0]),
	.prn(vcc));
// synopsys translate_off
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N8
cycloneive_lcell_comb \count[1]~2 (
// Equation(s):
// \count[1]~2_combout  = (!\always0~23_combout  & (count[1] $ (((!\LessThan1~0_combout  & count[0])))))

	.dataa(\LessThan1~0_combout ),
	.datab(count[0]),
	.datac(count[1]),
	.datad(\always0~23_combout ),
	.cin(gnd),
	.combout(\count[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \count[1]~2 .lut_mask = 16'h00B4;
defparam \count[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N9
dffeas \count[1] (
	.clk(CLK),
	.d(\count[1]~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[1]),
	.prn(vcc));
// synopsys translate_off
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N6
cycloneive_lcell_comb \Add0~1 (
// Equation(s):
// \Add0~1_combout  = count[2] $ (((count[1] & count[0])))

	.dataa(count[2]),
	.datab(count[1]),
	.datac(gnd),
	.datad(count[0]),
	.cin(gnd),
	.combout(\Add0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~1 .lut_mask = 16'h66AA;
defparam \Add0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N22
cycloneive_lcell_comb \count[2]~1 (
// Equation(s):
// \count[2]~1_combout  = (!\always0~23_combout  & ((\LessThan1~0_combout  & (count[2])) # (!\LessThan1~0_combout  & ((\Add0~1_combout )))))

	.dataa(\LessThan1~0_combout ),
	.datab(\always0~23_combout ),
	.datac(count[2]),
	.datad(\Add0~1_combout ),
	.cin(gnd),
	.combout(\count[2]~1_combout ),
	.cout());
// synopsys translate_off
defparam \count[2]~1 .lut_mask = 16'h3120;
defparam \count[2]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N23
dffeas \count[2] (
	.clk(CLK),
	.d(\count[2]~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[2]),
	.prn(vcc));
// synopsys translate_off
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N30
cycloneive_lcell_comb \Add0~0 (
// Equation(s):
// \Add0~0_combout  = count[3] $ (((count[2] & (count[0] & count[1]))))

	.dataa(count[2]),
	.datab(count[0]),
	.datac(count[1]),
	.datad(count[3]),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~0 .lut_mask = 16'h7F80;
defparam \Add0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N20
cycloneive_lcell_comb \count[3]~0 (
// Equation(s):
// \count[3]~0_combout  = (!\always0~23_combout  & ((\LessThan1~0_combout  & ((count[3]))) # (!\LessThan1~0_combout  & (\Add0~0_combout ))))

	.dataa(\LessThan1~0_combout ),
	.datab(\Add0~0_combout ),
	.datac(count[3]),
	.datad(\always0~23_combout ),
	.cin(gnd),
	.combout(\count[3]~0_combout ),
	.cout());
// synopsys translate_off
defparam \count[3]~0 .lut_mask = 16'h00E4;
defparam \count[3]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y37_N21
dffeas \count[3] (
	.clk(CLK),
	.d(\count[3]~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[3]),
	.prn(vcc));
// synopsys translate_off
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N26
cycloneive_lcell_comb \LessThan1~0 (
// Equation(s):
// \LessThan1~0_combout  = (count[3] & ((count[2]) # (count[1])))

	.dataa(count[2]),
	.datab(count[3]),
	.datac(count[1]),
	.datad(gnd),
	.cin(gnd),
	.combout(\LessThan1~0_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan1~0 .lut_mask = 16'hC8C8;
defparam \LessThan1~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module altsyncram_1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	data_a,
	ramaddr1,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	[31:0] data_a;
input 	ramaddr1;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



altsyncram_99f1 auto_generated(
	.ram_block3a32(ram_block3a32),
	.ram_block3a0(ram_block3a0),
	.ram_block3a33(ram_block3a33),
	.ram_block3a1(ram_block3a1),
	.ram_block3a34(ram_block3a34),
	.ram_block3a2(ram_block3a2),
	.ram_block3a35(ram_block3a35),
	.ram_block3a3(ram_block3a3),
	.ram_block3a36(ram_block3a36),
	.ram_block3a4(ram_block3a4),
	.ram_block3a37(ram_block3a37),
	.ram_block3a5(ram_block3a5),
	.ram_block3a38(ram_block3a38),
	.ram_block3a6(ram_block3a6),
	.ram_block3a39(ram_block3a39),
	.ram_block3a7(ram_block3a7),
	.ram_block3a40(ram_block3a40),
	.ram_block3a8(ram_block3a8),
	.ram_block3a41(ram_block3a41),
	.ram_block3a9(ram_block3a9),
	.ram_block3a42(ram_block3a42),
	.ram_block3a10(ram_block3a10),
	.ram_block3a43(ram_block3a43),
	.ram_block3a11(ram_block3a11),
	.ram_block3a44(ram_block3a44),
	.ram_block3a12(ram_block3a12),
	.ram_block3a45(ram_block3a45),
	.ram_block3a13(ram_block3a13),
	.ram_block3a46(ram_block3a46),
	.ram_block3a14(ram_block3a14),
	.ram_block3a47(ram_block3a47),
	.ram_block3a15(ram_block3a15),
	.ram_block3a48(ram_block3a48),
	.ram_block3a16(ram_block3a16),
	.ram_block3a49(ram_block3a49),
	.ram_block3a17(ram_block3a17),
	.ram_block3a50(ram_block3a50),
	.ram_block3a18(ram_block3a18),
	.ram_block3a51(ram_block3a51),
	.ram_block3a19(ram_block3a19),
	.ram_block3a52(ram_block3a52),
	.ram_block3a20(ram_block3a20),
	.ram_block3a53(ram_block3a53),
	.ram_block3a21(ram_block3a21),
	.ram_block3a54(ram_block3a54),
	.ram_block3a22(ram_block3a22),
	.ram_block3a55(ram_block3a55),
	.ram_block3a23(ram_block3a23),
	.ram_block3a56(ram_block3a56),
	.ram_block3a24(ram_block3a24),
	.ram_block3a57(ram_block3a57),
	.ram_block3a25(ram_block3a25),
	.ram_block3a58(ram_block3a58),
	.ram_block3a26(ram_block3a26),
	.ram_block3a59(ram_block3a59),
	.ram_block3a27(ram_block3a27),
	.ram_block3a60(ram_block3a60),
	.ram_block3a28(ram_block3a28),
	.ram_block3a61(ram_block3a61),
	.ram_block3a29(ram_block3a29),
	.ram_block3a62(ram_block3a62),
	.ram_block3a30(ram_block3a30),
	.ram_block3a63(ram_block3a63),
	.ram_block3a31(ram_block3a31),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(address_reg_a_0),
	.address_a({gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.ramaddr1(ramaddr1),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_99f1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	data_a,
	ramaddr1,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	[31:0] data_a;
input 	ramaddr1;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram1|ram_block3a32~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a0~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a33~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a1~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a34~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a2~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a35~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a3~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a36~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a4~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a37~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a5~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a38~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a6~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a39~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a7~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a40~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a8~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a41~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a9~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a42~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a10~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a43~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a11~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a44~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a12~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a45~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a13~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a46~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a14~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a47~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a15~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a48~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a16~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a49~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a17~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a50~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a18~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a51~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a19~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a52~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a20~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a53~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a21~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a54~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a22~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a55~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a23~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a56~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a24~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a57~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a25~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a58~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a26~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a59~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a27~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a60~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a28~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a61~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a29~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a62~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a30~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a63~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a31~PORTBDATAOUT0 ;
wire \mgl_prim2|sdr~0_combout ;
wire [0:0] \altsyncram1|address_reg_b ;
wire [31:0] \mgl_prim2|ram_rom_data_reg ;
wire [13:0] \mgl_prim2|ram_rom_addr_reg ;


sld_mod_ram_rom mgl_prim2(
	.ram_block3a32(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a0(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a33(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a1(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a34(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a2(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a35(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a3(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a36(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a4(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a37(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a5(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a38(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a6(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a39(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a7(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a40(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a8(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a41(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a9(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a42(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a10(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a43(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a11(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a44(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a12(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a45(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a13(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a46(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a14(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a47(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a15(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a48(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a16(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a49(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a17(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a50(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a18(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a51(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a19(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a52(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a20(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a53(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a21(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a54(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a22(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a55(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a23(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a56(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a24(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a57(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a25(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a58(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a26(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a59(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a27(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a60(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a28(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a61(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a29(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a62(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a30(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a63(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a31(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.is_in_use_reg1(is_in_use_reg),
	.ram_rom_data_reg_0(\mgl_prim2|ram_rom_data_reg [0]),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.ram_rom_addr_reg_0(\mgl_prim2|ram_rom_addr_reg [0]),
	.ram_rom_addr_reg_1(\mgl_prim2|ram_rom_addr_reg [1]),
	.ram_rom_addr_reg_2(\mgl_prim2|ram_rom_addr_reg [2]),
	.ram_rom_addr_reg_3(\mgl_prim2|ram_rom_addr_reg [3]),
	.ram_rom_addr_reg_4(\mgl_prim2|ram_rom_addr_reg [4]),
	.ram_rom_addr_reg_5(\mgl_prim2|ram_rom_addr_reg [5]),
	.ram_rom_addr_reg_6(\mgl_prim2|ram_rom_addr_reg [6]),
	.ram_rom_addr_reg_7(\mgl_prim2|ram_rom_addr_reg [7]),
	.ram_rom_addr_reg_8(\mgl_prim2|ram_rom_addr_reg [8]),
	.ram_rom_addr_reg_9(\mgl_prim2|ram_rom_addr_reg [9]),
	.ram_rom_addr_reg_10(\mgl_prim2|ram_rom_addr_reg [10]),
	.ram_rom_addr_reg_11(\mgl_prim2|ram_rom_addr_reg [11]),
	.ram_rom_addr_reg_12(\mgl_prim2|ram_rom_addr_reg [12]),
	.ram_rom_data_reg_1(\mgl_prim2|ram_rom_data_reg [1]),
	.ram_rom_data_reg_2(\mgl_prim2|ram_rom_data_reg [2]),
	.ram_rom_data_reg_3(\mgl_prim2|ram_rom_data_reg [3]),
	.ram_rom_data_reg_4(\mgl_prim2|ram_rom_data_reg [4]),
	.ram_rom_data_reg_5(\mgl_prim2|ram_rom_data_reg [5]),
	.ram_rom_data_reg_6(\mgl_prim2|ram_rom_data_reg [6]),
	.ram_rom_data_reg_7(\mgl_prim2|ram_rom_data_reg [7]),
	.ram_rom_data_reg_8(\mgl_prim2|ram_rom_data_reg [8]),
	.ram_rom_data_reg_9(\mgl_prim2|ram_rom_data_reg [9]),
	.ram_rom_data_reg_10(\mgl_prim2|ram_rom_data_reg [10]),
	.ram_rom_data_reg_11(\mgl_prim2|ram_rom_data_reg [11]),
	.ram_rom_data_reg_12(\mgl_prim2|ram_rom_data_reg [12]),
	.ram_rom_data_reg_13(\mgl_prim2|ram_rom_data_reg [13]),
	.ram_rom_data_reg_14(\mgl_prim2|ram_rom_data_reg [14]),
	.ram_rom_data_reg_15(\mgl_prim2|ram_rom_data_reg [15]),
	.ram_rom_data_reg_16(\mgl_prim2|ram_rom_data_reg [16]),
	.ram_rom_data_reg_17(\mgl_prim2|ram_rom_data_reg [17]),
	.ram_rom_data_reg_18(\mgl_prim2|ram_rom_data_reg [18]),
	.ram_rom_data_reg_19(\mgl_prim2|ram_rom_data_reg [19]),
	.ram_rom_data_reg_20(\mgl_prim2|ram_rom_data_reg [20]),
	.ram_rom_data_reg_21(\mgl_prim2|ram_rom_data_reg [21]),
	.ram_rom_data_reg_22(\mgl_prim2|ram_rom_data_reg [22]),
	.ram_rom_data_reg_23(\mgl_prim2|ram_rom_data_reg [23]),
	.ram_rom_data_reg_24(\mgl_prim2|ram_rom_data_reg [24]),
	.ram_rom_data_reg_25(\mgl_prim2|ram_rom_data_reg [25]),
	.ram_rom_data_reg_26(\mgl_prim2|ram_rom_data_reg [26]),
	.ram_rom_data_reg_27(\mgl_prim2|ram_rom_data_reg [27]),
	.ram_rom_data_reg_28(\mgl_prim2|ram_rom_data_reg [28]),
	.ram_rom_data_reg_29(\mgl_prim2|ram_rom_data_reg [29]),
	.ram_rom_data_reg_30(\mgl_prim2|ram_rom_data_reg [30]),
	.ram_rom_data_reg_31(\mgl_prim2|ram_rom_data_reg [31]),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.ir_in({gnd,irf_reg_3_1,gnd,gnd,irf_reg_0_1}),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.raw_tck(altera_internal_jtag1),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

altsyncram_fta2 altsyncram1(
	.ram_block3a321(ram_block3a32),
	.ram_block3a322(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a01(ram_block3a0),
	.ram_block3a02(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a331(ram_block3a33),
	.ram_block3a332(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a110(ram_block3a1),
	.ram_block3a111(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a341(ram_block3a34),
	.ram_block3a342(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a210(ram_block3a2),
	.ram_block3a211(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a351(ram_block3a35),
	.ram_block3a352(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a310(ram_block3a3),
	.ram_block3a311(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a361(ram_block3a36),
	.ram_block3a362(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a410(ram_block3a4),
	.ram_block3a411(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a371(ram_block3a37),
	.ram_block3a372(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a510(ram_block3a5),
	.ram_block3a511(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a381(ram_block3a38),
	.ram_block3a382(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a64(ram_block3a6),
	.ram_block3a65(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a391(ram_block3a39),
	.ram_block3a392(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a71(ram_block3a7),
	.ram_block3a72(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a401(ram_block3a40),
	.ram_block3a402(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a81(ram_block3a8),
	.ram_block3a82(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a412(ram_block3a41),
	.ram_block3a413(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a91(ram_block3a9),
	.ram_block3a92(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a421(ram_block3a42),
	.ram_block3a422(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a101(ram_block3a10),
	.ram_block3a102(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a431(ram_block3a43),
	.ram_block3a432(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a112(ram_block3a11),
	.ram_block3a113(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a441(ram_block3a44),
	.ram_block3a442(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a121(ram_block3a12),
	.ram_block3a122(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a451(ram_block3a45),
	.ram_block3a452(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a131(ram_block3a13),
	.ram_block3a132(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a461(ram_block3a46),
	.ram_block3a462(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a141(ram_block3a14),
	.ram_block3a142(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a471(ram_block3a47),
	.ram_block3a472(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a151(ram_block3a15),
	.ram_block3a152(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a481(ram_block3a48),
	.ram_block3a482(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a161(ram_block3a16),
	.ram_block3a162(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a491(ram_block3a49),
	.ram_block3a492(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a171(ram_block3a17),
	.ram_block3a172(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a501(ram_block3a50),
	.ram_block3a502(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a181(ram_block3a18),
	.ram_block3a182(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a512(ram_block3a51),
	.ram_block3a513(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a191(ram_block3a19),
	.ram_block3a192(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a521(ram_block3a52),
	.ram_block3a522(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a201(ram_block3a20),
	.ram_block3a202(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a531(ram_block3a53),
	.ram_block3a532(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a212(ram_block3a21),
	.ram_block3a213(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a541(ram_block3a54),
	.ram_block3a542(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a221(ram_block3a22),
	.ram_block3a222(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a551(ram_block3a55),
	.ram_block3a552(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a231(ram_block3a23),
	.ram_block3a232(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a561(ram_block3a56),
	.ram_block3a562(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a241(ram_block3a24),
	.ram_block3a242(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a571(ram_block3a57),
	.ram_block3a572(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a251(ram_block3a25),
	.ram_block3a252(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a581(ram_block3a58),
	.ram_block3a582(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a261(ram_block3a26),
	.ram_block3a262(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a591(ram_block3a59),
	.ram_block3a592(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a271(ram_block3a27),
	.ram_block3a272(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a601(ram_block3a60),
	.ram_block3a602(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a281(ram_block3a28),
	.ram_block3a282(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a611(ram_block3a61),
	.ram_block3a612(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a291(ram_block3a29),
	.ram_block3a292(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a621(ram_block3a62),
	.ram_block3a622(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a301(ram_block3a30),
	.ram_block3a302(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a631(ram_block3a63),
	.ram_block3a632(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a312(ram_block3a31),
	.ram_block3a313(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.data_b({\mgl_prim2|ram_rom_data_reg [31],\mgl_prim2|ram_rom_data_reg [30],\mgl_prim2|ram_rom_data_reg [29],\mgl_prim2|ram_rom_data_reg [28],\mgl_prim2|ram_rom_data_reg [27],\mgl_prim2|ram_rom_data_reg [26],\mgl_prim2|ram_rom_data_reg [25],\mgl_prim2|ram_rom_data_reg [24],\mgl_prim2|ram_rom_data_reg [23],
\mgl_prim2|ram_rom_data_reg [22],\mgl_prim2|ram_rom_data_reg [21],\mgl_prim2|ram_rom_data_reg [20],\mgl_prim2|ram_rom_data_reg [19],\mgl_prim2|ram_rom_data_reg [18],\mgl_prim2|ram_rom_data_reg [17],\mgl_prim2|ram_rom_data_reg [16],\mgl_prim2|ram_rom_data_reg [15],\mgl_prim2|ram_rom_data_reg [14],
\mgl_prim2|ram_rom_data_reg [13],\mgl_prim2|ram_rom_data_reg [12],\mgl_prim2|ram_rom_data_reg [11],\mgl_prim2|ram_rom_data_reg [10],\mgl_prim2|ram_rom_data_reg [9],\mgl_prim2|ram_rom_data_reg [8],\mgl_prim2|ram_rom_data_reg [7],\mgl_prim2|ram_rom_data_reg [6],\mgl_prim2|ram_rom_data_reg [5],
\mgl_prim2|ram_rom_data_reg [4],\mgl_prim2|ram_rom_data_reg [3],\mgl_prim2|ram_rom_data_reg [2],\mgl_prim2|ram_rom_data_reg [1],\mgl_prim2|ram_rom_data_reg [0]}),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.address_b({gnd,\mgl_prim2|ram_rom_addr_reg [12],\mgl_prim2|ram_rom_addr_reg [11],\mgl_prim2|ram_rom_addr_reg [10],\mgl_prim2|ram_rom_addr_reg [9],\mgl_prim2|ram_rom_addr_reg [8],\mgl_prim2|ram_rom_addr_reg [7],\mgl_prim2|ram_rom_addr_reg [6],\mgl_prim2|ram_rom_addr_reg [5],\mgl_prim2|ram_rom_addr_reg [4],
\mgl_prim2|ram_rom_addr_reg [3],\mgl_prim2|ram_rom_addr_reg [2],\mgl_prim2|ram_rom_addr_reg [1],\mgl_prim2|ram_rom_addr_reg [0]}),
	.address_reg_a_0(address_reg_a_0),
	.address_a({gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.ramaddr1(ramaddr1),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.clock1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_fta2 (
	ram_block3a321,
	ram_block3a322,
	ram_block3a01,
	ram_block3a02,
	ram_block3a331,
	ram_block3a332,
	ram_block3a110,
	ram_block3a111,
	ram_block3a341,
	ram_block3a342,
	ram_block3a210,
	ram_block3a211,
	ram_block3a351,
	ram_block3a352,
	ram_block3a310,
	ram_block3a311,
	ram_block3a361,
	ram_block3a362,
	ram_block3a410,
	ram_block3a411,
	ram_block3a371,
	ram_block3a372,
	ram_block3a510,
	ram_block3a511,
	ram_block3a381,
	ram_block3a382,
	ram_block3a64,
	ram_block3a65,
	ram_block3a391,
	ram_block3a392,
	ram_block3a71,
	ram_block3a72,
	ram_block3a401,
	ram_block3a402,
	ram_block3a81,
	ram_block3a82,
	ram_block3a412,
	ram_block3a413,
	ram_block3a91,
	ram_block3a92,
	ram_block3a421,
	ram_block3a422,
	ram_block3a101,
	ram_block3a102,
	ram_block3a431,
	ram_block3a432,
	ram_block3a112,
	ram_block3a113,
	ram_block3a441,
	ram_block3a442,
	ram_block3a121,
	ram_block3a122,
	ram_block3a451,
	ram_block3a452,
	ram_block3a131,
	ram_block3a132,
	ram_block3a461,
	ram_block3a462,
	ram_block3a141,
	ram_block3a142,
	ram_block3a471,
	ram_block3a472,
	ram_block3a151,
	ram_block3a152,
	ram_block3a481,
	ram_block3a482,
	ram_block3a161,
	ram_block3a162,
	ram_block3a491,
	ram_block3a492,
	ram_block3a171,
	ram_block3a172,
	ram_block3a501,
	ram_block3a502,
	ram_block3a181,
	ram_block3a182,
	ram_block3a512,
	ram_block3a513,
	ram_block3a191,
	ram_block3a192,
	ram_block3a521,
	ram_block3a522,
	ram_block3a201,
	ram_block3a202,
	ram_block3a531,
	ram_block3a532,
	ram_block3a212,
	ram_block3a213,
	ram_block3a541,
	ram_block3a542,
	ram_block3a221,
	ram_block3a222,
	ram_block3a551,
	ram_block3a552,
	ram_block3a231,
	ram_block3a232,
	ram_block3a561,
	ram_block3a562,
	ram_block3a241,
	ram_block3a242,
	ram_block3a571,
	ram_block3a572,
	ram_block3a251,
	ram_block3a252,
	ram_block3a581,
	ram_block3a582,
	ram_block3a261,
	ram_block3a262,
	ram_block3a591,
	ram_block3a592,
	ram_block3a271,
	ram_block3a272,
	ram_block3a601,
	ram_block3a602,
	ram_block3a281,
	ram_block3a282,
	ram_block3a611,
	ram_block3a612,
	ram_block3a291,
	ram_block3a292,
	ram_block3a621,
	ram_block3a622,
	ram_block3a301,
	ram_block3a302,
	ram_block3a631,
	ram_block3a632,
	ram_block3a312,
	ram_block3a313,
	data_b,
	ram_rom_addr_reg_13,
	address_b,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	sdr,
	data_a,
	address_reg_b_0,
	ramaddr1,
	irf_reg_2_1,
	state_5,
	clock1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a321;
output 	ram_block3a322;
output 	ram_block3a01;
output 	ram_block3a02;
output 	ram_block3a331;
output 	ram_block3a332;
output 	ram_block3a110;
output 	ram_block3a111;
output 	ram_block3a341;
output 	ram_block3a342;
output 	ram_block3a210;
output 	ram_block3a211;
output 	ram_block3a351;
output 	ram_block3a352;
output 	ram_block3a310;
output 	ram_block3a311;
output 	ram_block3a361;
output 	ram_block3a362;
output 	ram_block3a410;
output 	ram_block3a411;
output 	ram_block3a371;
output 	ram_block3a372;
output 	ram_block3a510;
output 	ram_block3a511;
output 	ram_block3a381;
output 	ram_block3a382;
output 	ram_block3a64;
output 	ram_block3a65;
output 	ram_block3a391;
output 	ram_block3a392;
output 	ram_block3a71;
output 	ram_block3a72;
output 	ram_block3a401;
output 	ram_block3a402;
output 	ram_block3a81;
output 	ram_block3a82;
output 	ram_block3a412;
output 	ram_block3a413;
output 	ram_block3a91;
output 	ram_block3a92;
output 	ram_block3a421;
output 	ram_block3a422;
output 	ram_block3a101;
output 	ram_block3a102;
output 	ram_block3a431;
output 	ram_block3a432;
output 	ram_block3a112;
output 	ram_block3a113;
output 	ram_block3a441;
output 	ram_block3a442;
output 	ram_block3a121;
output 	ram_block3a122;
output 	ram_block3a451;
output 	ram_block3a452;
output 	ram_block3a131;
output 	ram_block3a132;
output 	ram_block3a461;
output 	ram_block3a462;
output 	ram_block3a141;
output 	ram_block3a142;
output 	ram_block3a471;
output 	ram_block3a472;
output 	ram_block3a151;
output 	ram_block3a152;
output 	ram_block3a481;
output 	ram_block3a482;
output 	ram_block3a161;
output 	ram_block3a162;
output 	ram_block3a491;
output 	ram_block3a492;
output 	ram_block3a171;
output 	ram_block3a172;
output 	ram_block3a501;
output 	ram_block3a502;
output 	ram_block3a181;
output 	ram_block3a182;
output 	ram_block3a512;
output 	ram_block3a513;
output 	ram_block3a191;
output 	ram_block3a192;
output 	ram_block3a521;
output 	ram_block3a522;
output 	ram_block3a201;
output 	ram_block3a202;
output 	ram_block3a531;
output 	ram_block3a532;
output 	ram_block3a212;
output 	ram_block3a213;
output 	ram_block3a541;
output 	ram_block3a542;
output 	ram_block3a221;
output 	ram_block3a222;
output 	ram_block3a551;
output 	ram_block3a552;
output 	ram_block3a231;
output 	ram_block3a232;
output 	ram_block3a561;
output 	ram_block3a562;
output 	ram_block3a241;
output 	ram_block3a242;
output 	ram_block3a571;
output 	ram_block3a572;
output 	ram_block3a251;
output 	ram_block3a252;
output 	ram_block3a581;
output 	ram_block3a582;
output 	ram_block3a261;
output 	ram_block3a262;
output 	ram_block3a591;
output 	ram_block3a592;
output 	ram_block3a271;
output 	ram_block3a272;
output 	ram_block3a601;
output 	ram_block3a602;
output 	ram_block3a281;
output 	ram_block3a282;
output 	ram_block3a611;
output 	ram_block3a612;
output 	ram_block3a291;
output 	ram_block3a292;
output 	ram_block3a621;
output 	ram_block3a622;
output 	ram_block3a301;
output 	ram_block3a302;
output 	ram_block3a631;
output 	ram_block3a632;
output 	ram_block3a312;
output 	ram_block3a313;
input 	[31:0] data_b;
input 	ram_rom_addr_reg_13;
input 	[13:0] address_b;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
input 	sdr;
input 	[31:0] data_a;
output 	address_reg_b_0;
input 	ramaddr1;
input 	irf_reg_2_1;
input 	state_5;
input 	clock1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \decode4|eq_node[1]~0_combout ;
wire \decode5|eq_node[1]~0_combout ;
wire \decode4|eq_node[0]~1_combout ;
wire \decode5|eq_node[0]~1_combout ;
wire \address_reg_b[0]~feeder_combout ;

wire [0:0] ram_block3a32_PORTADATAOUT_bus;
wire [0:0] ram_block3a32_PORTBDATAOUT_bus;
wire [0:0] ram_block3a0_PORTADATAOUT_bus;
wire [0:0] ram_block3a0_PORTBDATAOUT_bus;
wire [0:0] ram_block3a33_PORTADATAOUT_bus;
wire [0:0] ram_block3a33_PORTBDATAOUT_bus;
wire [0:0] ram_block3a1_PORTADATAOUT_bus;
wire [0:0] ram_block3a1_PORTBDATAOUT_bus;
wire [0:0] ram_block3a34_PORTADATAOUT_bus;
wire [0:0] ram_block3a34_PORTBDATAOUT_bus;
wire [0:0] ram_block3a2_PORTADATAOUT_bus;
wire [0:0] ram_block3a2_PORTBDATAOUT_bus;
wire [0:0] ram_block3a35_PORTADATAOUT_bus;
wire [0:0] ram_block3a35_PORTBDATAOUT_bus;
wire [0:0] ram_block3a3_PORTADATAOUT_bus;
wire [0:0] ram_block3a3_PORTBDATAOUT_bus;
wire [0:0] ram_block3a36_PORTADATAOUT_bus;
wire [0:0] ram_block3a36_PORTBDATAOUT_bus;
wire [0:0] ram_block3a4_PORTADATAOUT_bus;
wire [0:0] ram_block3a4_PORTBDATAOUT_bus;
wire [0:0] ram_block3a37_PORTADATAOUT_bus;
wire [0:0] ram_block3a37_PORTBDATAOUT_bus;
wire [0:0] ram_block3a5_PORTADATAOUT_bus;
wire [0:0] ram_block3a5_PORTBDATAOUT_bus;
wire [0:0] ram_block3a38_PORTADATAOUT_bus;
wire [0:0] ram_block3a38_PORTBDATAOUT_bus;
wire [0:0] ram_block3a6_PORTADATAOUT_bus;
wire [0:0] ram_block3a6_PORTBDATAOUT_bus;
wire [0:0] ram_block3a39_PORTADATAOUT_bus;
wire [0:0] ram_block3a39_PORTBDATAOUT_bus;
wire [0:0] ram_block3a7_PORTADATAOUT_bus;
wire [0:0] ram_block3a7_PORTBDATAOUT_bus;
wire [0:0] ram_block3a40_PORTADATAOUT_bus;
wire [0:0] ram_block3a40_PORTBDATAOUT_bus;
wire [0:0] ram_block3a8_PORTADATAOUT_bus;
wire [0:0] ram_block3a8_PORTBDATAOUT_bus;
wire [0:0] ram_block3a41_PORTADATAOUT_bus;
wire [0:0] ram_block3a41_PORTBDATAOUT_bus;
wire [0:0] ram_block3a9_PORTADATAOUT_bus;
wire [0:0] ram_block3a9_PORTBDATAOUT_bus;
wire [0:0] ram_block3a42_PORTADATAOUT_bus;
wire [0:0] ram_block3a42_PORTBDATAOUT_bus;
wire [0:0] ram_block3a10_PORTADATAOUT_bus;
wire [0:0] ram_block3a10_PORTBDATAOUT_bus;
wire [0:0] ram_block3a43_PORTADATAOUT_bus;
wire [0:0] ram_block3a43_PORTBDATAOUT_bus;
wire [0:0] ram_block3a11_PORTADATAOUT_bus;
wire [0:0] ram_block3a11_PORTBDATAOUT_bus;
wire [0:0] ram_block3a44_PORTADATAOUT_bus;
wire [0:0] ram_block3a44_PORTBDATAOUT_bus;
wire [0:0] ram_block3a12_PORTADATAOUT_bus;
wire [0:0] ram_block3a12_PORTBDATAOUT_bus;
wire [0:0] ram_block3a45_PORTADATAOUT_bus;
wire [0:0] ram_block3a45_PORTBDATAOUT_bus;
wire [0:0] ram_block3a13_PORTADATAOUT_bus;
wire [0:0] ram_block3a13_PORTBDATAOUT_bus;
wire [0:0] ram_block3a46_PORTADATAOUT_bus;
wire [0:0] ram_block3a46_PORTBDATAOUT_bus;
wire [0:0] ram_block3a14_PORTADATAOUT_bus;
wire [0:0] ram_block3a14_PORTBDATAOUT_bus;
wire [0:0] ram_block3a47_PORTADATAOUT_bus;
wire [0:0] ram_block3a47_PORTBDATAOUT_bus;
wire [0:0] ram_block3a15_PORTADATAOUT_bus;
wire [0:0] ram_block3a15_PORTBDATAOUT_bus;
wire [0:0] ram_block3a48_PORTADATAOUT_bus;
wire [0:0] ram_block3a48_PORTBDATAOUT_bus;
wire [0:0] ram_block3a16_PORTADATAOUT_bus;
wire [0:0] ram_block3a16_PORTBDATAOUT_bus;
wire [0:0] ram_block3a49_PORTADATAOUT_bus;
wire [0:0] ram_block3a49_PORTBDATAOUT_bus;
wire [0:0] ram_block3a17_PORTADATAOUT_bus;
wire [0:0] ram_block3a17_PORTBDATAOUT_bus;
wire [0:0] ram_block3a50_PORTADATAOUT_bus;
wire [0:0] ram_block3a50_PORTBDATAOUT_bus;
wire [0:0] ram_block3a18_PORTADATAOUT_bus;
wire [0:0] ram_block3a18_PORTBDATAOUT_bus;
wire [0:0] ram_block3a51_PORTADATAOUT_bus;
wire [0:0] ram_block3a51_PORTBDATAOUT_bus;
wire [0:0] ram_block3a19_PORTADATAOUT_bus;
wire [0:0] ram_block3a19_PORTBDATAOUT_bus;
wire [0:0] ram_block3a52_PORTADATAOUT_bus;
wire [0:0] ram_block3a52_PORTBDATAOUT_bus;
wire [0:0] ram_block3a20_PORTADATAOUT_bus;
wire [0:0] ram_block3a20_PORTBDATAOUT_bus;
wire [0:0] ram_block3a53_PORTADATAOUT_bus;
wire [0:0] ram_block3a53_PORTBDATAOUT_bus;
wire [0:0] ram_block3a21_PORTADATAOUT_bus;
wire [0:0] ram_block3a21_PORTBDATAOUT_bus;
wire [0:0] ram_block3a54_PORTADATAOUT_bus;
wire [0:0] ram_block3a54_PORTBDATAOUT_bus;
wire [0:0] ram_block3a22_PORTADATAOUT_bus;
wire [0:0] ram_block3a22_PORTBDATAOUT_bus;
wire [0:0] ram_block3a55_PORTADATAOUT_bus;
wire [0:0] ram_block3a55_PORTBDATAOUT_bus;
wire [0:0] ram_block3a23_PORTADATAOUT_bus;
wire [0:0] ram_block3a23_PORTBDATAOUT_bus;
wire [0:0] ram_block3a56_PORTADATAOUT_bus;
wire [0:0] ram_block3a56_PORTBDATAOUT_bus;
wire [0:0] ram_block3a24_PORTADATAOUT_bus;
wire [0:0] ram_block3a24_PORTBDATAOUT_bus;
wire [0:0] ram_block3a57_PORTADATAOUT_bus;
wire [0:0] ram_block3a57_PORTBDATAOUT_bus;
wire [0:0] ram_block3a25_PORTADATAOUT_bus;
wire [0:0] ram_block3a25_PORTBDATAOUT_bus;
wire [0:0] ram_block3a58_PORTADATAOUT_bus;
wire [0:0] ram_block3a58_PORTBDATAOUT_bus;
wire [0:0] ram_block3a26_PORTADATAOUT_bus;
wire [0:0] ram_block3a26_PORTBDATAOUT_bus;
wire [0:0] ram_block3a59_PORTADATAOUT_bus;
wire [0:0] ram_block3a59_PORTBDATAOUT_bus;
wire [0:0] ram_block3a27_PORTADATAOUT_bus;
wire [0:0] ram_block3a27_PORTBDATAOUT_bus;
wire [0:0] ram_block3a60_PORTADATAOUT_bus;
wire [0:0] ram_block3a60_PORTBDATAOUT_bus;
wire [0:0] ram_block3a28_PORTADATAOUT_bus;
wire [0:0] ram_block3a28_PORTBDATAOUT_bus;
wire [0:0] ram_block3a61_PORTADATAOUT_bus;
wire [0:0] ram_block3a61_PORTBDATAOUT_bus;
wire [0:0] ram_block3a29_PORTADATAOUT_bus;
wire [0:0] ram_block3a29_PORTBDATAOUT_bus;
wire [0:0] ram_block3a62_PORTADATAOUT_bus;
wire [0:0] ram_block3a62_PORTBDATAOUT_bus;
wire [0:0] ram_block3a30_PORTADATAOUT_bus;
wire [0:0] ram_block3a30_PORTBDATAOUT_bus;
wire [0:0] ram_block3a63_PORTADATAOUT_bus;
wire [0:0] ram_block3a63_PORTBDATAOUT_bus;
wire [0:0] ram_block3a31_PORTADATAOUT_bus;
wire [0:0] ram_block3a31_PORTBDATAOUT_bus;

assign ram_block3a321 = ram_block3a32_PORTADATAOUT_bus[0];

assign ram_block3a322 = ram_block3a32_PORTBDATAOUT_bus[0];

assign ram_block3a01 = ram_block3a0_PORTADATAOUT_bus[0];

assign ram_block3a02 = ram_block3a0_PORTBDATAOUT_bus[0];

assign ram_block3a331 = ram_block3a33_PORTADATAOUT_bus[0];

assign ram_block3a332 = ram_block3a33_PORTBDATAOUT_bus[0];

assign ram_block3a110 = ram_block3a1_PORTADATAOUT_bus[0];

assign ram_block3a111 = ram_block3a1_PORTBDATAOUT_bus[0];

assign ram_block3a341 = ram_block3a34_PORTADATAOUT_bus[0];

assign ram_block3a342 = ram_block3a34_PORTBDATAOUT_bus[0];

assign ram_block3a210 = ram_block3a2_PORTADATAOUT_bus[0];

assign ram_block3a211 = ram_block3a2_PORTBDATAOUT_bus[0];

assign ram_block3a351 = ram_block3a35_PORTADATAOUT_bus[0];

assign ram_block3a352 = ram_block3a35_PORTBDATAOUT_bus[0];

assign ram_block3a310 = ram_block3a3_PORTADATAOUT_bus[0];

assign ram_block3a311 = ram_block3a3_PORTBDATAOUT_bus[0];

assign ram_block3a361 = ram_block3a36_PORTADATAOUT_bus[0];

assign ram_block3a362 = ram_block3a36_PORTBDATAOUT_bus[0];

assign ram_block3a410 = ram_block3a4_PORTADATAOUT_bus[0];

assign ram_block3a411 = ram_block3a4_PORTBDATAOUT_bus[0];

assign ram_block3a371 = ram_block3a37_PORTADATAOUT_bus[0];

assign ram_block3a372 = ram_block3a37_PORTBDATAOUT_bus[0];

assign ram_block3a510 = ram_block3a5_PORTADATAOUT_bus[0];

assign ram_block3a511 = ram_block3a5_PORTBDATAOUT_bus[0];

assign ram_block3a381 = ram_block3a38_PORTADATAOUT_bus[0];

assign ram_block3a382 = ram_block3a38_PORTBDATAOUT_bus[0];

assign ram_block3a64 = ram_block3a6_PORTADATAOUT_bus[0];

assign ram_block3a65 = ram_block3a6_PORTBDATAOUT_bus[0];

assign ram_block3a391 = ram_block3a39_PORTADATAOUT_bus[0];

assign ram_block3a392 = ram_block3a39_PORTBDATAOUT_bus[0];

assign ram_block3a71 = ram_block3a7_PORTADATAOUT_bus[0];

assign ram_block3a72 = ram_block3a7_PORTBDATAOUT_bus[0];

assign ram_block3a401 = ram_block3a40_PORTADATAOUT_bus[0];

assign ram_block3a402 = ram_block3a40_PORTBDATAOUT_bus[0];

assign ram_block3a81 = ram_block3a8_PORTADATAOUT_bus[0];

assign ram_block3a82 = ram_block3a8_PORTBDATAOUT_bus[0];

assign ram_block3a412 = ram_block3a41_PORTADATAOUT_bus[0];

assign ram_block3a413 = ram_block3a41_PORTBDATAOUT_bus[0];

assign ram_block3a91 = ram_block3a9_PORTADATAOUT_bus[0];

assign ram_block3a92 = ram_block3a9_PORTBDATAOUT_bus[0];

assign ram_block3a421 = ram_block3a42_PORTADATAOUT_bus[0];

assign ram_block3a422 = ram_block3a42_PORTBDATAOUT_bus[0];

assign ram_block3a101 = ram_block3a10_PORTADATAOUT_bus[0];

assign ram_block3a102 = ram_block3a10_PORTBDATAOUT_bus[0];

assign ram_block3a431 = ram_block3a43_PORTADATAOUT_bus[0];

assign ram_block3a432 = ram_block3a43_PORTBDATAOUT_bus[0];

assign ram_block3a112 = ram_block3a11_PORTADATAOUT_bus[0];

assign ram_block3a113 = ram_block3a11_PORTBDATAOUT_bus[0];

assign ram_block3a441 = ram_block3a44_PORTADATAOUT_bus[0];

assign ram_block3a442 = ram_block3a44_PORTBDATAOUT_bus[0];

assign ram_block3a121 = ram_block3a12_PORTADATAOUT_bus[0];

assign ram_block3a122 = ram_block3a12_PORTBDATAOUT_bus[0];

assign ram_block3a451 = ram_block3a45_PORTADATAOUT_bus[0];

assign ram_block3a452 = ram_block3a45_PORTBDATAOUT_bus[0];

assign ram_block3a131 = ram_block3a13_PORTADATAOUT_bus[0];

assign ram_block3a132 = ram_block3a13_PORTBDATAOUT_bus[0];

assign ram_block3a461 = ram_block3a46_PORTADATAOUT_bus[0];

assign ram_block3a462 = ram_block3a46_PORTBDATAOUT_bus[0];

assign ram_block3a141 = ram_block3a14_PORTADATAOUT_bus[0];

assign ram_block3a142 = ram_block3a14_PORTBDATAOUT_bus[0];

assign ram_block3a471 = ram_block3a47_PORTADATAOUT_bus[0];

assign ram_block3a472 = ram_block3a47_PORTBDATAOUT_bus[0];

assign ram_block3a151 = ram_block3a15_PORTADATAOUT_bus[0];

assign ram_block3a152 = ram_block3a15_PORTBDATAOUT_bus[0];

assign ram_block3a481 = ram_block3a48_PORTADATAOUT_bus[0];

assign ram_block3a482 = ram_block3a48_PORTBDATAOUT_bus[0];

assign ram_block3a161 = ram_block3a16_PORTADATAOUT_bus[0];

assign ram_block3a162 = ram_block3a16_PORTBDATAOUT_bus[0];

assign ram_block3a491 = ram_block3a49_PORTADATAOUT_bus[0];

assign ram_block3a492 = ram_block3a49_PORTBDATAOUT_bus[0];

assign ram_block3a171 = ram_block3a17_PORTADATAOUT_bus[0];

assign ram_block3a172 = ram_block3a17_PORTBDATAOUT_bus[0];

assign ram_block3a501 = ram_block3a50_PORTADATAOUT_bus[0];

assign ram_block3a502 = ram_block3a50_PORTBDATAOUT_bus[0];

assign ram_block3a181 = ram_block3a18_PORTADATAOUT_bus[0];

assign ram_block3a182 = ram_block3a18_PORTBDATAOUT_bus[0];

assign ram_block3a512 = ram_block3a51_PORTADATAOUT_bus[0];

assign ram_block3a513 = ram_block3a51_PORTBDATAOUT_bus[0];

assign ram_block3a191 = ram_block3a19_PORTADATAOUT_bus[0];

assign ram_block3a192 = ram_block3a19_PORTBDATAOUT_bus[0];

assign ram_block3a521 = ram_block3a52_PORTADATAOUT_bus[0];

assign ram_block3a522 = ram_block3a52_PORTBDATAOUT_bus[0];

assign ram_block3a201 = ram_block3a20_PORTADATAOUT_bus[0];

assign ram_block3a202 = ram_block3a20_PORTBDATAOUT_bus[0];

assign ram_block3a531 = ram_block3a53_PORTADATAOUT_bus[0];

assign ram_block3a532 = ram_block3a53_PORTBDATAOUT_bus[0];

assign ram_block3a212 = ram_block3a21_PORTADATAOUT_bus[0];

assign ram_block3a213 = ram_block3a21_PORTBDATAOUT_bus[0];

assign ram_block3a541 = ram_block3a54_PORTADATAOUT_bus[0];

assign ram_block3a542 = ram_block3a54_PORTBDATAOUT_bus[0];

assign ram_block3a221 = ram_block3a22_PORTADATAOUT_bus[0];

assign ram_block3a222 = ram_block3a22_PORTBDATAOUT_bus[0];

assign ram_block3a551 = ram_block3a55_PORTADATAOUT_bus[0];

assign ram_block3a552 = ram_block3a55_PORTBDATAOUT_bus[0];

assign ram_block3a231 = ram_block3a23_PORTADATAOUT_bus[0];

assign ram_block3a232 = ram_block3a23_PORTBDATAOUT_bus[0];

assign ram_block3a561 = ram_block3a56_PORTADATAOUT_bus[0];

assign ram_block3a562 = ram_block3a56_PORTBDATAOUT_bus[0];

assign ram_block3a241 = ram_block3a24_PORTADATAOUT_bus[0];

assign ram_block3a242 = ram_block3a24_PORTBDATAOUT_bus[0];

assign ram_block3a571 = ram_block3a57_PORTADATAOUT_bus[0];

assign ram_block3a572 = ram_block3a57_PORTBDATAOUT_bus[0];

assign ram_block3a251 = ram_block3a25_PORTADATAOUT_bus[0];

assign ram_block3a252 = ram_block3a25_PORTBDATAOUT_bus[0];

assign ram_block3a581 = ram_block3a58_PORTADATAOUT_bus[0];

assign ram_block3a582 = ram_block3a58_PORTBDATAOUT_bus[0];

assign ram_block3a261 = ram_block3a26_PORTADATAOUT_bus[0];

assign ram_block3a262 = ram_block3a26_PORTBDATAOUT_bus[0];

assign ram_block3a591 = ram_block3a59_PORTADATAOUT_bus[0];

assign ram_block3a592 = ram_block3a59_PORTBDATAOUT_bus[0];

assign ram_block3a271 = ram_block3a27_PORTADATAOUT_bus[0];

assign ram_block3a272 = ram_block3a27_PORTBDATAOUT_bus[0];

assign ram_block3a601 = ram_block3a60_PORTADATAOUT_bus[0];

assign ram_block3a602 = ram_block3a60_PORTBDATAOUT_bus[0];

assign ram_block3a281 = ram_block3a28_PORTADATAOUT_bus[0];

assign ram_block3a282 = ram_block3a28_PORTBDATAOUT_bus[0];

assign ram_block3a611 = ram_block3a61_PORTADATAOUT_bus[0];

assign ram_block3a612 = ram_block3a61_PORTBDATAOUT_bus[0];

assign ram_block3a291 = ram_block3a29_PORTADATAOUT_bus[0];

assign ram_block3a292 = ram_block3a29_PORTBDATAOUT_bus[0];

assign ram_block3a621 = ram_block3a62_PORTADATAOUT_bus[0];

assign ram_block3a622 = ram_block3a62_PORTBDATAOUT_bus[0];

assign ram_block3a301 = ram_block3a30_PORTADATAOUT_bus[0];

assign ram_block3a302 = ram_block3a30_PORTBDATAOUT_bus[0];

assign ram_block3a631 = ram_block3a63_PORTADATAOUT_bus[0];

assign ram_block3a632 = ram_block3a63_PORTBDATAOUT_bus[0];

assign ram_block3a312 = ram_block3a31_PORTADATAOUT_bus[0];

assign ram_block3a313 = ram_block3a31_PORTBDATAOUT_bus[0];

decode_jsa_1 decode5(
	.ram_rom_addr_reg_13(ram_rom_addr_reg_13),
	.sdr(sdr),
	.eq_node_1(\decode5|eq_node[1]~0_combout ),
	.eq_node_0(\decode5|eq_node[0]~1_combout ),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

decode_jsa decode4(
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.eq_node_1(\decode4|eq_node[1]~0_combout ),
	.eq_node_0(\decode4|eq_node[0]~1_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: M9K_X78_Y32_N0
cycloneive_ram_block ram_block3a32(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a32_PORTADATAOUT_bus),
	.portbdataout(ram_block3a32_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a32.clk0_core_clock_enable = "ena0";
defparam ram_block3a32.clk1_core_clock_enable = "ena1";
defparam ram_block3a32.data_interleave_offset_in_bits = 1;
defparam ram_block3a32.data_interleave_width_in_bits = 1;
defparam ram_block3a32.init_file = "meminit.hex";
defparam ram_block3a32.init_file_layout = "port_a";
defparam ram_block3a32.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a32.operation_mode = "bidir_dual_port";
defparam ram_block3a32.port_a_address_clear = "none";
defparam ram_block3a32.port_a_address_width = 13;
defparam ram_block3a32.port_a_byte_enable_clock = "none";
defparam ram_block3a32.port_a_data_out_clear = "none";
defparam ram_block3a32.port_a_data_out_clock = "none";
defparam ram_block3a32.port_a_data_width = 1;
defparam ram_block3a32.port_a_first_address = 0;
defparam ram_block3a32.port_a_first_bit_number = 0;
defparam ram_block3a32.port_a_last_address = 8191;
defparam ram_block3a32.port_a_logical_ram_depth = 16384;
defparam ram_block3a32.port_a_logical_ram_width = 32;
defparam ram_block3a32.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_address_clear = "none";
defparam ram_block3a32.port_b_address_clock = "clock1";
defparam ram_block3a32.port_b_address_width = 13;
defparam ram_block3a32.port_b_data_in_clock = "clock1";
defparam ram_block3a32.port_b_data_out_clear = "none";
defparam ram_block3a32.port_b_data_out_clock = "none";
defparam ram_block3a32.port_b_data_width = 1;
defparam ram_block3a32.port_b_first_address = 0;
defparam ram_block3a32.port_b_first_bit_number = 0;
defparam ram_block3a32.port_b_last_address = 8191;
defparam ram_block3a32.port_b_logical_ram_depth = 16384;
defparam ram_block3a32.port_b_logical_ram_width = 32;
defparam ram_block3a32.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_read_enable_clock = "clock1";
defparam ram_block3a32.port_b_write_enable_clock = "clock1";
defparam ram_block3a32.ram_block_type = "M9K";
defparam ram_block3a32.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y35_N0
cycloneive_ram_block ram_block3a0(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a0_PORTADATAOUT_bus),
	.portbdataout(ram_block3a0_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a0.clk0_core_clock_enable = "ena0";
defparam ram_block3a0.clk1_core_clock_enable = "ena1";
defparam ram_block3a0.data_interleave_offset_in_bits = 1;
defparam ram_block3a0.data_interleave_width_in_bits = 1;
defparam ram_block3a0.init_file = "meminit.hex";
defparam ram_block3a0.init_file_layout = "port_a";
defparam ram_block3a0.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a0.operation_mode = "bidir_dual_port";
defparam ram_block3a0.port_a_address_clear = "none";
defparam ram_block3a0.port_a_address_width = 13;
defparam ram_block3a0.port_a_byte_enable_clock = "none";
defparam ram_block3a0.port_a_data_out_clear = "none";
defparam ram_block3a0.port_a_data_out_clock = "none";
defparam ram_block3a0.port_a_data_width = 1;
defparam ram_block3a0.port_a_first_address = 0;
defparam ram_block3a0.port_a_first_bit_number = 0;
defparam ram_block3a0.port_a_last_address = 8191;
defparam ram_block3a0.port_a_logical_ram_depth = 16384;
defparam ram_block3a0.port_a_logical_ram_width = 32;
defparam ram_block3a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_address_clear = "none";
defparam ram_block3a0.port_b_address_clock = "clock1";
defparam ram_block3a0.port_b_address_width = 13;
defparam ram_block3a0.port_b_data_in_clock = "clock1";
defparam ram_block3a0.port_b_data_out_clear = "none";
defparam ram_block3a0.port_b_data_out_clock = "none";
defparam ram_block3a0.port_b_data_width = 1;
defparam ram_block3a0.port_b_first_address = 0;
defparam ram_block3a0.port_b_first_bit_number = 0;
defparam ram_block3a0.port_b_last_address = 8191;
defparam ram_block3a0.port_b_logical_ram_depth = 16384;
defparam ram_block3a0.port_b_logical_ram_width = 32;
defparam ram_block3a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_read_enable_clock = "clock1";
defparam ram_block3a0.port_b_write_enable_clock = "clock1";
defparam ram_block3a0.ram_block_type = "M9K";
defparam ram_block3a0.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004004AD3;
// synopsys translate_on

// Location: M9K_X51_Y28_N0
cycloneive_ram_block ram_block3a33(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a33_PORTADATAOUT_bus),
	.portbdataout(ram_block3a33_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a33.clk0_core_clock_enable = "ena0";
defparam ram_block3a33.clk1_core_clock_enable = "ena1";
defparam ram_block3a33.data_interleave_offset_in_bits = 1;
defparam ram_block3a33.data_interleave_width_in_bits = 1;
defparam ram_block3a33.init_file = "meminit.hex";
defparam ram_block3a33.init_file_layout = "port_a";
defparam ram_block3a33.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a33.operation_mode = "bidir_dual_port";
defparam ram_block3a33.port_a_address_clear = "none";
defparam ram_block3a33.port_a_address_width = 13;
defparam ram_block3a33.port_a_byte_enable_clock = "none";
defparam ram_block3a33.port_a_data_out_clear = "none";
defparam ram_block3a33.port_a_data_out_clock = "none";
defparam ram_block3a33.port_a_data_width = 1;
defparam ram_block3a33.port_a_first_address = 0;
defparam ram_block3a33.port_a_first_bit_number = 1;
defparam ram_block3a33.port_a_last_address = 8191;
defparam ram_block3a33.port_a_logical_ram_depth = 16384;
defparam ram_block3a33.port_a_logical_ram_width = 32;
defparam ram_block3a33.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_address_clear = "none";
defparam ram_block3a33.port_b_address_clock = "clock1";
defparam ram_block3a33.port_b_address_width = 13;
defparam ram_block3a33.port_b_data_in_clock = "clock1";
defparam ram_block3a33.port_b_data_out_clear = "none";
defparam ram_block3a33.port_b_data_out_clock = "none";
defparam ram_block3a33.port_b_data_width = 1;
defparam ram_block3a33.port_b_first_address = 0;
defparam ram_block3a33.port_b_first_bit_number = 1;
defparam ram_block3a33.port_b_last_address = 8191;
defparam ram_block3a33.port_b_logical_ram_depth = 16384;
defparam ram_block3a33.port_b_logical_ram_width = 32;
defparam ram_block3a33.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_read_enable_clock = "clock1";
defparam ram_block3a33.port_b_write_enable_clock = "clock1";
defparam ram_block3a33.ram_block_type = "M9K";
defparam ram_block3a33.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y28_N0
cycloneive_ram_block ram_block3a1(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a1_PORTADATAOUT_bus),
	.portbdataout(ram_block3a1_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a1.clk0_core_clock_enable = "ena0";
defparam ram_block3a1.clk1_core_clock_enable = "ena1";
defparam ram_block3a1.data_interleave_offset_in_bits = 1;
defparam ram_block3a1.data_interleave_width_in_bits = 1;
defparam ram_block3a1.init_file = "meminit.hex";
defparam ram_block3a1.init_file_layout = "port_a";
defparam ram_block3a1.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a1.operation_mode = "bidir_dual_port";
defparam ram_block3a1.port_a_address_clear = "none";
defparam ram_block3a1.port_a_address_width = 13;
defparam ram_block3a1.port_a_byte_enable_clock = "none";
defparam ram_block3a1.port_a_data_out_clear = "none";
defparam ram_block3a1.port_a_data_out_clock = "none";
defparam ram_block3a1.port_a_data_width = 1;
defparam ram_block3a1.port_a_first_address = 0;
defparam ram_block3a1.port_a_first_bit_number = 1;
defparam ram_block3a1.port_a_last_address = 8191;
defparam ram_block3a1.port_a_logical_ram_depth = 16384;
defparam ram_block3a1.port_a_logical_ram_width = 32;
defparam ram_block3a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_address_clear = "none";
defparam ram_block3a1.port_b_address_clock = "clock1";
defparam ram_block3a1.port_b_address_width = 13;
defparam ram_block3a1.port_b_data_in_clock = "clock1";
defparam ram_block3a1.port_b_data_out_clear = "none";
defparam ram_block3a1.port_b_data_out_clock = "none";
defparam ram_block3a1.port_b_data_width = 1;
defparam ram_block3a1.port_b_first_address = 0;
defparam ram_block3a1.port_b_first_bit_number = 1;
defparam ram_block3a1.port_b_last_address = 8191;
defparam ram_block3a1.port_b_logical_ram_depth = 16384;
defparam ram_block3a1.port_b_logical_ram_width = 32;
defparam ram_block3a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_read_enable_clock = "clock1";
defparam ram_block3a1.port_b_write_enable_clock = "clock1";
defparam ram_block3a1.ram_block_type = "M9K";
defparam ram_block3a1.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004006E40;
// synopsys translate_on

// Location: M9K_X37_Y31_N0
cycloneive_ram_block ram_block3a34(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a34_PORTADATAOUT_bus),
	.portbdataout(ram_block3a34_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a34.clk0_core_clock_enable = "ena0";
defparam ram_block3a34.clk1_core_clock_enable = "ena1";
defparam ram_block3a34.data_interleave_offset_in_bits = 1;
defparam ram_block3a34.data_interleave_width_in_bits = 1;
defparam ram_block3a34.init_file = "meminit.hex";
defparam ram_block3a34.init_file_layout = "port_a";
defparam ram_block3a34.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a34.operation_mode = "bidir_dual_port";
defparam ram_block3a34.port_a_address_clear = "none";
defparam ram_block3a34.port_a_address_width = 13;
defparam ram_block3a34.port_a_byte_enable_clock = "none";
defparam ram_block3a34.port_a_data_out_clear = "none";
defparam ram_block3a34.port_a_data_out_clock = "none";
defparam ram_block3a34.port_a_data_width = 1;
defparam ram_block3a34.port_a_first_address = 0;
defparam ram_block3a34.port_a_first_bit_number = 2;
defparam ram_block3a34.port_a_last_address = 8191;
defparam ram_block3a34.port_a_logical_ram_depth = 16384;
defparam ram_block3a34.port_a_logical_ram_width = 32;
defparam ram_block3a34.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_address_clear = "none";
defparam ram_block3a34.port_b_address_clock = "clock1";
defparam ram_block3a34.port_b_address_width = 13;
defparam ram_block3a34.port_b_data_in_clock = "clock1";
defparam ram_block3a34.port_b_data_out_clear = "none";
defparam ram_block3a34.port_b_data_out_clock = "none";
defparam ram_block3a34.port_b_data_width = 1;
defparam ram_block3a34.port_b_first_address = 0;
defparam ram_block3a34.port_b_first_bit_number = 2;
defparam ram_block3a34.port_b_last_address = 8191;
defparam ram_block3a34.port_b_logical_ram_depth = 16384;
defparam ram_block3a34.port_b_logical_ram_width = 32;
defparam ram_block3a34.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_read_enable_clock = "clock1";
defparam ram_block3a34.port_b_write_enable_clock = "clock1";
defparam ram_block3a34.ram_block_type = "M9K";
defparam ram_block3a34.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y22_N0
cycloneive_ram_block ram_block3a2(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a2_PORTADATAOUT_bus),
	.portbdataout(ram_block3a2_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a2.clk0_core_clock_enable = "ena0";
defparam ram_block3a2.clk1_core_clock_enable = "ena1";
defparam ram_block3a2.data_interleave_offset_in_bits = 1;
defparam ram_block3a2.data_interleave_width_in_bits = 1;
defparam ram_block3a2.init_file = "meminit.hex";
defparam ram_block3a2.init_file_layout = "port_a";
defparam ram_block3a2.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a2.operation_mode = "bidir_dual_port";
defparam ram_block3a2.port_a_address_clear = "none";
defparam ram_block3a2.port_a_address_width = 13;
defparam ram_block3a2.port_a_byte_enable_clock = "none";
defparam ram_block3a2.port_a_data_out_clear = "none";
defparam ram_block3a2.port_a_data_out_clock = "none";
defparam ram_block3a2.port_a_data_width = 1;
defparam ram_block3a2.port_a_first_address = 0;
defparam ram_block3a2.port_a_first_bit_number = 2;
defparam ram_block3a2.port_a_last_address = 8191;
defparam ram_block3a2.port_a_logical_ram_depth = 16384;
defparam ram_block3a2.port_a_logical_ram_width = 32;
defparam ram_block3a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_address_clear = "none";
defparam ram_block3a2.port_b_address_clock = "clock1";
defparam ram_block3a2.port_b_address_width = 13;
defparam ram_block3a2.port_b_data_in_clock = "clock1";
defparam ram_block3a2.port_b_data_out_clear = "none";
defparam ram_block3a2.port_b_data_out_clock = "none";
defparam ram_block3a2.port_b_data_width = 1;
defparam ram_block3a2.port_b_first_address = 0;
defparam ram_block3a2.port_b_first_bit_number = 2;
defparam ram_block3a2.port_b_last_address = 8191;
defparam ram_block3a2.port_b_logical_ram_depth = 16384;
defparam ram_block3a2.port_b_logical_ram_width = 32;
defparam ram_block3a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_read_enable_clock = "clock1";
defparam ram_block3a2.port_b_write_enable_clock = "clock1";
defparam ram_block3a2.ram_block_type = "M9K";
defparam ram_block3a2.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006AA4C70;
// synopsys translate_on

// Location: M9K_X64_Y26_N0
cycloneive_ram_block ram_block3a35(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a35_PORTADATAOUT_bus),
	.portbdataout(ram_block3a35_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a35.clk0_core_clock_enable = "ena0";
defparam ram_block3a35.clk1_core_clock_enable = "ena1";
defparam ram_block3a35.data_interleave_offset_in_bits = 1;
defparam ram_block3a35.data_interleave_width_in_bits = 1;
defparam ram_block3a35.init_file = "meminit.hex";
defparam ram_block3a35.init_file_layout = "port_a";
defparam ram_block3a35.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a35.operation_mode = "bidir_dual_port";
defparam ram_block3a35.port_a_address_clear = "none";
defparam ram_block3a35.port_a_address_width = 13;
defparam ram_block3a35.port_a_byte_enable_clock = "none";
defparam ram_block3a35.port_a_data_out_clear = "none";
defparam ram_block3a35.port_a_data_out_clock = "none";
defparam ram_block3a35.port_a_data_width = 1;
defparam ram_block3a35.port_a_first_address = 0;
defparam ram_block3a35.port_a_first_bit_number = 3;
defparam ram_block3a35.port_a_last_address = 8191;
defparam ram_block3a35.port_a_logical_ram_depth = 16384;
defparam ram_block3a35.port_a_logical_ram_width = 32;
defparam ram_block3a35.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_address_clear = "none";
defparam ram_block3a35.port_b_address_clock = "clock1";
defparam ram_block3a35.port_b_address_width = 13;
defparam ram_block3a35.port_b_data_in_clock = "clock1";
defparam ram_block3a35.port_b_data_out_clear = "none";
defparam ram_block3a35.port_b_data_out_clock = "none";
defparam ram_block3a35.port_b_data_width = 1;
defparam ram_block3a35.port_b_first_address = 0;
defparam ram_block3a35.port_b_first_bit_number = 3;
defparam ram_block3a35.port_b_last_address = 8191;
defparam ram_block3a35.port_b_logical_ram_depth = 16384;
defparam ram_block3a35.port_b_logical_ram_width = 32;
defparam ram_block3a35.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_read_enable_clock = "clock1";
defparam ram_block3a35.port_b_write_enable_clock = "clock1";
defparam ram_block3a35.ram_block_type = "M9K";
defparam ram_block3a35.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y42_N0
cycloneive_ram_block ram_block3a3(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a3_PORTADATAOUT_bus),
	.portbdataout(ram_block3a3_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a3.clk0_core_clock_enable = "ena0";
defparam ram_block3a3.clk1_core_clock_enable = "ena1";
defparam ram_block3a3.data_interleave_offset_in_bits = 1;
defparam ram_block3a3.data_interleave_width_in_bits = 1;
defparam ram_block3a3.init_file = "meminit.hex";
defparam ram_block3a3.init_file_layout = "port_a";
defparam ram_block3a3.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a3.operation_mode = "bidir_dual_port";
defparam ram_block3a3.port_a_address_clear = "none";
defparam ram_block3a3.port_a_address_width = 13;
defparam ram_block3a3.port_a_byte_enable_clock = "none";
defparam ram_block3a3.port_a_data_out_clear = "none";
defparam ram_block3a3.port_a_data_out_clock = "none";
defparam ram_block3a3.port_a_data_width = 1;
defparam ram_block3a3.port_a_first_address = 0;
defparam ram_block3a3.port_a_first_bit_number = 3;
defparam ram_block3a3.port_a_last_address = 8191;
defparam ram_block3a3.port_a_logical_ram_depth = 16384;
defparam ram_block3a3.port_a_logical_ram_width = 32;
defparam ram_block3a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_address_clear = "none";
defparam ram_block3a3.port_b_address_clock = "clock1";
defparam ram_block3a3.port_b_address_width = 13;
defparam ram_block3a3.port_b_data_in_clock = "clock1";
defparam ram_block3a3.port_b_data_out_clear = "none";
defparam ram_block3a3.port_b_data_out_clock = "none";
defparam ram_block3a3.port_b_data_width = 1;
defparam ram_block3a3.port_b_first_address = 0;
defparam ram_block3a3.port_b_first_bit_number = 3;
defparam ram_block3a3.port_b_last_address = 8191;
defparam ram_block3a3.port_b_logical_ram_depth = 16384;
defparam ram_block3a3.port_b_logical_ram_width = 32;
defparam ram_block3a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_read_enable_clock = "clock1";
defparam ram_block3a3.port_b_write_enable_clock = "clock1";
defparam ram_block3a3.ram_block_type = "M9K";
defparam ram_block3a3.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004CC0841;
// synopsys translate_on

// Location: M9K_X78_Y38_N0
cycloneive_ram_block ram_block3a36(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a36_PORTADATAOUT_bus),
	.portbdataout(ram_block3a36_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a36.clk0_core_clock_enable = "ena0";
defparam ram_block3a36.clk1_core_clock_enable = "ena1";
defparam ram_block3a36.data_interleave_offset_in_bits = 1;
defparam ram_block3a36.data_interleave_width_in_bits = 1;
defparam ram_block3a36.init_file = "meminit.hex";
defparam ram_block3a36.init_file_layout = "port_a";
defparam ram_block3a36.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a36.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a36.operation_mode = "bidir_dual_port";
defparam ram_block3a36.port_a_address_clear = "none";
defparam ram_block3a36.port_a_address_width = 13;
defparam ram_block3a36.port_a_byte_enable_clock = "none";
defparam ram_block3a36.port_a_data_out_clear = "none";
defparam ram_block3a36.port_a_data_out_clock = "none";
defparam ram_block3a36.port_a_data_width = 1;
defparam ram_block3a36.port_a_first_address = 0;
defparam ram_block3a36.port_a_first_bit_number = 4;
defparam ram_block3a36.port_a_last_address = 8191;
defparam ram_block3a36.port_a_logical_ram_depth = 16384;
defparam ram_block3a36.port_a_logical_ram_width = 32;
defparam ram_block3a36.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_address_clear = "none";
defparam ram_block3a36.port_b_address_clock = "clock1";
defparam ram_block3a36.port_b_address_width = 13;
defparam ram_block3a36.port_b_data_in_clock = "clock1";
defparam ram_block3a36.port_b_data_out_clear = "none";
defparam ram_block3a36.port_b_data_out_clock = "none";
defparam ram_block3a36.port_b_data_width = 1;
defparam ram_block3a36.port_b_first_address = 0;
defparam ram_block3a36.port_b_first_bit_number = 4;
defparam ram_block3a36.port_b_last_address = 8191;
defparam ram_block3a36.port_b_logical_ram_depth = 16384;
defparam ram_block3a36.port_b_logical_ram_width = 32;
defparam ram_block3a36.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_read_enable_clock = "clock1";
defparam ram_block3a36.port_b_write_enable_clock = "clock1";
defparam ram_block3a36.ram_block_type = "M9K";
defparam ram_block3a36.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y30_N0
cycloneive_ram_block ram_block3a4(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a4_PORTADATAOUT_bus),
	.portbdataout(ram_block3a4_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a4.clk0_core_clock_enable = "ena0";
defparam ram_block3a4.clk1_core_clock_enable = "ena1";
defparam ram_block3a4.data_interleave_offset_in_bits = 1;
defparam ram_block3a4.data_interleave_width_in_bits = 1;
defparam ram_block3a4.init_file = "meminit.hex";
defparam ram_block3a4.init_file_layout = "port_a";
defparam ram_block3a4.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a4.operation_mode = "bidir_dual_port";
defparam ram_block3a4.port_a_address_clear = "none";
defparam ram_block3a4.port_a_address_width = 13;
defparam ram_block3a4.port_a_byte_enable_clock = "none";
defparam ram_block3a4.port_a_data_out_clear = "none";
defparam ram_block3a4.port_a_data_out_clock = "none";
defparam ram_block3a4.port_a_data_width = 1;
defparam ram_block3a4.port_a_first_address = 0;
defparam ram_block3a4.port_a_first_bit_number = 4;
defparam ram_block3a4.port_a_last_address = 8191;
defparam ram_block3a4.port_a_logical_ram_depth = 16384;
defparam ram_block3a4.port_a_logical_ram_width = 32;
defparam ram_block3a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_address_clear = "none";
defparam ram_block3a4.port_b_address_clock = "clock1";
defparam ram_block3a4.port_b_address_width = 13;
defparam ram_block3a4.port_b_data_in_clock = "clock1";
defparam ram_block3a4.port_b_data_out_clear = "none";
defparam ram_block3a4.port_b_data_out_clock = "none";
defparam ram_block3a4.port_b_data_width = 1;
defparam ram_block3a4.port_b_first_address = 0;
defparam ram_block3a4.port_b_first_bit_number = 4;
defparam ram_block3a4.port_b_last_address = 8191;
defparam ram_block3a4.port_b_logical_ram_depth = 16384;
defparam ram_block3a4.port_b_logical_ram_width = 32;
defparam ram_block3a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_read_enable_clock = "clock1";
defparam ram_block3a4.port_b_write_enable_clock = "clock1";
defparam ram_block3a4.ram_block_type = "M9K";
defparam ram_block3a4.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004F0080A;
// synopsys translate_on

// Location: M9K_X64_Y27_N0
cycloneive_ram_block ram_block3a37(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a37_PORTADATAOUT_bus),
	.portbdataout(ram_block3a37_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a37.clk0_core_clock_enable = "ena0";
defparam ram_block3a37.clk1_core_clock_enable = "ena1";
defparam ram_block3a37.data_interleave_offset_in_bits = 1;
defparam ram_block3a37.data_interleave_width_in_bits = 1;
defparam ram_block3a37.init_file = "meminit.hex";
defparam ram_block3a37.init_file_layout = "port_a";
defparam ram_block3a37.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a37.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a37.operation_mode = "bidir_dual_port";
defparam ram_block3a37.port_a_address_clear = "none";
defparam ram_block3a37.port_a_address_width = 13;
defparam ram_block3a37.port_a_byte_enable_clock = "none";
defparam ram_block3a37.port_a_data_out_clear = "none";
defparam ram_block3a37.port_a_data_out_clock = "none";
defparam ram_block3a37.port_a_data_width = 1;
defparam ram_block3a37.port_a_first_address = 0;
defparam ram_block3a37.port_a_first_bit_number = 5;
defparam ram_block3a37.port_a_last_address = 8191;
defparam ram_block3a37.port_a_logical_ram_depth = 16384;
defparam ram_block3a37.port_a_logical_ram_width = 32;
defparam ram_block3a37.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_address_clear = "none";
defparam ram_block3a37.port_b_address_clock = "clock1";
defparam ram_block3a37.port_b_address_width = 13;
defparam ram_block3a37.port_b_data_in_clock = "clock1";
defparam ram_block3a37.port_b_data_out_clear = "none";
defparam ram_block3a37.port_b_data_out_clock = "none";
defparam ram_block3a37.port_b_data_width = 1;
defparam ram_block3a37.port_b_first_address = 0;
defparam ram_block3a37.port_b_first_bit_number = 5;
defparam ram_block3a37.port_b_last_address = 8191;
defparam ram_block3a37.port_b_logical_ram_depth = 16384;
defparam ram_block3a37.port_b_logical_ram_width = 32;
defparam ram_block3a37.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_read_enable_clock = "clock1";
defparam ram_block3a37.port_b_write_enable_clock = "clock1";
defparam ram_block3a37.ram_block_type = "M9K";
defparam ram_block3a37.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y31_N0
cycloneive_ram_block ram_block3a5(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a5_PORTADATAOUT_bus),
	.portbdataout(ram_block3a5_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a5.clk0_core_clock_enable = "ena0";
defparam ram_block3a5.clk1_core_clock_enable = "ena1";
defparam ram_block3a5.data_interleave_offset_in_bits = 1;
defparam ram_block3a5.data_interleave_width_in_bits = 1;
defparam ram_block3a5.init_file = "meminit.hex";
defparam ram_block3a5.init_file_layout = "port_a";
defparam ram_block3a5.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a5.operation_mode = "bidir_dual_port";
defparam ram_block3a5.port_a_address_clear = "none";
defparam ram_block3a5.port_a_address_width = 13;
defparam ram_block3a5.port_a_byte_enable_clock = "none";
defparam ram_block3a5.port_a_data_out_clear = "none";
defparam ram_block3a5.port_a_data_out_clock = "none";
defparam ram_block3a5.port_a_data_width = 1;
defparam ram_block3a5.port_a_first_address = 0;
defparam ram_block3a5.port_a_first_bit_number = 5;
defparam ram_block3a5.port_a_last_address = 8191;
defparam ram_block3a5.port_a_logical_ram_depth = 16384;
defparam ram_block3a5.port_a_logical_ram_width = 32;
defparam ram_block3a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_address_clear = "none";
defparam ram_block3a5.port_b_address_clock = "clock1";
defparam ram_block3a5.port_b_address_width = 13;
defparam ram_block3a5.port_b_data_in_clock = "clock1";
defparam ram_block3a5.port_b_data_out_clear = "none";
defparam ram_block3a5.port_b_data_out_clock = "none";
defparam ram_block3a5.port_b_data_width = 1;
defparam ram_block3a5.port_b_first_address = 0;
defparam ram_block3a5.port_b_first_bit_number = 5;
defparam ram_block3a5.port_b_last_address = 8191;
defparam ram_block3a5.port_b_logical_ram_depth = 16384;
defparam ram_block3a5.port_b_logical_ram_width = 32;
defparam ram_block3a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_read_enable_clock = "clock1";
defparam ram_block3a5.port_b_write_enable_clock = "clock1";
defparam ram_block3a5.ram_block_type = "M9K";
defparam ram_block3a5.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007004EBB;
// synopsys translate_on

// Location: M9K_X37_Y32_N0
cycloneive_ram_block ram_block3a38(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a38_PORTADATAOUT_bus),
	.portbdataout(ram_block3a38_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a38.clk0_core_clock_enable = "ena0";
defparam ram_block3a38.clk1_core_clock_enable = "ena1";
defparam ram_block3a38.data_interleave_offset_in_bits = 1;
defparam ram_block3a38.data_interleave_width_in_bits = 1;
defparam ram_block3a38.init_file = "meminit.hex";
defparam ram_block3a38.init_file_layout = "port_a";
defparam ram_block3a38.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a38.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a38.operation_mode = "bidir_dual_port";
defparam ram_block3a38.port_a_address_clear = "none";
defparam ram_block3a38.port_a_address_width = 13;
defparam ram_block3a38.port_a_byte_enable_clock = "none";
defparam ram_block3a38.port_a_data_out_clear = "none";
defparam ram_block3a38.port_a_data_out_clock = "none";
defparam ram_block3a38.port_a_data_width = 1;
defparam ram_block3a38.port_a_first_address = 0;
defparam ram_block3a38.port_a_first_bit_number = 6;
defparam ram_block3a38.port_a_last_address = 8191;
defparam ram_block3a38.port_a_logical_ram_depth = 16384;
defparam ram_block3a38.port_a_logical_ram_width = 32;
defparam ram_block3a38.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_address_clear = "none";
defparam ram_block3a38.port_b_address_clock = "clock1";
defparam ram_block3a38.port_b_address_width = 13;
defparam ram_block3a38.port_b_data_in_clock = "clock1";
defparam ram_block3a38.port_b_data_out_clear = "none";
defparam ram_block3a38.port_b_data_out_clock = "none";
defparam ram_block3a38.port_b_data_width = 1;
defparam ram_block3a38.port_b_first_address = 0;
defparam ram_block3a38.port_b_first_bit_number = 6;
defparam ram_block3a38.port_b_last_address = 8191;
defparam ram_block3a38.port_b_logical_ram_depth = 16384;
defparam ram_block3a38.port_b_logical_ram_width = 32;
defparam ram_block3a38.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_read_enable_clock = "clock1";
defparam ram_block3a38.port_b_write_enable_clock = "clock1";
defparam ram_block3a38.ram_block_type = "M9K";
defparam ram_block3a38.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y25_N0
cycloneive_ram_block ram_block3a6(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a6_PORTADATAOUT_bus),
	.portbdataout(ram_block3a6_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a6.clk0_core_clock_enable = "ena0";
defparam ram_block3a6.clk1_core_clock_enable = "ena1";
defparam ram_block3a6.data_interleave_offset_in_bits = 1;
defparam ram_block3a6.data_interleave_width_in_bits = 1;
defparam ram_block3a6.init_file = "meminit.hex";
defparam ram_block3a6.init_file_layout = "port_a";
defparam ram_block3a6.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a6.operation_mode = "bidir_dual_port";
defparam ram_block3a6.port_a_address_clear = "none";
defparam ram_block3a6.port_a_address_width = 13;
defparam ram_block3a6.port_a_byte_enable_clock = "none";
defparam ram_block3a6.port_a_data_out_clear = "none";
defparam ram_block3a6.port_a_data_out_clock = "none";
defparam ram_block3a6.port_a_data_width = 1;
defparam ram_block3a6.port_a_first_address = 0;
defparam ram_block3a6.port_a_first_bit_number = 6;
defparam ram_block3a6.port_a_last_address = 8191;
defparam ram_block3a6.port_a_logical_ram_depth = 16384;
defparam ram_block3a6.port_a_logical_ram_width = 32;
defparam ram_block3a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_address_clear = "none";
defparam ram_block3a6.port_b_address_clock = "clock1";
defparam ram_block3a6.port_b_address_width = 13;
defparam ram_block3a6.port_b_data_in_clock = "clock1";
defparam ram_block3a6.port_b_data_out_clear = "none";
defparam ram_block3a6.port_b_data_out_clock = "none";
defparam ram_block3a6.port_b_data_width = 1;
defparam ram_block3a6.port_b_first_address = 0;
defparam ram_block3a6.port_b_first_bit_number = 6;
defparam ram_block3a6.port_b_last_address = 8191;
defparam ram_block3a6.port_b_logical_ram_depth = 16384;
defparam ram_block3a6.port_b_logical_ram_width = 32;
defparam ram_block3a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_read_enable_clock = "clock1";
defparam ram_block3a6.port_b_write_enable_clock = "clock1";
defparam ram_block3a6.ram_block_type = "M9K";
defparam ram_block3a6.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000400210B;
// synopsys translate_on

// Location: M9K_X78_Y39_N0
cycloneive_ram_block ram_block3a39(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a39_PORTADATAOUT_bus),
	.portbdataout(ram_block3a39_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a39.clk0_core_clock_enable = "ena0";
defparam ram_block3a39.clk1_core_clock_enable = "ena1";
defparam ram_block3a39.data_interleave_offset_in_bits = 1;
defparam ram_block3a39.data_interleave_width_in_bits = 1;
defparam ram_block3a39.init_file = "meminit.hex";
defparam ram_block3a39.init_file_layout = "port_a";
defparam ram_block3a39.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a39.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a39.operation_mode = "bidir_dual_port";
defparam ram_block3a39.port_a_address_clear = "none";
defparam ram_block3a39.port_a_address_width = 13;
defparam ram_block3a39.port_a_byte_enable_clock = "none";
defparam ram_block3a39.port_a_data_out_clear = "none";
defparam ram_block3a39.port_a_data_out_clock = "none";
defparam ram_block3a39.port_a_data_width = 1;
defparam ram_block3a39.port_a_first_address = 0;
defparam ram_block3a39.port_a_first_bit_number = 7;
defparam ram_block3a39.port_a_last_address = 8191;
defparam ram_block3a39.port_a_logical_ram_depth = 16384;
defparam ram_block3a39.port_a_logical_ram_width = 32;
defparam ram_block3a39.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_address_clear = "none";
defparam ram_block3a39.port_b_address_clock = "clock1";
defparam ram_block3a39.port_b_address_width = 13;
defparam ram_block3a39.port_b_data_in_clock = "clock1";
defparam ram_block3a39.port_b_data_out_clear = "none";
defparam ram_block3a39.port_b_data_out_clock = "none";
defparam ram_block3a39.port_b_data_width = 1;
defparam ram_block3a39.port_b_first_address = 0;
defparam ram_block3a39.port_b_first_bit_number = 7;
defparam ram_block3a39.port_b_last_address = 8191;
defparam ram_block3a39.port_b_logical_ram_depth = 16384;
defparam ram_block3a39.port_b_logical_ram_width = 32;
defparam ram_block3a39.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_read_enable_clock = "clock1";
defparam ram_block3a39.port_b_write_enable_clock = "clock1";
defparam ram_block3a39.ram_block_type = "M9K";
defparam ram_block3a39.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y36_N0
cycloneive_ram_block ram_block3a7(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a7_PORTADATAOUT_bus),
	.portbdataout(ram_block3a7_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a7.clk0_core_clock_enable = "ena0";
defparam ram_block3a7.clk1_core_clock_enable = "ena1";
defparam ram_block3a7.data_interleave_offset_in_bits = 1;
defparam ram_block3a7.data_interleave_width_in_bits = 1;
defparam ram_block3a7.init_file = "meminit.hex";
defparam ram_block3a7.init_file_layout = "port_a";
defparam ram_block3a7.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a7.operation_mode = "bidir_dual_port";
defparam ram_block3a7.port_a_address_clear = "none";
defparam ram_block3a7.port_a_address_width = 13;
defparam ram_block3a7.port_a_byte_enable_clock = "none";
defparam ram_block3a7.port_a_data_out_clear = "none";
defparam ram_block3a7.port_a_data_out_clock = "none";
defparam ram_block3a7.port_a_data_width = 1;
defparam ram_block3a7.port_a_first_address = 0;
defparam ram_block3a7.port_a_first_bit_number = 7;
defparam ram_block3a7.port_a_last_address = 8191;
defparam ram_block3a7.port_a_logical_ram_depth = 16384;
defparam ram_block3a7.port_a_logical_ram_width = 32;
defparam ram_block3a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_address_clear = "none";
defparam ram_block3a7.port_b_address_clock = "clock1";
defparam ram_block3a7.port_b_address_width = 13;
defparam ram_block3a7.port_b_data_in_clock = "clock1";
defparam ram_block3a7.port_b_data_out_clear = "none";
defparam ram_block3a7.port_b_data_out_clock = "none";
defparam ram_block3a7.port_b_data_width = 1;
defparam ram_block3a7.port_b_first_address = 0;
defparam ram_block3a7.port_b_first_bit_number = 7;
defparam ram_block3a7.port_b_last_address = 8191;
defparam ram_block3a7.port_b_logical_ram_depth = 16384;
defparam ram_block3a7.port_b_logical_ram_width = 32;
defparam ram_block3a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_read_enable_clock = "clock1";
defparam ram_block3a7.port_b_write_enable_clock = "clock1";
defparam ram_block3a7.ram_block_type = "M9K";
defparam ram_block3a7.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000400000E;
// synopsys translate_on

// Location: M9K_X64_Y24_N0
cycloneive_ram_block ram_block3a40(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a40_PORTADATAOUT_bus),
	.portbdataout(ram_block3a40_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a40.clk0_core_clock_enable = "ena0";
defparam ram_block3a40.clk1_core_clock_enable = "ena1";
defparam ram_block3a40.data_interleave_offset_in_bits = 1;
defparam ram_block3a40.data_interleave_width_in_bits = 1;
defparam ram_block3a40.init_file = "meminit.hex";
defparam ram_block3a40.init_file_layout = "port_a";
defparam ram_block3a40.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a40.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a40.operation_mode = "bidir_dual_port";
defparam ram_block3a40.port_a_address_clear = "none";
defparam ram_block3a40.port_a_address_width = 13;
defparam ram_block3a40.port_a_byte_enable_clock = "none";
defparam ram_block3a40.port_a_data_out_clear = "none";
defparam ram_block3a40.port_a_data_out_clock = "none";
defparam ram_block3a40.port_a_data_width = 1;
defparam ram_block3a40.port_a_first_address = 0;
defparam ram_block3a40.port_a_first_bit_number = 8;
defparam ram_block3a40.port_a_last_address = 8191;
defparam ram_block3a40.port_a_logical_ram_depth = 16384;
defparam ram_block3a40.port_a_logical_ram_width = 32;
defparam ram_block3a40.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_address_clear = "none";
defparam ram_block3a40.port_b_address_clock = "clock1";
defparam ram_block3a40.port_b_address_width = 13;
defparam ram_block3a40.port_b_data_in_clock = "clock1";
defparam ram_block3a40.port_b_data_out_clear = "none";
defparam ram_block3a40.port_b_data_out_clock = "none";
defparam ram_block3a40.port_b_data_width = 1;
defparam ram_block3a40.port_b_first_address = 0;
defparam ram_block3a40.port_b_first_bit_number = 8;
defparam ram_block3a40.port_b_last_address = 8191;
defparam ram_block3a40.port_b_logical_ram_depth = 16384;
defparam ram_block3a40.port_b_logical_ram_width = 32;
defparam ram_block3a40.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_read_enable_clock = "clock1";
defparam ram_block3a40.port_b_write_enable_clock = "clock1";
defparam ram_block3a40.ram_block_type = "M9K";
defparam ram_block3a40.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y33_N0
cycloneive_ram_block ram_block3a8(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a8_PORTADATAOUT_bus),
	.portbdataout(ram_block3a8_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a8.clk0_core_clock_enable = "ena0";
defparam ram_block3a8.clk1_core_clock_enable = "ena1";
defparam ram_block3a8.data_interleave_offset_in_bits = 1;
defparam ram_block3a8.data_interleave_width_in_bits = 1;
defparam ram_block3a8.init_file = "meminit.hex";
defparam ram_block3a8.init_file_layout = "port_a";
defparam ram_block3a8.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a8.operation_mode = "bidir_dual_port";
defparam ram_block3a8.port_a_address_clear = "none";
defparam ram_block3a8.port_a_address_width = 13;
defparam ram_block3a8.port_a_byte_enable_clock = "none";
defparam ram_block3a8.port_a_data_out_clear = "none";
defparam ram_block3a8.port_a_data_out_clock = "none";
defparam ram_block3a8.port_a_data_width = 1;
defparam ram_block3a8.port_a_first_address = 0;
defparam ram_block3a8.port_a_first_bit_number = 8;
defparam ram_block3a8.port_a_last_address = 8191;
defparam ram_block3a8.port_a_logical_ram_depth = 16384;
defparam ram_block3a8.port_a_logical_ram_width = 32;
defparam ram_block3a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_address_clear = "none";
defparam ram_block3a8.port_b_address_clock = "clock1";
defparam ram_block3a8.port_b_address_width = 13;
defparam ram_block3a8.port_b_data_in_clock = "clock1";
defparam ram_block3a8.port_b_data_out_clear = "none";
defparam ram_block3a8.port_b_data_out_clock = "none";
defparam ram_block3a8.port_b_data_width = 1;
defparam ram_block3a8.port_b_first_address = 0;
defparam ram_block3a8.port_b_first_bit_number = 8;
defparam ram_block3a8.port_b_last_address = 8191;
defparam ram_block3a8.port_b_logical_ram_depth = 16384;
defparam ram_block3a8.port_b_logical_ram_width = 32;
defparam ram_block3a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_read_enable_clock = "clock1";
defparam ram_block3a8.port_b_write_enable_clock = "clock1";
defparam ram_block3a8.ram_block_type = "M9K";
defparam ram_block3a8.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004003902;
// synopsys translate_on

// Location: M9K_X78_Y27_N0
cycloneive_ram_block ram_block3a41(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a41_PORTADATAOUT_bus),
	.portbdataout(ram_block3a41_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a41.clk0_core_clock_enable = "ena0";
defparam ram_block3a41.clk1_core_clock_enable = "ena1";
defparam ram_block3a41.data_interleave_offset_in_bits = 1;
defparam ram_block3a41.data_interleave_width_in_bits = 1;
defparam ram_block3a41.init_file = "meminit.hex";
defparam ram_block3a41.init_file_layout = "port_a";
defparam ram_block3a41.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a41.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a41.operation_mode = "bidir_dual_port";
defparam ram_block3a41.port_a_address_clear = "none";
defparam ram_block3a41.port_a_address_width = 13;
defparam ram_block3a41.port_a_byte_enable_clock = "none";
defparam ram_block3a41.port_a_data_out_clear = "none";
defparam ram_block3a41.port_a_data_out_clock = "none";
defparam ram_block3a41.port_a_data_width = 1;
defparam ram_block3a41.port_a_first_address = 0;
defparam ram_block3a41.port_a_first_bit_number = 9;
defparam ram_block3a41.port_a_last_address = 8191;
defparam ram_block3a41.port_a_logical_ram_depth = 16384;
defparam ram_block3a41.port_a_logical_ram_width = 32;
defparam ram_block3a41.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_address_clear = "none";
defparam ram_block3a41.port_b_address_clock = "clock1";
defparam ram_block3a41.port_b_address_width = 13;
defparam ram_block3a41.port_b_data_in_clock = "clock1";
defparam ram_block3a41.port_b_data_out_clear = "none";
defparam ram_block3a41.port_b_data_out_clock = "none";
defparam ram_block3a41.port_b_data_width = 1;
defparam ram_block3a41.port_b_first_address = 0;
defparam ram_block3a41.port_b_first_bit_number = 9;
defparam ram_block3a41.port_b_last_address = 8191;
defparam ram_block3a41.port_b_logical_ram_depth = 16384;
defparam ram_block3a41.port_b_logical_ram_width = 32;
defparam ram_block3a41.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_read_enable_clock = "clock1";
defparam ram_block3a41.port_b_write_enable_clock = "clock1";
defparam ram_block3a41.ram_block_type = "M9K";
defparam ram_block3a41.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y30_N0
cycloneive_ram_block ram_block3a9(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a9_PORTADATAOUT_bus),
	.portbdataout(ram_block3a9_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a9.clk0_core_clock_enable = "ena0";
defparam ram_block3a9.clk1_core_clock_enable = "ena1";
defparam ram_block3a9.data_interleave_offset_in_bits = 1;
defparam ram_block3a9.data_interleave_width_in_bits = 1;
defparam ram_block3a9.init_file = "meminit.hex";
defparam ram_block3a9.init_file_layout = "port_a";
defparam ram_block3a9.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a9.operation_mode = "bidir_dual_port";
defparam ram_block3a9.port_a_address_clear = "none";
defparam ram_block3a9.port_a_address_width = 13;
defparam ram_block3a9.port_a_byte_enable_clock = "none";
defparam ram_block3a9.port_a_data_out_clear = "none";
defparam ram_block3a9.port_a_data_out_clock = "none";
defparam ram_block3a9.port_a_data_width = 1;
defparam ram_block3a9.port_a_first_address = 0;
defparam ram_block3a9.port_a_first_bit_number = 9;
defparam ram_block3a9.port_a_last_address = 8191;
defparam ram_block3a9.port_a_logical_ram_depth = 16384;
defparam ram_block3a9.port_a_logical_ram_width = 32;
defparam ram_block3a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_address_clear = "none";
defparam ram_block3a9.port_b_address_clock = "clock1";
defparam ram_block3a9.port_b_address_width = 13;
defparam ram_block3a9.port_b_data_in_clock = "clock1";
defparam ram_block3a9.port_b_data_out_clear = "none";
defparam ram_block3a9.port_b_data_out_clock = "none";
defparam ram_block3a9.port_b_data_width = 1;
defparam ram_block3a9.port_b_first_address = 0;
defparam ram_block3a9.port_b_first_bit_number = 9;
defparam ram_block3a9.port_b_last_address = 8191;
defparam ram_block3a9.port_b_logical_ram_depth = 16384;
defparam ram_block3a9.port_b_logical_ram_width = 32;
defparam ram_block3a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_read_enable_clock = "clock1";
defparam ram_block3a9.port_b_write_enable_clock = "clock1";
defparam ram_block3a9.ram_block_type = "M9K";
defparam ram_block3a9.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004000903;
// synopsys translate_on

// Location: M9K_X64_Y43_N0
cycloneive_ram_block ram_block3a42(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a42_PORTADATAOUT_bus),
	.portbdataout(ram_block3a42_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a42.clk0_core_clock_enable = "ena0";
defparam ram_block3a42.clk1_core_clock_enable = "ena1";
defparam ram_block3a42.data_interleave_offset_in_bits = 1;
defparam ram_block3a42.data_interleave_width_in_bits = 1;
defparam ram_block3a42.init_file = "meminit.hex";
defparam ram_block3a42.init_file_layout = "port_a";
defparam ram_block3a42.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a42.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a42.operation_mode = "bidir_dual_port";
defparam ram_block3a42.port_a_address_clear = "none";
defparam ram_block3a42.port_a_address_width = 13;
defparam ram_block3a42.port_a_byte_enable_clock = "none";
defparam ram_block3a42.port_a_data_out_clear = "none";
defparam ram_block3a42.port_a_data_out_clock = "none";
defparam ram_block3a42.port_a_data_width = 1;
defparam ram_block3a42.port_a_first_address = 0;
defparam ram_block3a42.port_a_first_bit_number = 10;
defparam ram_block3a42.port_a_last_address = 8191;
defparam ram_block3a42.port_a_logical_ram_depth = 16384;
defparam ram_block3a42.port_a_logical_ram_width = 32;
defparam ram_block3a42.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_address_clear = "none";
defparam ram_block3a42.port_b_address_clock = "clock1";
defparam ram_block3a42.port_b_address_width = 13;
defparam ram_block3a42.port_b_data_in_clock = "clock1";
defparam ram_block3a42.port_b_data_out_clear = "none";
defparam ram_block3a42.port_b_data_out_clock = "none";
defparam ram_block3a42.port_b_data_width = 1;
defparam ram_block3a42.port_b_first_address = 0;
defparam ram_block3a42.port_b_first_bit_number = 10;
defparam ram_block3a42.port_b_last_address = 8191;
defparam ram_block3a42.port_b_logical_ram_depth = 16384;
defparam ram_block3a42.port_b_logical_ram_width = 32;
defparam ram_block3a42.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_read_enable_clock = "clock1";
defparam ram_block3a42.port_b_write_enable_clock = "clock1";
defparam ram_block3a42.ram_block_type = "M9K";
defparam ram_block3a42.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y43_N0
cycloneive_ram_block ram_block3a10(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a10_PORTADATAOUT_bus),
	.portbdataout(ram_block3a10_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a10.clk0_core_clock_enable = "ena0";
defparam ram_block3a10.clk1_core_clock_enable = "ena1";
defparam ram_block3a10.data_interleave_offset_in_bits = 1;
defparam ram_block3a10.data_interleave_width_in_bits = 1;
defparam ram_block3a10.init_file = "meminit.hex";
defparam ram_block3a10.init_file_layout = "port_a";
defparam ram_block3a10.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a10.operation_mode = "bidir_dual_port";
defparam ram_block3a10.port_a_address_clear = "none";
defparam ram_block3a10.port_a_address_width = 13;
defparam ram_block3a10.port_a_byte_enable_clock = "none";
defparam ram_block3a10.port_a_data_out_clear = "none";
defparam ram_block3a10.port_a_data_out_clock = "none";
defparam ram_block3a10.port_a_data_width = 1;
defparam ram_block3a10.port_a_first_address = 0;
defparam ram_block3a10.port_a_first_bit_number = 10;
defparam ram_block3a10.port_a_last_address = 8191;
defparam ram_block3a10.port_a_logical_ram_depth = 16384;
defparam ram_block3a10.port_a_logical_ram_width = 32;
defparam ram_block3a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_address_clear = "none";
defparam ram_block3a10.port_b_address_clock = "clock1";
defparam ram_block3a10.port_b_address_width = 13;
defparam ram_block3a10.port_b_data_in_clock = "clock1";
defparam ram_block3a10.port_b_data_out_clear = "none";
defparam ram_block3a10.port_b_data_out_clock = "none";
defparam ram_block3a10.port_b_data_width = 1;
defparam ram_block3a10.port_b_first_address = 0;
defparam ram_block3a10.port_b_first_bit_number = 10;
defparam ram_block3a10.port_b_last_address = 8191;
defparam ram_block3a10.port_b_logical_ram_depth = 16384;
defparam ram_block3a10.port_b_logical_ram_width = 32;
defparam ram_block3a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_read_enable_clock = "clock1";
defparam ram_block3a10.port_b_write_enable_clock = "clock1";
defparam ram_block3a10.ram_block_type = "M9K";
defparam ram_block3a10.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004000102;
// synopsys translate_on

// Location: M9K_X51_Y29_N0
cycloneive_ram_block ram_block3a43(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a43_PORTADATAOUT_bus),
	.portbdataout(ram_block3a43_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a43.clk0_core_clock_enable = "ena0";
defparam ram_block3a43.clk1_core_clock_enable = "ena1";
defparam ram_block3a43.data_interleave_offset_in_bits = 1;
defparam ram_block3a43.data_interleave_width_in_bits = 1;
defparam ram_block3a43.init_file = "meminit.hex";
defparam ram_block3a43.init_file_layout = "port_a";
defparam ram_block3a43.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a43.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a43.operation_mode = "bidir_dual_port";
defparam ram_block3a43.port_a_address_clear = "none";
defparam ram_block3a43.port_a_address_width = 13;
defparam ram_block3a43.port_a_byte_enable_clock = "none";
defparam ram_block3a43.port_a_data_out_clear = "none";
defparam ram_block3a43.port_a_data_out_clock = "none";
defparam ram_block3a43.port_a_data_width = 1;
defparam ram_block3a43.port_a_first_address = 0;
defparam ram_block3a43.port_a_first_bit_number = 11;
defparam ram_block3a43.port_a_last_address = 8191;
defparam ram_block3a43.port_a_logical_ram_depth = 16384;
defparam ram_block3a43.port_a_logical_ram_width = 32;
defparam ram_block3a43.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_address_clear = "none";
defparam ram_block3a43.port_b_address_clock = "clock1";
defparam ram_block3a43.port_b_address_width = 13;
defparam ram_block3a43.port_b_data_in_clock = "clock1";
defparam ram_block3a43.port_b_data_out_clear = "none";
defparam ram_block3a43.port_b_data_out_clock = "none";
defparam ram_block3a43.port_b_data_width = 1;
defparam ram_block3a43.port_b_first_address = 0;
defparam ram_block3a43.port_b_first_bit_number = 11;
defparam ram_block3a43.port_b_last_address = 8191;
defparam ram_block3a43.port_b_logical_ram_depth = 16384;
defparam ram_block3a43.port_b_logical_ram_width = 32;
defparam ram_block3a43.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_read_enable_clock = "clock1";
defparam ram_block3a43.port_b_write_enable_clock = "clock1";
defparam ram_block3a43.ram_block_type = "M9K";
defparam ram_block3a43.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y32_N0
cycloneive_ram_block ram_block3a11(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a11_PORTADATAOUT_bus),
	.portbdataout(ram_block3a11_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a11.clk0_core_clock_enable = "ena0";
defparam ram_block3a11.clk1_core_clock_enable = "ena1";
defparam ram_block3a11.data_interleave_offset_in_bits = 1;
defparam ram_block3a11.data_interleave_width_in_bits = 1;
defparam ram_block3a11.init_file = "meminit.hex";
defparam ram_block3a11.init_file_layout = "port_a";
defparam ram_block3a11.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a11.operation_mode = "bidir_dual_port";
defparam ram_block3a11.port_a_address_clear = "none";
defparam ram_block3a11.port_a_address_width = 13;
defparam ram_block3a11.port_a_byte_enable_clock = "none";
defparam ram_block3a11.port_a_data_out_clear = "none";
defparam ram_block3a11.port_a_data_out_clock = "none";
defparam ram_block3a11.port_a_data_width = 1;
defparam ram_block3a11.port_a_first_address = 0;
defparam ram_block3a11.port_a_first_bit_number = 11;
defparam ram_block3a11.port_a_last_address = 8191;
defparam ram_block3a11.port_a_logical_ram_depth = 16384;
defparam ram_block3a11.port_a_logical_ram_width = 32;
defparam ram_block3a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_address_clear = "none";
defparam ram_block3a11.port_b_address_clock = "clock1";
defparam ram_block3a11.port_b_address_width = 13;
defparam ram_block3a11.port_b_data_in_clock = "clock1";
defparam ram_block3a11.port_b_data_out_clear = "none";
defparam ram_block3a11.port_b_data_out_clock = "none";
defparam ram_block3a11.port_b_data_width = 1;
defparam ram_block3a11.port_b_first_address = 0;
defparam ram_block3a11.port_b_first_bit_number = 11;
defparam ram_block3a11.port_b_last_address = 8191;
defparam ram_block3a11.port_b_logical_ram_depth = 16384;
defparam ram_block3a11.port_b_logical_ram_width = 32;
defparam ram_block3a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_read_enable_clock = "clock1";
defparam ram_block3a11.port_b_write_enable_clock = "clock1";
defparam ram_block3a11.ram_block_type = "M9K";
defparam ram_block3a11.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004005410;
// synopsys translate_on

// Location: M9K_X64_Y29_N0
cycloneive_ram_block ram_block3a44(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a44_PORTADATAOUT_bus),
	.portbdataout(ram_block3a44_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a44.clk0_core_clock_enable = "ena0";
defparam ram_block3a44.clk1_core_clock_enable = "ena1";
defparam ram_block3a44.data_interleave_offset_in_bits = 1;
defparam ram_block3a44.data_interleave_width_in_bits = 1;
defparam ram_block3a44.init_file = "meminit.hex";
defparam ram_block3a44.init_file_layout = "port_a";
defparam ram_block3a44.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a44.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a44.operation_mode = "bidir_dual_port";
defparam ram_block3a44.port_a_address_clear = "none";
defparam ram_block3a44.port_a_address_width = 13;
defparam ram_block3a44.port_a_byte_enable_clock = "none";
defparam ram_block3a44.port_a_data_out_clear = "none";
defparam ram_block3a44.port_a_data_out_clock = "none";
defparam ram_block3a44.port_a_data_width = 1;
defparam ram_block3a44.port_a_first_address = 0;
defparam ram_block3a44.port_a_first_bit_number = 12;
defparam ram_block3a44.port_a_last_address = 8191;
defparam ram_block3a44.port_a_logical_ram_depth = 16384;
defparam ram_block3a44.port_a_logical_ram_width = 32;
defparam ram_block3a44.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_address_clear = "none";
defparam ram_block3a44.port_b_address_clock = "clock1";
defparam ram_block3a44.port_b_address_width = 13;
defparam ram_block3a44.port_b_data_in_clock = "clock1";
defparam ram_block3a44.port_b_data_out_clear = "none";
defparam ram_block3a44.port_b_data_out_clock = "none";
defparam ram_block3a44.port_b_data_width = 1;
defparam ram_block3a44.port_b_first_address = 0;
defparam ram_block3a44.port_b_first_bit_number = 12;
defparam ram_block3a44.port_b_last_address = 8191;
defparam ram_block3a44.port_b_logical_ram_depth = 16384;
defparam ram_block3a44.port_b_logical_ram_width = 32;
defparam ram_block3a44.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_read_enable_clock = "clock1";
defparam ram_block3a44.port_b_write_enable_clock = "clock1";
defparam ram_block3a44.ram_block_type = "M9K";
defparam ram_block3a44.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y33_N0
cycloneive_ram_block ram_block3a12(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a12_PORTADATAOUT_bus),
	.portbdataout(ram_block3a12_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a12.clk0_core_clock_enable = "ena0";
defparam ram_block3a12.clk1_core_clock_enable = "ena1";
defparam ram_block3a12.data_interleave_offset_in_bits = 1;
defparam ram_block3a12.data_interleave_width_in_bits = 1;
defparam ram_block3a12.init_file = "meminit.hex";
defparam ram_block3a12.init_file_layout = "port_a";
defparam ram_block3a12.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a12.operation_mode = "bidir_dual_port";
defparam ram_block3a12.port_a_address_clear = "none";
defparam ram_block3a12.port_a_address_width = 13;
defparam ram_block3a12.port_a_byte_enable_clock = "none";
defparam ram_block3a12.port_a_data_out_clear = "none";
defparam ram_block3a12.port_a_data_out_clock = "none";
defparam ram_block3a12.port_a_data_width = 1;
defparam ram_block3a12.port_a_first_address = 0;
defparam ram_block3a12.port_a_first_bit_number = 12;
defparam ram_block3a12.port_a_last_address = 8191;
defparam ram_block3a12.port_a_logical_ram_depth = 16384;
defparam ram_block3a12.port_a_logical_ram_width = 32;
defparam ram_block3a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_address_clear = "none";
defparam ram_block3a12.port_b_address_clock = "clock1";
defparam ram_block3a12.port_b_address_width = 13;
defparam ram_block3a12.port_b_data_in_clock = "clock1";
defparam ram_block3a12.port_b_data_out_clear = "none";
defparam ram_block3a12.port_b_data_out_clock = "none";
defparam ram_block3a12.port_b_data_width = 1;
defparam ram_block3a12.port_b_first_address = 0;
defparam ram_block3a12.port_b_first_bit_number = 12;
defparam ram_block3a12.port_b_last_address = 8191;
defparam ram_block3a12.port_b_logical_ram_depth = 16384;
defparam ram_block3a12.port_b_logical_ram_width = 32;
defparam ram_block3a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_read_enable_clock = "clock1";
defparam ram_block3a12.port_b_write_enable_clock = "clock1";
defparam ram_block3a12.ram_block_type = "M9K";
defparam ram_block3a12.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004001893;
// synopsys translate_on

// Location: M9K_X78_Y29_N0
cycloneive_ram_block ram_block3a45(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a45_PORTADATAOUT_bus),
	.portbdataout(ram_block3a45_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a45.clk0_core_clock_enable = "ena0";
defparam ram_block3a45.clk1_core_clock_enable = "ena1";
defparam ram_block3a45.data_interleave_offset_in_bits = 1;
defparam ram_block3a45.data_interleave_width_in_bits = 1;
defparam ram_block3a45.init_file = "meminit.hex";
defparam ram_block3a45.init_file_layout = "port_a";
defparam ram_block3a45.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a45.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a45.operation_mode = "bidir_dual_port";
defparam ram_block3a45.port_a_address_clear = "none";
defparam ram_block3a45.port_a_address_width = 13;
defparam ram_block3a45.port_a_byte_enable_clock = "none";
defparam ram_block3a45.port_a_data_out_clear = "none";
defparam ram_block3a45.port_a_data_out_clock = "none";
defparam ram_block3a45.port_a_data_width = 1;
defparam ram_block3a45.port_a_first_address = 0;
defparam ram_block3a45.port_a_first_bit_number = 13;
defparam ram_block3a45.port_a_last_address = 8191;
defparam ram_block3a45.port_a_logical_ram_depth = 16384;
defparam ram_block3a45.port_a_logical_ram_width = 32;
defparam ram_block3a45.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_address_clear = "none";
defparam ram_block3a45.port_b_address_clock = "clock1";
defparam ram_block3a45.port_b_address_width = 13;
defparam ram_block3a45.port_b_data_in_clock = "clock1";
defparam ram_block3a45.port_b_data_out_clear = "none";
defparam ram_block3a45.port_b_data_out_clock = "none";
defparam ram_block3a45.port_b_data_width = 1;
defparam ram_block3a45.port_b_first_address = 0;
defparam ram_block3a45.port_b_first_bit_number = 13;
defparam ram_block3a45.port_b_last_address = 8191;
defparam ram_block3a45.port_b_logical_ram_depth = 16384;
defparam ram_block3a45.port_b_logical_ram_width = 32;
defparam ram_block3a45.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_read_enable_clock = "clock1";
defparam ram_block3a45.port_b_write_enable_clock = "clock1";
defparam ram_block3a45.ram_block_type = "M9K";
defparam ram_block3a45.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y28_N0
cycloneive_ram_block ram_block3a13(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a13_PORTADATAOUT_bus),
	.portbdataout(ram_block3a13_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a13.clk0_core_clock_enable = "ena0";
defparam ram_block3a13.clk1_core_clock_enable = "ena1";
defparam ram_block3a13.data_interleave_offset_in_bits = 1;
defparam ram_block3a13.data_interleave_width_in_bits = 1;
defparam ram_block3a13.init_file = "meminit.hex";
defparam ram_block3a13.init_file_layout = "port_a";
defparam ram_block3a13.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a13.operation_mode = "bidir_dual_port";
defparam ram_block3a13.port_a_address_clear = "none";
defparam ram_block3a13.port_a_address_width = 13;
defparam ram_block3a13.port_a_byte_enable_clock = "none";
defparam ram_block3a13.port_a_data_out_clear = "none";
defparam ram_block3a13.port_a_data_out_clock = "none";
defparam ram_block3a13.port_a_data_width = 1;
defparam ram_block3a13.port_a_first_address = 0;
defparam ram_block3a13.port_a_first_bit_number = 13;
defparam ram_block3a13.port_a_last_address = 8191;
defparam ram_block3a13.port_a_logical_ram_depth = 16384;
defparam ram_block3a13.port_a_logical_ram_width = 32;
defparam ram_block3a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_address_clear = "none";
defparam ram_block3a13.port_b_address_clock = "clock1";
defparam ram_block3a13.port_b_address_width = 13;
defparam ram_block3a13.port_b_data_in_clock = "clock1";
defparam ram_block3a13.port_b_data_out_clear = "none";
defparam ram_block3a13.port_b_data_out_clock = "none";
defparam ram_block3a13.port_b_data_width = 1;
defparam ram_block3a13.port_b_first_address = 0;
defparam ram_block3a13.port_b_first_bit_number = 13;
defparam ram_block3a13.port_b_last_address = 8191;
defparam ram_block3a13.port_b_logical_ram_depth = 16384;
defparam ram_block3a13.port_b_logical_ram_width = 32;
defparam ram_block3a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_read_enable_clock = "clock1";
defparam ram_block3a13.port_b_write_enable_clock = "clock1";
defparam ram_block3a13.ram_block_type = "M9K";
defparam ram_block3a13.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000040068A2;
// synopsys translate_on

// Location: M9K_X51_Y23_N0
cycloneive_ram_block ram_block3a46(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a46_PORTADATAOUT_bus),
	.portbdataout(ram_block3a46_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a46.clk0_core_clock_enable = "ena0";
defparam ram_block3a46.clk1_core_clock_enable = "ena1";
defparam ram_block3a46.data_interleave_offset_in_bits = 1;
defparam ram_block3a46.data_interleave_width_in_bits = 1;
defparam ram_block3a46.init_file = "meminit.hex";
defparam ram_block3a46.init_file_layout = "port_a";
defparam ram_block3a46.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a46.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a46.operation_mode = "bidir_dual_port";
defparam ram_block3a46.port_a_address_clear = "none";
defparam ram_block3a46.port_a_address_width = 13;
defparam ram_block3a46.port_a_byte_enable_clock = "none";
defparam ram_block3a46.port_a_data_out_clear = "none";
defparam ram_block3a46.port_a_data_out_clock = "none";
defparam ram_block3a46.port_a_data_width = 1;
defparam ram_block3a46.port_a_first_address = 0;
defparam ram_block3a46.port_a_first_bit_number = 14;
defparam ram_block3a46.port_a_last_address = 8191;
defparam ram_block3a46.port_a_logical_ram_depth = 16384;
defparam ram_block3a46.port_a_logical_ram_width = 32;
defparam ram_block3a46.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_address_clear = "none";
defparam ram_block3a46.port_b_address_clock = "clock1";
defparam ram_block3a46.port_b_address_width = 13;
defparam ram_block3a46.port_b_data_in_clock = "clock1";
defparam ram_block3a46.port_b_data_out_clear = "none";
defparam ram_block3a46.port_b_data_out_clock = "none";
defparam ram_block3a46.port_b_data_width = 1;
defparam ram_block3a46.port_b_first_address = 0;
defparam ram_block3a46.port_b_first_bit_number = 14;
defparam ram_block3a46.port_b_last_address = 8191;
defparam ram_block3a46.port_b_logical_ram_depth = 16384;
defparam ram_block3a46.port_b_logical_ram_width = 32;
defparam ram_block3a46.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_read_enable_clock = "clock1";
defparam ram_block3a46.port_b_write_enable_clock = "clock1";
defparam ram_block3a46.ram_block_type = "M9K";
defparam ram_block3a46.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y37_N0
cycloneive_ram_block ram_block3a14(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a14_PORTADATAOUT_bus),
	.portbdataout(ram_block3a14_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a14.clk0_core_clock_enable = "ena0";
defparam ram_block3a14.clk1_core_clock_enable = "ena1";
defparam ram_block3a14.data_interleave_offset_in_bits = 1;
defparam ram_block3a14.data_interleave_width_in_bits = 1;
defparam ram_block3a14.init_file = "meminit.hex";
defparam ram_block3a14.init_file_layout = "port_a";
defparam ram_block3a14.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a14.operation_mode = "bidir_dual_port";
defparam ram_block3a14.port_a_address_clear = "none";
defparam ram_block3a14.port_a_address_width = 13;
defparam ram_block3a14.port_a_byte_enable_clock = "none";
defparam ram_block3a14.port_a_data_out_clear = "none";
defparam ram_block3a14.port_a_data_out_clock = "none";
defparam ram_block3a14.port_a_data_width = 1;
defparam ram_block3a14.port_a_first_address = 0;
defparam ram_block3a14.port_a_first_bit_number = 14;
defparam ram_block3a14.port_a_last_address = 8191;
defparam ram_block3a14.port_a_logical_ram_depth = 16384;
defparam ram_block3a14.port_a_logical_ram_width = 32;
defparam ram_block3a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_address_clear = "none";
defparam ram_block3a14.port_b_address_clock = "clock1";
defparam ram_block3a14.port_b_address_width = 13;
defparam ram_block3a14.port_b_data_in_clock = "clock1";
defparam ram_block3a14.port_b_data_out_clear = "none";
defparam ram_block3a14.port_b_data_out_clock = "none";
defparam ram_block3a14.port_b_data_width = 1;
defparam ram_block3a14.port_b_first_address = 0;
defparam ram_block3a14.port_b_first_bit_number = 14;
defparam ram_block3a14.port_b_last_address = 8191;
defparam ram_block3a14.port_b_logical_ram_depth = 16384;
defparam ram_block3a14.port_b_logical_ram_width = 32;
defparam ram_block3a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_read_enable_clock = "clock1";
defparam ram_block3a14.port_b_write_enable_clock = "clock1";
defparam ram_block3a14.ram_block_type = "M9K";
defparam ram_block3a14.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004007E01;
// synopsys translate_on

// Location: M9K_X51_Y42_N0
cycloneive_ram_block ram_block3a47(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a47_PORTADATAOUT_bus),
	.portbdataout(ram_block3a47_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a47.clk0_core_clock_enable = "ena0";
defparam ram_block3a47.clk1_core_clock_enable = "ena1";
defparam ram_block3a47.data_interleave_offset_in_bits = 1;
defparam ram_block3a47.data_interleave_width_in_bits = 1;
defparam ram_block3a47.init_file = "meminit.hex";
defparam ram_block3a47.init_file_layout = "port_a";
defparam ram_block3a47.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a47.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a47.operation_mode = "bidir_dual_port";
defparam ram_block3a47.port_a_address_clear = "none";
defparam ram_block3a47.port_a_address_width = 13;
defparam ram_block3a47.port_a_byte_enable_clock = "none";
defparam ram_block3a47.port_a_data_out_clear = "none";
defparam ram_block3a47.port_a_data_out_clock = "none";
defparam ram_block3a47.port_a_data_width = 1;
defparam ram_block3a47.port_a_first_address = 0;
defparam ram_block3a47.port_a_first_bit_number = 15;
defparam ram_block3a47.port_a_last_address = 8191;
defparam ram_block3a47.port_a_logical_ram_depth = 16384;
defparam ram_block3a47.port_a_logical_ram_width = 32;
defparam ram_block3a47.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_address_clear = "none";
defparam ram_block3a47.port_b_address_clock = "clock1";
defparam ram_block3a47.port_b_address_width = 13;
defparam ram_block3a47.port_b_data_in_clock = "clock1";
defparam ram_block3a47.port_b_data_out_clear = "none";
defparam ram_block3a47.port_b_data_out_clock = "none";
defparam ram_block3a47.port_b_data_width = 1;
defparam ram_block3a47.port_b_first_address = 0;
defparam ram_block3a47.port_b_first_bit_number = 15;
defparam ram_block3a47.port_b_last_address = 8191;
defparam ram_block3a47.port_b_logical_ram_depth = 16384;
defparam ram_block3a47.port_b_logical_ram_width = 32;
defparam ram_block3a47.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_read_enable_clock = "clock1";
defparam ram_block3a47.port_b_write_enable_clock = "clock1";
defparam ram_block3a47.ram_block_type = "M9K";
defparam ram_block3a47.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y41_N0
cycloneive_ram_block ram_block3a15(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a15_PORTADATAOUT_bus),
	.portbdataout(ram_block3a15_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a15.clk0_core_clock_enable = "ena0";
defparam ram_block3a15.clk1_core_clock_enable = "ena1";
defparam ram_block3a15.data_interleave_offset_in_bits = 1;
defparam ram_block3a15.data_interleave_width_in_bits = 1;
defparam ram_block3a15.init_file = "meminit.hex";
defparam ram_block3a15.init_file_layout = "port_a";
defparam ram_block3a15.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a15.operation_mode = "bidir_dual_port";
defparam ram_block3a15.port_a_address_clear = "none";
defparam ram_block3a15.port_a_address_width = 13;
defparam ram_block3a15.port_a_byte_enable_clock = "none";
defparam ram_block3a15.port_a_data_out_clear = "none";
defparam ram_block3a15.port_a_data_out_clock = "none";
defparam ram_block3a15.port_a_data_width = 1;
defparam ram_block3a15.port_a_first_address = 0;
defparam ram_block3a15.port_a_first_bit_number = 15;
defparam ram_block3a15.port_a_last_address = 8191;
defparam ram_block3a15.port_a_logical_ram_depth = 16384;
defparam ram_block3a15.port_a_logical_ram_width = 32;
defparam ram_block3a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_address_clear = "none";
defparam ram_block3a15.port_b_address_clock = "clock1";
defparam ram_block3a15.port_b_address_width = 13;
defparam ram_block3a15.port_b_data_in_clock = "clock1";
defparam ram_block3a15.port_b_data_out_clear = "none";
defparam ram_block3a15.port_b_data_out_clock = "none";
defparam ram_block3a15.port_b_data_width = 1;
defparam ram_block3a15.port_b_first_address = 0;
defparam ram_block3a15.port_b_first_bit_number = 15;
defparam ram_block3a15.port_b_last_address = 8191;
defparam ram_block3a15.port_b_logical_ram_depth = 16384;
defparam ram_block3a15.port_b_logical_ram_width = 32;
defparam ram_block3a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_read_enable_clock = "clock1";
defparam ram_block3a15.port_b_write_enable_clock = "clock1";
defparam ram_block3a15.ram_block_type = "M9K";
defparam ram_block3a15.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004000901;
// synopsys translate_on

// Location: M9K_X51_Y39_N0
cycloneive_ram_block ram_block3a48(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a48_PORTADATAOUT_bus),
	.portbdataout(ram_block3a48_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a48.clk0_core_clock_enable = "ena0";
defparam ram_block3a48.clk1_core_clock_enable = "ena1";
defparam ram_block3a48.data_interleave_offset_in_bits = 1;
defparam ram_block3a48.data_interleave_width_in_bits = 1;
defparam ram_block3a48.init_file = "meminit.hex";
defparam ram_block3a48.init_file_layout = "port_a";
defparam ram_block3a48.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a48.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a48.operation_mode = "bidir_dual_port";
defparam ram_block3a48.port_a_address_clear = "none";
defparam ram_block3a48.port_a_address_width = 13;
defparam ram_block3a48.port_a_byte_enable_clock = "none";
defparam ram_block3a48.port_a_data_out_clear = "none";
defparam ram_block3a48.port_a_data_out_clock = "none";
defparam ram_block3a48.port_a_data_width = 1;
defparam ram_block3a48.port_a_first_address = 0;
defparam ram_block3a48.port_a_first_bit_number = 16;
defparam ram_block3a48.port_a_last_address = 8191;
defparam ram_block3a48.port_a_logical_ram_depth = 16384;
defparam ram_block3a48.port_a_logical_ram_width = 32;
defparam ram_block3a48.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_address_clear = "none";
defparam ram_block3a48.port_b_address_clock = "clock1";
defparam ram_block3a48.port_b_address_width = 13;
defparam ram_block3a48.port_b_data_in_clock = "clock1";
defparam ram_block3a48.port_b_data_out_clear = "none";
defparam ram_block3a48.port_b_data_out_clock = "none";
defparam ram_block3a48.port_b_data_width = 1;
defparam ram_block3a48.port_b_first_address = 0;
defparam ram_block3a48.port_b_first_bit_number = 16;
defparam ram_block3a48.port_b_last_address = 8191;
defparam ram_block3a48.port_b_logical_ram_depth = 16384;
defparam ram_block3a48.port_b_logical_ram_width = 32;
defparam ram_block3a48.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_read_enable_clock = "clock1";
defparam ram_block3a48.port_b_write_enable_clock = "clock1";
defparam ram_block3a48.ram_block_type = "M9K";
defparam ram_block3a48.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y37_N0
cycloneive_ram_block ram_block3a16(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a16_PORTADATAOUT_bus),
	.portbdataout(ram_block3a16_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a16.clk0_core_clock_enable = "ena0";
defparam ram_block3a16.clk1_core_clock_enable = "ena1";
defparam ram_block3a16.data_interleave_offset_in_bits = 1;
defparam ram_block3a16.data_interleave_width_in_bits = 1;
defparam ram_block3a16.init_file = "meminit.hex";
defparam ram_block3a16.init_file_layout = "port_a";
defparam ram_block3a16.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a16.operation_mode = "bidir_dual_port";
defparam ram_block3a16.port_a_address_clear = "none";
defparam ram_block3a16.port_a_address_width = 13;
defparam ram_block3a16.port_a_byte_enable_clock = "none";
defparam ram_block3a16.port_a_data_out_clear = "none";
defparam ram_block3a16.port_a_data_out_clock = "none";
defparam ram_block3a16.port_a_data_width = 1;
defparam ram_block3a16.port_a_first_address = 0;
defparam ram_block3a16.port_a_first_bit_number = 16;
defparam ram_block3a16.port_a_last_address = 8191;
defparam ram_block3a16.port_a_logical_ram_depth = 16384;
defparam ram_block3a16.port_a_logical_ram_width = 32;
defparam ram_block3a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_address_clear = "none";
defparam ram_block3a16.port_b_address_clock = "clock1";
defparam ram_block3a16.port_b_address_width = 13;
defparam ram_block3a16.port_b_data_in_clock = "clock1";
defparam ram_block3a16.port_b_data_out_clear = "none";
defparam ram_block3a16.port_b_data_out_clock = "none";
defparam ram_block3a16.port_b_data_width = 1;
defparam ram_block3a16.port_b_first_address = 0;
defparam ram_block3a16.port_b_first_bit_number = 16;
defparam ram_block3a16.port_b_last_address = 8191;
defparam ram_block3a16.port_b_logical_ram_depth = 16384;
defparam ram_block3a16.port_b_logical_ram_width = 32;
defparam ram_block3a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_read_enable_clock = "clock1";
defparam ram_block3a16.port_b_write_enable_clock = "clock1";
defparam ram_block3a16.ram_block_type = "M9K";
defparam ram_block3a16.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005558145;
// synopsys translate_on

// Location: M9K_X51_Y34_N0
cycloneive_ram_block ram_block3a49(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a49_PORTADATAOUT_bus),
	.portbdataout(ram_block3a49_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a49.clk0_core_clock_enable = "ena0";
defparam ram_block3a49.clk1_core_clock_enable = "ena1";
defparam ram_block3a49.data_interleave_offset_in_bits = 1;
defparam ram_block3a49.data_interleave_width_in_bits = 1;
defparam ram_block3a49.init_file = "meminit.hex";
defparam ram_block3a49.init_file_layout = "port_a";
defparam ram_block3a49.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a49.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a49.operation_mode = "bidir_dual_port";
defparam ram_block3a49.port_a_address_clear = "none";
defparam ram_block3a49.port_a_address_width = 13;
defparam ram_block3a49.port_a_byte_enable_clock = "none";
defparam ram_block3a49.port_a_data_out_clear = "none";
defparam ram_block3a49.port_a_data_out_clock = "none";
defparam ram_block3a49.port_a_data_width = 1;
defparam ram_block3a49.port_a_first_address = 0;
defparam ram_block3a49.port_a_first_bit_number = 17;
defparam ram_block3a49.port_a_last_address = 8191;
defparam ram_block3a49.port_a_logical_ram_depth = 16384;
defparam ram_block3a49.port_a_logical_ram_width = 32;
defparam ram_block3a49.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_address_clear = "none";
defparam ram_block3a49.port_b_address_clock = "clock1";
defparam ram_block3a49.port_b_address_width = 13;
defparam ram_block3a49.port_b_data_in_clock = "clock1";
defparam ram_block3a49.port_b_data_out_clear = "none";
defparam ram_block3a49.port_b_data_out_clock = "none";
defparam ram_block3a49.port_b_data_width = 1;
defparam ram_block3a49.port_b_first_address = 0;
defparam ram_block3a49.port_b_first_bit_number = 17;
defparam ram_block3a49.port_b_last_address = 8191;
defparam ram_block3a49.port_b_logical_ram_depth = 16384;
defparam ram_block3a49.port_b_logical_ram_width = 32;
defparam ram_block3a49.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_read_enable_clock = "clock1";
defparam ram_block3a49.port_b_write_enable_clock = "clock1";
defparam ram_block3a49.ram_block_type = "M9K";
defparam ram_block3a49.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y37_N0
cycloneive_ram_block ram_block3a17(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a17_PORTADATAOUT_bus),
	.portbdataout(ram_block3a17_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a17.clk0_core_clock_enable = "ena0";
defparam ram_block3a17.clk1_core_clock_enable = "ena1";
defparam ram_block3a17.data_interleave_offset_in_bits = 1;
defparam ram_block3a17.data_interleave_width_in_bits = 1;
defparam ram_block3a17.init_file = "meminit.hex";
defparam ram_block3a17.init_file_layout = "port_a";
defparam ram_block3a17.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a17.operation_mode = "bidir_dual_port";
defparam ram_block3a17.port_a_address_clear = "none";
defparam ram_block3a17.port_a_address_width = 13;
defparam ram_block3a17.port_a_byte_enable_clock = "none";
defparam ram_block3a17.port_a_data_out_clear = "none";
defparam ram_block3a17.port_a_data_out_clock = "none";
defparam ram_block3a17.port_a_data_width = 1;
defparam ram_block3a17.port_a_first_address = 0;
defparam ram_block3a17.port_a_first_bit_number = 17;
defparam ram_block3a17.port_a_last_address = 8191;
defparam ram_block3a17.port_a_logical_ram_depth = 16384;
defparam ram_block3a17.port_a_logical_ram_width = 32;
defparam ram_block3a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_address_clear = "none";
defparam ram_block3a17.port_b_address_clock = "clock1";
defparam ram_block3a17.port_b_address_width = 13;
defparam ram_block3a17.port_b_data_in_clock = "clock1";
defparam ram_block3a17.port_b_data_out_clear = "none";
defparam ram_block3a17.port_b_data_out_clock = "none";
defparam ram_block3a17.port_b_data_width = 1;
defparam ram_block3a17.port_b_first_address = 0;
defparam ram_block3a17.port_b_first_bit_number = 17;
defparam ram_block3a17.port_b_last_address = 8191;
defparam ram_block3a17.port_b_logical_ram_depth = 16384;
defparam ram_block3a17.port_b_logical_ram_width = 32;
defparam ram_block3a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_read_enable_clock = "clock1";
defparam ram_block3a17.port_b_write_enable_clock = "clock1";
defparam ram_block3a17.ram_block_type = "M9K";
defparam ram_block3a17.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005994FBA;
// synopsys translate_on

// Location: M9K_X51_Y26_N0
cycloneive_ram_block ram_block3a50(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a50_PORTADATAOUT_bus),
	.portbdataout(ram_block3a50_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a50.clk0_core_clock_enable = "ena0";
defparam ram_block3a50.clk1_core_clock_enable = "ena1";
defparam ram_block3a50.data_interleave_offset_in_bits = 1;
defparam ram_block3a50.data_interleave_width_in_bits = 1;
defparam ram_block3a50.init_file = "meminit.hex";
defparam ram_block3a50.init_file_layout = "port_a";
defparam ram_block3a50.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a50.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a50.operation_mode = "bidir_dual_port";
defparam ram_block3a50.port_a_address_clear = "none";
defparam ram_block3a50.port_a_address_width = 13;
defparam ram_block3a50.port_a_byte_enable_clock = "none";
defparam ram_block3a50.port_a_data_out_clear = "none";
defparam ram_block3a50.port_a_data_out_clock = "none";
defparam ram_block3a50.port_a_data_width = 1;
defparam ram_block3a50.port_a_first_address = 0;
defparam ram_block3a50.port_a_first_bit_number = 18;
defparam ram_block3a50.port_a_last_address = 8191;
defparam ram_block3a50.port_a_logical_ram_depth = 16384;
defparam ram_block3a50.port_a_logical_ram_width = 32;
defparam ram_block3a50.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_address_clear = "none";
defparam ram_block3a50.port_b_address_clock = "clock1";
defparam ram_block3a50.port_b_address_width = 13;
defparam ram_block3a50.port_b_data_in_clock = "clock1";
defparam ram_block3a50.port_b_data_out_clear = "none";
defparam ram_block3a50.port_b_data_out_clock = "none";
defparam ram_block3a50.port_b_data_width = 1;
defparam ram_block3a50.port_b_first_address = 0;
defparam ram_block3a50.port_b_first_bit_number = 18;
defparam ram_block3a50.port_b_last_address = 8191;
defparam ram_block3a50.port_b_logical_ram_depth = 16384;
defparam ram_block3a50.port_b_logical_ram_width = 32;
defparam ram_block3a50.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_read_enable_clock = "clock1";
defparam ram_block3a50.port_b_write_enable_clock = "clock1";
defparam ram_block3a50.ram_block_type = "M9K";
defparam ram_block3a50.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y40_N0
cycloneive_ram_block ram_block3a18(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a18_PORTADATAOUT_bus),
	.portbdataout(ram_block3a18_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a18.clk0_core_clock_enable = "ena0";
defparam ram_block3a18.clk1_core_clock_enable = "ena1";
defparam ram_block3a18.data_interleave_offset_in_bits = 1;
defparam ram_block3a18.data_interleave_width_in_bits = 1;
defparam ram_block3a18.init_file = "meminit.hex";
defparam ram_block3a18.init_file_layout = "port_a";
defparam ram_block3a18.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a18.operation_mode = "bidir_dual_port";
defparam ram_block3a18.port_a_address_clear = "none";
defparam ram_block3a18.port_a_address_width = 13;
defparam ram_block3a18.port_a_byte_enable_clock = "none";
defparam ram_block3a18.port_a_data_out_clear = "none";
defparam ram_block3a18.port_a_data_out_clock = "none";
defparam ram_block3a18.port_a_data_width = 1;
defparam ram_block3a18.port_a_first_address = 0;
defparam ram_block3a18.port_a_first_bit_number = 18;
defparam ram_block3a18.port_a_last_address = 8191;
defparam ram_block3a18.port_a_logical_ram_depth = 16384;
defparam ram_block3a18.port_a_logical_ram_width = 32;
defparam ram_block3a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_address_clear = "none";
defparam ram_block3a18.port_b_address_clock = "clock1";
defparam ram_block3a18.port_b_address_width = 13;
defparam ram_block3a18.port_b_data_in_clock = "clock1";
defparam ram_block3a18.port_b_data_out_clear = "none";
defparam ram_block3a18.port_b_data_out_clock = "none";
defparam ram_block3a18.port_b_data_width = 1;
defparam ram_block3a18.port_b_first_address = 0;
defparam ram_block3a18.port_b_first_bit_number = 18;
defparam ram_block3a18.port_b_last_address = 8191;
defparam ram_block3a18.port_b_logical_ram_depth = 16384;
defparam ram_block3a18.port_b_logical_ram_width = 32;
defparam ram_block3a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_read_enable_clock = "clock1";
defparam ram_block3a18.port_b_write_enable_clock = "clock1";
defparam ram_block3a18.ram_block_type = "M9K";
defparam ram_block3a18.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000061E814C;
// synopsys translate_on

// Location: M9K_X64_Y38_N0
cycloneive_ram_block ram_block3a51(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a51_PORTADATAOUT_bus),
	.portbdataout(ram_block3a51_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a51.clk0_core_clock_enable = "ena0";
defparam ram_block3a51.clk1_core_clock_enable = "ena1";
defparam ram_block3a51.data_interleave_offset_in_bits = 1;
defparam ram_block3a51.data_interleave_width_in_bits = 1;
defparam ram_block3a51.init_file = "meminit.hex";
defparam ram_block3a51.init_file_layout = "port_a";
defparam ram_block3a51.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a51.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a51.operation_mode = "bidir_dual_port";
defparam ram_block3a51.port_a_address_clear = "none";
defparam ram_block3a51.port_a_address_width = 13;
defparam ram_block3a51.port_a_byte_enable_clock = "none";
defparam ram_block3a51.port_a_data_out_clear = "none";
defparam ram_block3a51.port_a_data_out_clock = "none";
defparam ram_block3a51.port_a_data_width = 1;
defparam ram_block3a51.port_a_first_address = 0;
defparam ram_block3a51.port_a_first_bit_number = 19;
defparam ram_block3a51.port_a_last_address = 8191;
defparam ram_block3a51.port_a_logical_ram_depth = 16384;
defparam ram_block3a51.port_a_logical_ram_width = 32;
defparam ram_block3a51.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_address_clear = "none";
defparam ram_block3a51.port_b_address_clock = "clock1";
defparam ram_block3a51.port_b_address_width = 13;
defparam ram_block3a51.port_b_data_in_clock = "clock1";
defparam ram_block3a51.port_b_data_out_clear = "none";
defparam ram_block3a51.port_b_data_out_clock = "none";
defparam ram_block3a51.port_b_data_width = 1;
defparam ram_block3a51.port_b_first_address = 0;
defparam ram_block3a51.port_b_first_bit_number = 19;
defparam ram_block3a51.port_b_last_address = 8191;
defparam ram_block3a51.port_b_logical_ram_depth = 16384;
defparam ram_block3a51.port_b_logical_ram_width = 32;
defparam ram_block3a51.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_read_enable_clock = "clock1";
defparam ram_block3a51.port_b_write_enable_clock = "clock1";
defparam ram_block3a51.ram_block_type = "M9K";
defparam ram_block3a51.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y38_N0
cycloneive_ram_block ram_block3a19(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a19_PORTADATAOUT_bus),
	.portbdataout(ram_block3a19_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a19.clk0_core_clock_enable = "ena0";
defparam ram_block3a19.clk1_core_clock_enable = "ena1";
defparam ram_block3a19.data_interleave_offset_in_bits = 1;
defparam ram_block3a19.data_interleave_width_in_bits = 1;
defparam ram_block3a19.init_file = "meminit.hex";
defparam ram_block3a19.init_file_layout = "port_a";
defparam ram_block3a19.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a19.operation_mode = "bidir_dual_port";
defparam ram_block3a19.port_a_address_clear = "none";
defparam ram_block3a19.port_a_address_width = 13;
defparam ram_block3a19.port_a_byte_enable_clock = "none";
defparam ram_block3a19.port_a_data_out_clear = "none";
defparam ram_block3a19.port_a_data_out_clock = "none";
defparam ram_block3a19.port_a_data_width = 1;
defparam ram_block3a19.port_a_first_address = 0;
defparam ram_block3a19.port_a_first_bit_number = 19;
defparam ram_block3a19.port_a_last_address = 8191;
defparam ram_block3a19.port_a_logical_ram_depth = 16384;
defparam ram_block3a19.port_a_logical_ram_width = 32;
defparam ram_block3a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_address_clear = "none";
defparam ram_block3a19.port_b_address_clock = "clock1";
defparam ram_block3a19.port_b_address_width = 13;
defparam ram_block3a19.port_b_data_in_clock = "clock1";
defparam ram_block3a19.port_b_data_out_clear = "none";
defparam ram_block3a19.port_b_data_out_clock = "none";
defparam ram_block3a19.port_b_data_width = 1;
defparam ram_block3a19.port_b_first_address = 0;
defparam ram_block3a19.port_b_first_bit_number = 19;
defparam ram_block3a19.port_b_last_address = 8191;
defparam ram_block3a19.port_b_logical_ram_depth = 16384;
defparam ram_block3a19.port_b_logical_ram_width = 32;
defparam ram_block3a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_read_enable_clock = "clock1";
defparam ram_block3a19.port_b_write_enable_clock = "clock1";
defparam ram_block3a19.ram_block_type = "M9K";
defparam ram_block3a19.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007E08800;
// synopsys translate_on

// Location: M9K_X64_Y25_N0
cycloneive_ram_block ram_block3a52(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a52_PORTADATAOUT_bus),
	.portbdataout(ram_block3a52_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a52.clk0_core_clock_enable = "ena0";
defparam ram_block3a52.clk1_core_clock_enable = "ena1";
defparam ram_block3a52.data_interleave_offset_in_bits = 1;
defparam ram_block3a52.data_interleave_width_in_bits = 1;
defparam ram_block3a52.init_file = "meminit.hex";
defparam ram_block3a52.init_file_layout = "port_a";
defparam ram_block3a52.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a52.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a52.operation_mode = "bidir_dual_port";
defparam ram_block3a52.port_a_address_clear = "none";
defparam ram_block3a52.port_a_address_width = 13;
defparam ram_block3a52.port_a_byte_enable_clock = "none";
defparam ram_block3a52.port_a_data_out_clear = "none";
defparam ram_block3a52.port_a_data_out_clock = "none";
defparam ram_block3a52.port_a_data_width = 1;
defparam ram_block3a52.port_a_first_address = 0;
defparam ram_block3a52.port_a_first_bit_number = 20;
defparam ram_block3a52.port_a_last_address = 8191;
defparam ram_block3a52.port_a_logical_ram_depth = 16384;
defparam ram_block3a52.port_a_logical_ram_width = 32;
defparam ram_block3a52.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_address_clear = "none";
defparam ram_block3a52.port_b_address_clock = "clock1";
defparam ram_block3a52.port_b_address_width = 13;
defparam ram_block3a52.port_b_data_in_clock = "clock1";
defparam ram_block3a52.port_b_data_out_clear = "none";
defparam ram_block3a52.port_b_data_out_clock = "none";
defparam ram_block3a52.port_b_data_width = 1;
defparam ram_block3a52.port_b_first_address = 0;
defparam ram_block3a52.port_b_first_bit_number = 20;
defparam ram_block3a52.port_b_last_address = 8191;
defparam ram_block3a52.port_b_logical_ram_depth = 16384;
defparam ram_block3a52.port_b_logical_ram_width = 32;
defparam ram_block3a52.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_read_enable_clock = "clock1";
defparam ram_block3a52.port_b_write_enable_clock = "clock1";
defparam ram_block3a52.ram_block_type = "M9K";
defparam ram_block3a52.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y22_N0
cycloneive_ram_block ram_block3a20(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a20_PORTADATAOUT_bus),
	.portbdataout(ram_block3a20_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a20.clk0_core_clock_enable = "ena0";
defparam ram_block3a20.clk1_core_clock_enable = "ena1";
defparam ram_block3a20.data_interleave_offset_in_bits = 1;
defparam ram_block3a20.data_interleave_width_in_bits = 1;
defparam ram_block3a20.init_file = "meminit.hex";
defparam ram_block3a20.init_file_layout = "port_a";
defparam ram_block3a20.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a20.operation_mode = "bidir_dual_port";
defparam ram_block3a20.port_a_address_clear = "none";
defparam ram_block3a20.port_a_address_width = 13;
defparam ram_block3a20.port_a_byte_enable_clock = "none";
defparam ram_block3a20.port_a_data_out_clear = "none";
defparam ram_block3a20.port_a_data_out_clock = "none";
defparam ram_block3a20.port_a_data_width = 1;
defparam ram_block3a20.port_a_first_address = 0;
defparam ram_block3a20.port_a_first_bit_number = 20;
defparam ram_block3a20.port_a_last_address = 8191;
defparam ram_block3a20.port_a_logical_ram_depth = 16384;
defparam ram_block3a20.port_a_logical_ram_width = 32;
defparam ram_block3a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_address_clear = "none";
defparam ram_block3a20.port_b_address_clock = "clock1";
defparam ram_block3a20.port_b_address_width = 13;
defparam ram_block3a20.port_b_data_in_clock = "clock1";
defparam ram_block3a20.port_b_data_out_clear = "none";
defparam ram_block3a20.port_b_data_out_clock = "none";
defparam ram_block3a20.port_b_data_width = 1;
defparam ram_block3a20.port_b_first_address = 0;
defparam ram_block3a20.port_b_first_bit_number = 20;
defparam ram_block3a20.port_b_last_address = 8191;
defparam ram_block3a20.port_b_logical_ram_depth = 16384;
defparam ram_block3a20.port_b_logical_ram_width = 32;
defparam ram_block3a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_read_enable_clock = "clock1";
defparam ram_block3a20.port_b_write_enable_clock = "clock1";
defparam ram_block3a20.ram_block_type = "M9K";
defparam ram_block3a20.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000400000C;
// synopsys translate_on

// Location: M9K_X51_Y24_N0
cycloneive_ram_block ram_block3a53(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a53_PORTADATAOUT_bus),
	.portbdataout(ram_block3a53_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a53.clk0_core_clock_enable = "ena0";
defparam ram_block3a53.clk1_core_clock_enable = "ena1";
defparam ram_block3a53.data_interleave_offset_in_bits = 1;
defparam ram_block3a53.data_interleave_width_in_bits = 1;
defparam ram_block3a53.init_file = "meminit.hex";
defparam ram_block3a53.init_file_layout = "port_a";
defparam ram_block3a53.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a53.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a53.operation_mode = "bidir_dual_port";
defparam ram_block3a53.port_a_address_clear = "none";
defparam ram_block3a53.port_a_address_width = 13;
defparam ram_block3a53.port_a_byte_enable_clock = "none";
defparam ram_block3a53.port_a_data_out_clear = "none";
defparam ram_block3a53.port_a_data_out_clock = "none";
defparam ram_block3a53.port_a_data_width = 1;
defparam ram_block3a53.port_a_first_address = 0;
defparam ram_block3a53.port_a_first_bit_number = 21;
defparam ram_block3a53.port_a_last_address = 8191;
defparam ram_block3a53.port_a_logical_ram_depth = 16384;
defparam ram_block3a53.port_a_logical_ram_width = 32;
defparam ram_block3a53.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_address_clear = "none";
defparam ram_block3a53.port_b_address_clock = "clock1";
defparam ram_block3a53.port_b_address_width = 13;
defparam ram_block3a53.port_b_data_in_clock = "clock1";
defparam ram_block3a53.port_b_data_out_clear = "none";
defparam ram_block3a53.port_b_data_out_clock = "none";
defparam ram_block3a53.port_b_data_width = 1;
defparam ram_block3a53.port_b_first_address = 0;
defparam ram_block3a53.port_b_first_bit_number = 21;
defparam ram_block3a53.port_b_last_address = 8191;
defparam ram_block3a53.port_b_logical_ram_depth = 16384;
defparam ram_block3a53.port_b_logical_ram_width = 32;
defparam ram_block3a53.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_read_enable_clock = "clock1";
defparam ram_block3a53.port_b_write_enable_clock = "clock1";
defparam ram_block3a53.ram_block_type = "M9K";
defparam ram_block3a53.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y27_N0
cycloneive_ram_block ram_block3a21(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a21_PORTADATAOUT_bus),
	.portbdataout(ram_block3a21_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a21.clk0_core_clock_enable = "ena0";
defparam ram_block3a21.clk1_core_clock_enable = "ena1";
defparam ram_block3a21.data_interleave_offset_in_bits = 1;
defparam ram_block3a21.data_interleave_width_in_bits = 1;
defparam ram_block3a21.init_file = "meminit.hex";
defparam ram_block3a21.init_file_layout = "port_a";
defparam ram_block3a21.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a21.operation_mode = "bidir_dual_port";
defparam ram_block3a21.port_a_address_clear = "none";
defparam ram_block3a21.port_a_address_width = 13;
defparam ram_block3a21.port_a_byte_enable_clock = "none";
defparam ram_block3a21.port_a_data_out_clear = "none";
defparam ram_block3a21.port_a_data_out_clock = "none";
defparam ram_block3a21.port_a_data_width = 1;
defparam ram_block3a21.port_a_first_address = 0;
defparam ram_block3a21.port_a_first_bit_number = 21;
defparam ram_block3a21.port_a_last_address = 8191;
defparam ram_block3a21.port_a_logical_ram_depth = 16384;
defparam ram_block3a21.port_a_logical_ram_width = 32;
defparam ram_block3a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_address_clear = "none";
defparam ram_block3a21.port_b_address_clock = "clock1";
defparam ram_block3a21.port_b_address_width = 13;
defparam ram_block3a21.port_b_data_in_clock = "clock1";
defparam ram_block3a21.port_b_data_out_clear = "none";
defparam ram_block3a21.port_b_data_out_clock = "none";
defparam ram_block3a21.port_b_data_width = 1;
defparam ram_block3a21.port_b_first_address = 0;
defparam ram_block3a21.port_b_first_bit_number = 21;
defparam ram_block3a21.port_b_last_address = 8191;
defparam ram_block3a21.port_b_logical_ram_depth = 16384;
defparam ram_block3a21.port_b_logical_ram_width = 32;
defparam ram_block3a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_read_enable_clock = "clock1";
defparam ram_block3a21.port_b_write_enable_clock = "clock1";
defparam ram_block3a21.ram_block_type = "M9K";
defparam ram_block3a21.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FF7DF0;
// synopsys translate_on

// Location: M9K_X51_Y33_N0
cycloneive_ram_block ram_block3a54(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a54_PORTADATAOUT_bus),
	.portbdataout(ram_block3a54_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a54.clk0_core_clock_enable = "ena0";
defparam ram_block3a54.clk1_core_clock_enable = "ena1";
defparam ram_block3a54.data_interleave_offset_in_bits = 1;
defparam ram_block3a54.data_interleave_width_in_bits = 1;
defparam ram_block3a54.init_file = "meminit.hex";
defparam ram_block3a54.init_file_layout = "port_a";
defparam ram_block3a54.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a54.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a54.operation_mode = "bidir_dual_port";
defparam ram_block3a54.port_a_address_clear = "none";
defparam ram_block3a54.port_a_address_width = 13;
defparam ram_block3a54.port_a_byte_enable_clock = "none";
defparam ram_block3a54.port_a_data_out_clear = "none";
defparam ram_block3a54.port_a_data_out_clock = "none";
defparam ram_block3a54.port_a_data_width = 1;
defparam ram_block3a54.port_a_first_address = 0;
defparam ram_block3a54.port_a_first_bit_number = 22;
defparam ram_block3a54.port_a_last_address = 8191;
defparam ram_block3a54.port_a_logical_ram_depth = 16384;
defparam ram_block3a54.port_a_logical_ram_width = 32;
defparam ram_block3a54.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_address_clear = "none";
defparam ram_block3a54.port_b_address_clock = "clock1";
defparam ram_block3a54.port_b_address_width = 13;
defparam ram_block3a54.port_b_data_in_clock = "clock1";
defparam ram_block3a54.port_b_data_out_clear = "none";
defparam ram_block3a54.port_b_data_out_clock = "none";
defparam ram_block3a54.port_b_data_width = 1;
defparam ram_block3a54.port_b_first_address = 0;
defparam ram_block3a54.port_b_first_bit_number = 22;
defparam ram_block3a54.port_b_last_address = 8191;
defparam ram_block3a54.port_b_logical_ram_depth = 16384;
defparam ram_block3a54.port_b_logical_ram_width = 32;
defparam ram_block3a54.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_read_enable_clock = "clock1";
defparam ram_block3a54.port_b_write_enable_clock = "clock1";
defparam ram_block3a54.ram_block_type = "M9K";
defparam ram_block3a54.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y31_N0
cycloneive_ram_block ram_block3a22(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a22_PORTADATAOUT_bus),
	.portbdataout(ram_block3a22_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a22.clk0_core_clock_enable = "ena0";
defparam ram_block3a22.clk1_core_clock_enable = "ena1";
defparam ram_block3a22.data_interleave_offset_in_bits = 1;
defparam ram_block3a22.data_interleave_width_in_bits = 1;
defparam ram_block3a22.init_file = "meminit.hex";
defparam ram_block3a22.init_file_layout = "port_a";
defparam ram_block3a22.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a22.operation_mode = "bidir_dual_port";
defparam ram_block3a22.port_a_address_clear = "none";
defparam ram_block3a22.port_a_address_width = 13;
defparam ram_block3a22.port_a_byte_enable_clock = "none";
defparam ram_block3a22.port_a_data_out_clear = "none";
defparam ram_block3a22.port_a_data_out_clock = "none";
defparam ram_block3a22.port_a_data_width = 1;
defparam ram_block3a22.port_a_first_address = 0;
defparam ram_block3a22.port_a_first_bit_number = 22;
defparam ram_block3a22.port_a_last_address = 8191;
defparam ram_block3a22.port_a_logical_ram_depth = 16384;
defparam ram_block3a22.port_a_logical_ram_width = 32;
defparam ram_block3a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_address_clear = "none";
defparam ram_block3a22.port_b_address_clock = "clock1";
defparam ram_block3a22.port_b_address_width = 13;
defparam ram_block3a22.port_b_data_in_clock = "clock1";
defparam ram_block3a22.port_b_data_out_clear = "none";
defparam ram_block3a22.port_b_data_out_clock = "none";
defparam ram_block3a22.port_b_data_width = 1;
defparam ram_block3a22.port_b_first_address = 0;
defparam ram_block3a22.port_b_first_bit_number = 22;
defparam ram_block3a22.port_b_last_address = 8191;
defparam ram_block3a22.port_b_logical_ram_depth = 16384;
defparam ram_block3a22.port_b_logical_ram_width = 32;
defparam ram_block3a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_read_enable_clock = "clock1";
defparam ram_block3a22.port_b_write_enable_clock = "clock1";
defparam ram_block3a22.ram_block_type = "M9K";
defparam ram_block3a22.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004008100;
// synopsys translate_on

// Location: M9K_X64_Y30_N0
cycloneive_ram_block ram_block3a55(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a55_PORTADATAOUT_bus),
	.portbdataout(ram_block3a55_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a55.clk0_core_clock_enable = "ena0";
defparam ram_block3a55.clk1_core_clock_enable = "ena1";
defparam ram_block3a55.data_interleave_offset_in_bits = 1;
defparam ram_block3a55.data_interleave_width_in_bits = 1;
defparam ram_block3a55.init_file = "meminit.hex";
defparam ram_block3a55.init_file_layout = "port_a";
defparam ram_block3a55.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a55.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a55.operation_mode = "bidir_dual_port";
defparam ram_block3a55.port_a_address_clear = "none";
defparam ram_block3a55.port_a_address_width = 13;
defparam ram_block3a55.port_a_byte_enable_clock = "none";
defparam ram_block3a55.port_a_data_out_clear = "none";
defparam ram_block3a55.port_a_data_out_clock = "none";
defparam ram_block3a55.port_a_data_width = 1;
defparam ram_block3a55.port_a_first_address = 0;
defparam ram_block3a55.port_a_first_bit_number = 23;
defparam ram_block3a55.port_a_last_address = 8191;
defparam ram_block3a55.port_a_logical_ram_depth = 16384;
defparam ram_block3a55.port_a_logical_ram_width = 32;
defparam ram_block3a55.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_address_clear = "none";
defparam ram_block3a55.port_b_address_clock = "clock1";
defparam ram_block3a55.port_b_address_width = 13;
defparam ram_block3a55.port_b_data_in_clock = "clock1";
defparam ram_block3a55.port_b_data_out_clear = "none";
defparam ram_block3a55.port_b_data_out_clock = "none";
defparam ram_block3a55.port_b_data_width = 1;
defparam ram_block3a55.port_b_first_address = 0;
defparam ram_block3a55.port_b_first_bit_number = 23;
defparam ram_block3a55.port_b_last_address = 8191;
defparam ram_block3a55.port_b_logical_ram_depth = 16384;
defparam ram_block3a55.port_b_logical_ram_width = 32;
defparam ram_block3a55.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_read_enable_clock = "clock1";
defparam ram_block3a55.port_b_write_enable_clock = "clock1";
defparam ram_block3a55.ram_block_type = "M9K";
defparam ram_block3a55.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y34_N0
cycloneive_ram_block ram_block3a23(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a23_PORTADATAOUT_bus),
	.portbdataout(ram_block3a23_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a23.clk0_core_clock_enable = "ena0";
defparam ram_block3a23.clk1_core_clock_enable = "ena1";
defparam ram_block3a23.data_interleave_offset_in_bits = 1;
defparam ram_block3a23.data_interleave_width_in_bits = 1;
defparam ram_block3a23.init_file = "meminit.hex";
defparam ram_block3a23.init_file_layout = "port_a";
defparam ram_block3a23.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a23.operation_mode = "bidir_dual_port";
defparam ram_block3a23.port_a_address_clear = "none";
defparam ram_block3a23.port_a_address_width = 13;
defparam ram_block3a23.port_a_byte_enable_clock = "none";
defparam ram_block3a23.port_a_data_out_clear = "none";
defparam ram_block3a23.port_a_data_out_clock = "none";
defparam ram_block3a23.port_a_data_width = 1;
defparam ram_block3a23.port_a_first_address = 0;
defparam ram_block3a23.port_a_first_bit_number = 23;
defparam ram_block3a23.port_a_last_address = 8191;
defparam ram_block3a23.port_a_logical_ram_depth = 16384;
defparam ram_block3a23.port_a_logical_ram_width = 32;
defparam ram_block3a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_address_clear = "none";
defparam ram_block3a23.port_b_address_clock = "clock1";
defparam ram_block3a23.port_b_address_width = 13;
defparam ram_block3a23.port_b_data_in_clock = "clock1";
defparam ram_block3a23.port_b_data_out_clear = "none";
defparam ram_block3a23.port_b_data_out_clock = "none";
defparam ram_block3a23.port_b_data_width = 1;
defparam ram_block3a23.port_b_first_address = 0;
defparam ram_block3a23.port_b_first_bit_number = 23;
defparam ram_block3a23.port_b_last_address = 8191;
defparam ram_block3a23.port_b_logical_ram_depth = 16384;
defparam ram_block3a23.port_b_logical_ram_width = 32;
defparam ram_block3a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_read_enable_clock = "clock1";
defparam ram_block3a23.port_b_write_enable_clock = "clock1";
defparam ram_block3a23.ram_block_type = "M9K";
defparam ram_block3a23.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FF8600;
// synopsys translate_on

// Location: M9K_X78_Y36_N0
cycloneive_ram_block ram_block3a56(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a56_PORTADATAOUT_bus),
	.portbdataout(ram_block3a56_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a56.clk0_core_clock_enable = "ena0";
defparam ram_block3a56.clk1_core_clock_enable = "ena1";
defparam ram_block3a56.data_interleave_offset_in_bits = 1;
defparam ram_block3a56.data_interleave_width_in_bits = 1;
defparam ram_block3a56.init_file = "meminit.hex";
defparam ram_block3a56.init_file_layout = "port_a";
defparam ram_block3a56.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a56.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a56.operation_mode = "bidir_dual_port";
defparam ram_block3a56.port_a_address_clear = "none";
defparam ram_block3a56.port_a_address_width = 13;
defparam ram_block3a56.port_a_byte_enable_clock = "none";
defparam ram_block3a56.port_a_data_out_clear = "none";
defparam ram_block3a56.port_a_data_out_clock = "none";
defparam ram_block3a56.port_a_data_width = 1;
defparam ram_block3a56.port_a_first_address = 0;
defparam ram_block3a56.port_a_first_bit_number = 24;
defparam ram_block3a56.port_a_last_address = 8191;
defparam ram_block3a56.port_a_logical_ram_depth = 16384;
defparam ram_block3a56.port_a_logical_ram_width = 32;
defparam ram_block3a56.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_address_clear = "none";
defparam ram_block3a56.port_b_address_clock = "clock1";
defparam ram_block3a56.port_b_address_width = 13;
defparam ram_block3a56.port_b_data_in_clock = "clock1";
defparam ram_block3a56.port_b_data_out_clear = "none";
defparam ram_block3a56.port_b_data_out_clock = "none";
defparam ram_block3a56.port_b_data_width = 1;
defparam ram_block3a56.port_b_first_address = 0;
defparam ram_block3a56.port_b_first_bit_number = 24;
defparam ram_block3a56.port_b_last_address = 8191;
defparam ram_block3a56.port_b_logical_ram_depth = 16384;
defparam ram_block3a56.port_b_logical_ram_width = 32;
defparam ram_block3a56.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_read_enable_clock = "clock1";
defparam ram_block3a56.port_b_write_enable_clock = "clock1";
defparam ram_block3a56.ram_block_type = "M9K";
defparam ram_block3a56.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y40_N0
cycloneive_ram_block ram_block3a24(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a24_PORTADATAOUT_bus),
	.portbdataout(ram_block3a24_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a24.clk0_core_clock_enable = "ena0";
defparam ram_block3a24.clk1_core_clock_enable = "ena1";
defparam ram_block3a24.data_interleave_offset_in_bits = 1;
defparam ram_block3a24.data_interleave_width_in_bits = 1;
defparam ram_block3a24.init_file = "meminit.hex";
defparam ram_block3a24.init_file_layout = "port_a";
defparam ram_block3a24.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a24.operation_mode = "bidir_dual_port";
defparam ram_block3a24.port_a_address_clear = "none";
defparam ram_block3a24.port_a_address_width = 13;
defparam ram_block3a24.port_a_byte_enable_clock = "none";
defparam ram_block3a24.port_a_data_out_clear = "none";
defparam ram_block3a24.port_a_data_out_clock = "none";
defparam ram_block3a24.port_a_data_width = 1;
defparam ram_block3a24.port_a_first_address = 0;
defparam ram_block3a24.port_a_first_bit_number = 24;
defparam ram_block3a24.port_a_last_address = 8191;
defparam ram_block3a24.port_a_logical_ram_depth = 16384;
defparam ram_block3a24.port_a_logical_ram_width = 32;
defparam ram_block3a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_address_clear = "none";
defparam ram_block3a24.port_b_address_clock = "clock1";
defparam ram_block3a24.port_b_address_width = 13;
defparam ram_block3a24.port_b_data_in_clock = "clock1";
defparam ram_block3a24.port_b_data_out_clear = "none";
defparam ram_block3a24.port_b_data_out_clock = "none";
defparam ram_block3a24.port_b_data_width = 1;
defparam ram_block3a24.port_b_first_address = 0;
defparam ram_block3a24.port_b_first_bit_number = 24;
defparam ram_block3a24.port_b_last_address = 8191;
defparam ram_block3a24.port_b_logical_ram_depth = 16384;
defparam ram_block3a24.port_b_logical_ram_width = 32;
defparam ram_block3a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_read_enable_clock = "clock1";
defparam ram_block3a24.port_b_write_enable_clock = "clock1";
defparam ram_block3a24.ram_block_type = "M9K";
defparam ram_block3a24.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004000000;
// synopsys translate_on

// Location: M9K_X78_Y34_N0
cycloneive_ram_block ram_block3a57(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a57_PORTADATAOUT_bus),
	.portbdataout(ram_block3a57_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a57.clk0_core_clock_enable = "ena0";
defparam ram_block3a57.clk1_core_clock_enable = "ena1";
defparam ram_block3a57.data_interleave_offset_in_bits = 1;
defparam ram_block3a57.data_interleave_width_in_bits = 1;
defparam ram_block3a57.init_file = "meminit.hex";
defparam ram_block3a57.init_file_layout = "port_a";
defparam ram_block3a57.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a57.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a57.operation_mode = "bidir_dual_port";
defparam ram_block3a57.port_a_address_clear = "none";
defparam ram_block3a57.port_a_address_width = 13;
defparam ram_block3a57.port_a_byte_enable_clock = "none";
defparam ram_block3a57.port_a_data_out_clear = "none";
defparam ram_block3a57.port_a_data_out_clock = "none";
defparam ram_block3a57.port_a_data_width = 1;
defparam ram_block3a57.port_a_first_address = 0;
defparam ram_block3a57.port_a_first_bit_number = 25;
defparam ram_block3a57.port_a_last_address = 8191;
defparam ram_block3a57.port_a_logical_ram_depth = 16384;
defparam ram_block3a57.port_a_logical_ram_width = 32;
defparam ram_block3a57.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_address_clear = "none";
defparam ram_block3a57.port_b_address_clock = "clock1";
defparam ram_block3a57.port_b_address_width = 13;
defparam ram_block3a57.port_b_data_in_clock = "clock1";
defparam ram_block3a57.port_b_data_out_clear = "none";
defparam ram_block3a57.port_b_data_out_clock = "none";
defparam ram_block3a57.port_b_data_width = 1;
defparam ram_block3a57.port_b_first_address = 0;
defparam ram_block3a57.port_b_first_bit_number = 25;
defparam ram_block3a57.port_b_last_address = 8191;
defparam ram_block3a57.port_b_logical_ram_depth = 16384;
defparam ram_block3a57.port_b_logical_ram_width = 32;
defparam ram_block3a57.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_read_enable_clock = "clock1";
defparam ram_block3a57.port_b_write_enable_clock = "clock1";
defparam ram_block3a57.ram_block_type = "M9K";
defparam ram_block3a57.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y23_N0
cycloneive_ram_block ram_block3a25(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a25_PORTADATAOUT_bus),
	.portbdataout(ram_block3a25_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a25.clk0_core_clock_enable = "ena0";
defparam ram_block3a25.clk1_core_clock_enable = "ena1";
defparam ram_block3a25.data_interleave_offset_in_bits = 1;
defparam ram_block3a25.data_interleave_width_in_bits = 1;
defparam ram_block3a25.init_file = "meminit.hex";
defparam ram_block3a25.init_file_layout = "port_a";
defparam ram_block3a25.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a25.operation_mode = "bidir_dual_port";
defparam ram_block3a25.port_a_address_clear = "none";
defparam ram_block3a25.port_a_address_width = 13;
defparam ram_block3a25.port_a_byte_enable_clock = "none";
defparam ram_block3a25.port_a_data_out_clear = "none";
defparam ram_block3a25.port_a_data_out_clock = "none";
defparam ram_block3a25.port_a_data_width = 1;
defparam ram_block3a25.port_a_first_address = 0;
defparam ram_block3a25.port_a_first_bit_number = 25;
defparam ram_block3a25.port_a_last_address = 8191;
defparam ram_block3a25.port_a_logical_ram_depth = 16384;
defparam ram_block3a25.port_a_logical_ram_width = 32;
defparam ram_block3a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_address_clear = "none";
defparam ram_block3a25.port_b_address_clock = "clock1";
defparam ram_block3a25.port_b_address_width = 13;
defparam ram_block3a25.port_b_data_in_clock = "clock1";
defparam ram_block3a25.port_b_data_out_clear = "none";
defparam ram_block3a25.port_b_data_out_clock = "none";
defparam ram_block3a25.port_b_data_width = 1;
defparam ram_block3a25.port_b_first_address = 0;
defparam ram_block3a25.port_b_first_bit_number = 25;
defparam ram_block3a25.port_b_last_address = 8191;
defparam ram_block3a25.port_b_logical_ram_depth = 16384;
defparam ram_block3a25.port_b_logical_ram_width = 32;
defparam ram_block3a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_read_enable_clock = "clock1";
defparam ram_block3a25.port_b_write_enable_clock = "clock1";
defparam ram_block3a25.ram_block_type = "M9K";
defparam ram_block3a25.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FF8000;
// synopsys translate_on

// Location: M9K_X64_Y39_N0
cycloneive_ram_block ram_block3a58(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a58_PORTADATAOUT_bus),
	.portbdataout(ram_block3a58_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a58.clk0_core_clock_enable = "ena0";
defparam ram_block3a58.clk1_core_clock_enable = "ena1";
defparam ram_block3a58.data_interleave_offset_in_bits = 1;
defparam ram_block3a58.data_interleave_width_in_bits = 1;
defparam ram_block3a58.init_file = "meminit.hex";
defparam ram_block3a58.init_file_layout = "port_a";
defparam ram_block3a58.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a58.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a58.operation_mode = "bidir_dual_port";
defparam ram_block3a58.port_a_address_clear = "none";
defparam ram_block3a58.port_a_address_width = 13;
defparam ram_block3a58.port_a_byte_enable_clock = "none";
defparam ram_block3a58.port_a_data_out_clear = "none";
defparam ram_block3a58.port_a_data_out_clock = "none";
defparam ram_block3a58.port_a_data_width = 1;
defparam ram_block3a58.port_a_first_address = 0;
defparam ram_block3a58.port_a_first_bit_number = 26;
defparam ram_block3a58.port_a_last_address = 8191;
defparam ram_block3a58.port_a_logical_ram_depth = 16384;
defparam ram_block3a58.port_a_logical_ram_width = 32;
defparam ram_block3a58.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_address_clear = "none";
defparam ram_block3a58.port_b_address_clock = "clock1";
defparam ram_block3a58.port_b_address_width = 13;
defparam ram_block3a58.port_b_data_in_clock = "clock1";
defparam ram_block3a58.port_b_data_out_clear = "none";
defparam ram_block3a58.port_b_data_out_clock = "none";
defparam ram_block3a58.port_b_data_width = 1;
defparam ram_block3a58.port_b_first_address = 0;
defparam ram_block3a58.port_b_first_bit_number = 26;
defparam ram_block3a58.port_b_last_address = 8191;
defparam ram_block3a58.port_b_logical_ram_depth = 16384;
defparam ram_block3a58.port_b_logical_ram_width = 32;
defparam ram_block3a58.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_read_enable_clock = "clock1";
defparam ram_block3a58.port_b_write_enable_clock = "clock1";
defparam ram_block3a58.ram_block_type = "M9K";
defparam ram_block3a58.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y35_N0
cycloneive_ram_block ram_block3a26(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a26_PORTADATAOUT_bus),
	.portbdataout(ram_block3a26_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a26.clk0_core_clock_enable = "ena0";
defparam ram_block3a26.clk1_core_clock_enable = "ena1";
defparam ram_block3a26.data_interleave_offset_in_bits = 1;
defparam ram_block3a26.data_interleave_width_in_bits = 1;
defparam ram_block3a26.init_file = "meminit.hex";
defparam ram_block3a26.init_file_layout = "port_a";
defparam ram_block3a26.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a26.operation_mode = "bidir_dual_port";
defparam ram_block3a26.port_a_address_clear = "none";
defparam ram_block3a26.port_a_address_width = 13;
defparam ram_block3a26.port_a_byte_enable_clock = "none";
defparam ram_block3a26.port_a_data_out_clear = "none";
defparam ram_block3a26.port_a_data_out_clock = "none";
defparam ram_block3a26.port_a_data_width = 1;
defparam ram_block3a26.port_a_first_address = 0;
defparam ram_block3a26.port_a_first_bit_number = 26;
defparam ram_block3a26.port_a_last_address = 8191;
defparam ram_block3a26.port_a_logical_ram_depth = 16384;
defparam ram_block3a26.port_a_logical_ram_width = 32;
defparam ram_block3a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_address_clear = "none";
defparam ram_block3a26.port_b_address_clock = "clock1";
defparam ram_block3a26.port_b_address_width = 13;
defparam ram_block3a26.port_b_data_in_clock = "clock1";
defparam ram_block3a26.port_b_data_out_clear = "none";
defparam ram_block3a26.port_b_data_out_clock = "none";
defparam ram_block3a26.port_b_data_width = 1;
defparam ram_block3a26.port_b_first_address = 0;
defparam ram_block3a26.port_b_first_bit_number = 26;
defparam ram_block3a26.port_b_last_address = 8191;
defparam ram_block3a26.port_b_logical_ram_depth = 16384;
defparam ram_block3a26.port_b_logical_ram_width = 32;
defparam ram_block3a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_read_enable_clock = "clock1";
defparam ram_block3a26.port_b_write_enable_clock = "clock1";
defparam ram_block3a26.ram_block_type = "M9K";
defparam ram_block3a26.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FF810F;
// synopsys translate_on

// Location: M9K_X64_Y33_N0
cycloneive_ram_block ram_block3a59(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a59_PORTADATAOUT_bus),
	.portbdataout(ram_block3a59_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a59.clk0_core_clock_enable = "ena0";
defparam ram_block3a59.clk1_core_clock_enable = "ena1";
defparam ram_block3a59.data_interleave_offset_in_bits = 1;
defparam ram_block3a59.data_interleave_width_in_bits = 1;
defparam ram_block3a59.init_file = "meminit.hex";
defparam ram_block3a59.init_file_layout = "port_a";
defparam ram_block3a59.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a59.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a59.operation_mode = "bidir_dual_port";
defparam ram_block3a59.port_a_address_clear = "none";
defparam ram_block3a59.port_a_address_width = 13;
defparam ram_block3a59.port_a_byte_enable_clock = "none";
defparam ram_block3a59.port_a_data_out_clear = "none";
defparam ram_block3a59.port_a_data_out_clock = "none";
defparam ram_block3a59.port_a_data_width = 1;
defparam ram_block3a59.port_a_first_address = 0;
defparam ram_block3a59.port_a_first_bit_number = 27;
defparam ram_block3a59.port_a_last_address = 8191;
defparam ram_block3a59.port_a_logical_ram_depth = 16384;
defparam ram_block3a59.port_a_logical_ram_width = 32;
defparam ram_block3a59.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_address_clear = "none";
defparam ram_block3a59.port_b_address_clock = "clock1";
defparam ram_block3a59.port_b_address_width = 13;
defparam ram_block3a59.port_b_data_in_clock = "clock1";
defparam ram_block3a59.port_b_data_out_clear = "none";
defparam ram_block3a59.port_b_data_out_clock = "none";
defparam ram_block3a59.port_b_data_width = 1;
defparam ram_block3a59.port_b_first_address = 0;
defparam ram_block3a59.port_b_first_bit_number = 27;
defparam ram_block3a59.port_b_last_address = 8191;
defparam ram_block3a59.port_b_logical_ram_depth = 16384;
defparam ram_block3a59.port_b_logical_ram_width = 32;
defparam ram_block3a59.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_read_enable_clock = "clock1";
defparam ram_block3a59.port_b_write_enable_clock = "clock1";
defparam ram_block3a59.ram_block_type = "M9K";
defparam ram_block3a59.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y36_N0
cycloneive_ram_block ram_block3a27(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a27_PORTADATAOUT_bus),
	.portbdataout(ram_block3a27_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a27.clk0_core_clock_enable = "ena0";
defparam ram_block3a27.clk1_core_clock_enable = "ena1";
defparam ram_block3a27.data_interleave_offset_in_bits = 1;
defparam ram_block3a27.data_interleave_width_in_bits = 1;
defparam ram_block3a27.init_file = "meminit.hex";
defparam ram_block3a27.init_file_layout = "port_a";
defparam ram_block3a27.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a27.operation_mode = "bidir_dual_port";
defparam ram_block3a27.port_a_address_clear = "none";
defparam ram_block3a27.port_a_address_width = 13;
defparam ram_block3a27.port_a_byte_enable_clock = "none";
defparam ram_block3a27.port_a_data_out_clear = "none";
defparam ram_block3a27.port_a_data_out_clock = "none";
defparam ram_block3a27.port_a_data_width = 1;
defparam ram_block3a27.port_a_first_address = 0;
defparam ram_block3a27.port_a_first_bit_number = 27;
defparam ram_block3a27.port_a_last_address = 8191;
defparam ram_block3a27.port_a_logical_ram_depth = 16384;
defparam ram_block3a27.port_a_logical_ram_width = 32;
defparam ram_block3a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_address_clear = "none";
defparam ram_block3a27.port_b_address_clock = "clock1";
defparam ram_block3a27.port_b_address_width = 13;
defparam ram_block3a27.port_b_data_in_clock = "clock1";
defparam ram_block3a27.port_b_data_out_clear = "none";
defparam ram_block3a27.port_b_data_out_clock = "none";
defparam ram_block3a27.port_b_data_width = 1;
defparam ram_block3a27.port_b_first_address = 0;
defparam ram_block3a27.port_b_first_bit_number = 27;
defparam ram_block3a27.port_b_last_address = 8191;
defparam ram_block3a27.port_b_logical_ram_depth = 16384;
defparam ram_block3a27.port_b_logical_ram_width = 32;
defparam ram_block3a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_read_enable_clock = "clock1";
defparam ram_block3a27.port_b_write_enable_clock = "clock1";
defparam ram_block3a27.ram_block_type = "M9K";
defparam ram_block3a27.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FF8800;
// synopsys translate_on

// Location: M9K_X51_Y36_N0
cycloneive_ram_block ram_block3a60(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a60_PORTADATAOUT_bus),
	.portbdataout(ram_block3a60_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a60.clk0_core_clock_enable = "ena0";
defparam ram_block3a60.clk1_core_clock_enable = "ena1";
defparam ram_block3a60.data_interleave_offset_in_bits = 1;
defparam ram_block3a60.data_interleave_width_in_bits = 1;
defparam ram_block3a60.init_file = "meminit.hex";
defparam ram_block3a60.init_file_layout = "port_a";
defparam ram_block3a60.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a60.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a60.operation_mode = "bidir_dual_port";
defparam ram_block3a60.port_a_address_clear = "none";
defparam ram_block3a60.port_a_address_width = 13;
defparam ram_block3a60.port_a_byte_enable_clock = "none";
defparam ram_block3a60.port_a_data_out_clear = "none";
defparam ram_block3a60.port_a_data_out_clock = "none";
defparam ram_block3a60.port_a_data_width = 1;
defparam ram_block3a60.port_a_first_address = 0;
defparam ram_block3a60.port_a_first_bit_number = 28;
defparam ram_block3a60.port_a_last_address = 8191;
defparam ram_block3a60.port_a_logical_ram_depth = 16384;
defparam ram_block3a60.port_a_logical_ram_width = 32;
defparam ram_block3a60.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_address_clear = "none";
defparam ram_block3a60.port_b_address_clock = "clock1";
defparam ram_block3a60.port_b_address_width = 13;
defparam ram_block3a60.port_b_data_in_clock = "clock1";
defparam ram_block3a60.port_b_data_out_clear = "none";
defparam ram_block3a60.port_b_data_out_clock = "none";
defparam ram_block3a60.port_b_data_width = 1;
defparam ram_block3a60.port_b_first_address = 0;
defparam ram_block3a60.port_b_first_bit_number = 28;
defparam ram_block3a60.port_b_last_address = 8191;
defparam ram_block3a60.port_b_logical_ram_depth = 16384;
defparam ram_block3a60.port_b_logical_ram_width = 32;
defparam ram_block3a60.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_read_enable_clock = "clock1";
defparam ram_block3a60.port_b_write_enable_clock = "clock1";
defparam ram_block3a60.ram_block_type = "M9K";
defparam ram_block3a60.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y32_N0
cycloneive_ram_block ram_block3a28(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a28_PORTADATAOUT_bus),
	.portbdataout(ram_block3a28_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a28.clk0_core_clock_enable = "ena0";
defparam ram_block3a28.clk1_core_clock_enable = "ena1";
defparam ram_block3a28.data_interleave_offset_in_bits = 1;
defparam ram_block3a28.data_interleave_width_in_bits = 1;
defparam ram_block3a28.init_file = "meminit.hex";
defparam ram_block3a28.init_file_layout = "port_a";
defparam ram_block3a28.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a28.operation_mode = "bidir_dual_port";
defparam ram_block3a28.port_a_address_clear = "none";
defparam ram_block3a28.port_a_address_width = 13;
defparam ram_block3a28.port_a_byte_enable_clock = "none";
defparam ram_block3a28.port_a_data_out_clear = "none";
defparam ram_block3a28.port_a_data_out_clock = "none";
defparam ram_block3a28.port_a_data_width = 1;
defparam ram_block3a28.port_a_first_address = 0;
defparam ram_block3a28.port_a_first_bit_number = 28;
defparam ram_block3a28.port_a_last_address = 8191;
defparam ram_block3a28.port_a_logical_ram_depth = 16384;
defparam ram_block3a28.port_a_logical_ram_width = 32;
defparam ram_block3a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_address_clear = "none";
defparam ram_block3a28.port_b_address_clock = "clock1";
defparam ram_block3a28.port_b_address_width = 13;
defparam ram_block3a28.port_b_data_in_clock = "clock1";
defparam ram_block3a28.port_b_data_out_clear = "none";
defparam ram_block3a28.port_b_data_out_clock = "none";
defparam ram_block3a28.port_b_data_width = 1;
defparam ram_block3a28.port_b_first_address = 0;
defparam ram_block3a28.port_b_first_bit_number = 28;
defparam ram_block3a28.port_b_last_address = 8191;
defparam ram_block3a28.port_b_logical_ram_depth = 16384;
defparam ram_block3a28.port_b_logical_ram_width = 32;
defparam ram_block3a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_read_enable_clock = "clock1";
defparam ram_block3a28.port_b_write_enable_clock = "clock1";
defparam ram_block3a28.ram_block_type = "M9K";
defparam ram_block3a28.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000400084F;
// synopsys translate_on

// Location: M9K_X64_Y37_N0
cycloneive_ram_block ram_block3a61(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a61_PORTADATAOUT_bus),
	.portbdataout(ram_block3a61_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a61.clk0_core_clock_enable = "ena0";
defparam ram_block3a61.clk1_core_clock_enable = "ena1";
defparam ram_block3a61.data_interleave_offset_in_bits = 1;
defparam ram_block3a61.data_interleave_width_in_bits = 1;
defparam ram_block3a61.init_file = "meminit.hex";
defparam ram_block3a61.init_file_layout = "port_a";
defparam ram_block3a61.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a61.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a61.operation_mode = "bidir_dual_port";
defparam ram_block3a61.port_a_address_clear = "none";
defparam ram_block3a61.port_a_address_width = 13;
defparam ram_block3a61.port_a_byte_enable_clock = "none";
defparam ram_block3a61.port_a_data_out_clear = "none";
defparam ram_block3a61.port_a_data_out_clock = "none";
defparam ram_block3a61.port_a_data_width = 1;
defparam ram_block3a61.port_a_first_address = 0;
defparam ram_block3a61.port_a_first_bit_number = 29;
defparam ram_block3a61.port_a_last_address = 8191;
defparam ram_block3a61.port_a_logical_ram_depth = 16384;
defparam ram_block3a61.port_a_logical_ram_width = 32;
defparam ram_block3a61.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_address_clear = "none";
defparam ram_block3a61.port_b_address_clock = "clock1";
defparam ram_block3a61.port_b_address_width = 13;
defparam ram_block3a61.port_b_data_in_clock = "clock1";
defparam ram_block3a61.port_b_data_out_clear = "none";
defparam ram_block3a61.port_b_data_out_clock = "none";
defparam ram_block3a61.port_b_data_width = 1;
defparam ram_block3a61.port_b_first_address = 0;
defparam ram_block3a61.port_b_first_bit_number = 29;
defparam ram_block3a61.port_b_last_address = 8191;
defparam ram_block3a61.port_b_logical_ram_depth = 16384;
defparam ram_block3a61.port_b_logical_ram_width = 32;
defparam ram_block3a61.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_read_enable_clock = "clock1";
defparam ram_block3a61.port_b_write_enable_clock = "clock1";
defparam ram_block3a61.ram_block_type = "M9K";
defparam ram_block3a61.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y41_N0
cycloneive_ram_block ram_block3a29(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a29_PORTADATAOUT_bus),
	.portbdataout(ram_block3a29_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a29.clk0_core_clock_enable = "ena0";
defparam ram_block3a29.clk1_core_clock_enable = "ena1";
defparam ram_block3a29.data_interleave_offset_in_bits = 1;
defparam ram_block3a29.data_interleave_width_in_bits = 1;
defparam ram_block3a29.init_file = "meminit.hex";
defparam ram_block3a29.init_file_layout = "port_a";
defparam ram_block3a29.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a29.operation_mode = "bidir_dual_port";
defparam ram_block3a29.port_a_address_clear = "none";
defparam ram_block3a29.port_a_address_width = 13;
defparam ram_block3a29.port_a_byte_enable_clock = "none";
defparam ram_block3a29.port_a_data_out_clear = "none";
defparam ram_block3a29.port_a_data_out_clock = "none";
defparam ram_block3a29.port_a_data_width = 1;
defparam ram_block3a29.port_a_first_address = 0;
defparam ram_block3a29.port_a_first_bit_number = 29;
defparam ram_block3a29.port_a_last_address = 8191;
defparam ram_block3a29.port_a_logical_ram_depth = 16384;
defparam ram_block3a29.port_a_logical_ram_width = 32;
defparam ram_block3a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_address_clear = "none";
defparam ram_block3a29.port_b_address_clock = "clock1";
defparam ram_block3a29.port_b_address_width = 13;
defparam ram_block3a29.port_b_data_in_clock = "clock1";
defparam ram_block3a29.port_b_data_out_clear = "none";
defparam ram_block3a29.port_b_data_out_clock = "none";
defparam ram_block3a29.port_b_data_width = 1;
defparam ram_block3a29.port_b_first_address = 0;
defparam ram_block3a29.port_b_first_bit_number = 29;
defparam ram_block3a29.port_b_last_address = 8191;
defparam ram_block3a29.port_b_logical_ram_depth = 16384;
defparam ram_block3a29.port_b_logical_ram_width = 32;
defparam ram_block3a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_read_enable_clock = "clock1";
defparam ram_block3a29.port_b_write_enable_clock = "clock1";
defparam ram_block3a29.ram_block_type = "M9K";
defparam ram_block3a29.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FF894F;
// synopsys translate_on

// Location: M9K_X64_Y35_N0
cycloneive_ram_block ram_block3a62(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a62_PORTADATAOUT_bus),
	.portbdataout(ram_block3a62_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a62.clk0_core_clock_enable = "ena0";
defparam ram_block3a62.clk1_core_clock_enable = "ena1";
defparam ram_block3a62.data_interleave_offset_in_bits = 1;
defparam ram_block3a62.data_interleave_width_in_bits = 1;
defparam ram_block3a62.init_file = "meminit.hex";
defparam ram_block3a62.init_file_layout = "port_a";
defparam ram_block3a62.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a62.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a62.operation_mode = "bidir_dual_port";
defparam ram_block3a62.port_a_address_clear = "none";
defparam ram_block3a62.port_a_address_width = 13;
defparam ram_block3a62.port_a_byte_enable_clock = "none";
defparam ram_block3a62.port_a_data_out_clear = "none";
defparam ram_block3a62.port_a_data_out_clock = "none";
defparam ram_block3a62.port_a_data_width = 1;
defparam ram_block3a62.port_a_first_address = 0;
defparam ram_block3a62.port_a_first_bit_number = 30;
defparam ram_block3a62.port_a_last_address = 8191;
defparam ram_block3a62.port_a_logical_ram_depth = 16384;
defparam ram_block3a62.port_a_logical_ram_width = 32;
defparam ram_block3a62.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_address_clear = "none";
defparam ram_block3a62.port_b_address_clock = "clock1";
defparam ram_block3a62.port_b_address_width = 13;
defparam ram_block3a62.port_b_data_in_clock = "clock1";
defparam ram_block3a62.port_b_data_out_clear = "none";
defparam ram_block3a62.port_b_data_out_clock = "none";
defparam ram_block3a62.port_b_data_width = 1;
defparam ram_block3a62.port_b_first_address = 0;
defparam ram_block3a62.port_b_first_bit_number = 30;
defparam ram_block3a62.port_b_last_address = 8191;
defparam ram_block3a62.port_b_logical_ram_depth = 16384;
defparam ram_block3a62.port_b_logical_ram_width = 32;
defparam ram_block3a62.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_read_enable_clock = "clock1";
defparam ram_block3a62.port_b_write_enable_clock = "clock1";
defparam ram_block3a62.ram_block_type = "M9K";
defparam ram_block3a62.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y35_N0
cycloneive_ram_block ram_block3a30(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a30_PORTADATAOUT_bus),
	.portbdataout(ram_block3a30_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a30.clk0_core_clock_enable = "ena0";
defparam ram_block3a30.clk1_core_clock_enable = "ena1";
defparam ram_block3a30.data_interleave_offset_in_bits = 1;
defparam ram_block3a30.data_interleave_width_in_bits = 1;
defparam ram_block3a30.init_file = "meminit.hex";
defparam ram_block3a30.init_file_layout = "port_a";
defparam ram_block3a30.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a30.operation_mode = "bidir_dual_port";
defparam ram_block3a30.port_a_address_clear = "none";
defparam ram_block3a30.port_a_address_width = 13;
defparam ram_block3a30.port_a_byte_enable_clock = "none";
defparam ram_block3a30.port_a_data_out_clear = "none";
defparam ram_block3a30.port_a_data_out_clock = "none";
defparam ram_block3a30.port_a_data_width = 1;
defparam ram_block3a30.port_a_first_address = 0;
defparam ram_block3a30.port_a_first_bit_number = 30;
defparam ram_block3a30.port_a_last_address = 8191;
defparam ram_block3a30.port_a_logical_ram_depth = 16384;
defparam ram_block3a30.port_a_logical_ram_width = 32;
defparam ram_block3a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_address_clear = "none";
defparam ram_block3a30.port_b_address_clock = "clock1";
defparam ram_block3a30.port_b_address_width = 13;
defparam ram_block3a30.port_b_data_in_clock = "clock1";
defparam ram_block3a30.port_b_data_out_clear = "none";
defparam ram_block3a30.port_b_data_out_clock = "none";
defparam ram_block3a30.port_b_data_width = 1;
defparam ram_block3a30.port_b_first_address = 0;
defparam ram_block3a30.port_b_first_bit_number = 30;
defparam ram_block3a30.port_b_last_address = 8191;
defparam ram_block3a30.port_b_logical_ram_depth = 16384;
defparam ram_block3a30.port_b_logical_ram_width = 32;
defparam ram_block3a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_read_enable_clock = "clock1";
defparam ram_block3a30.port_b_write_enable_clock = "clock1";
defparam ram_block3a30.ram_block_type = "M9K";
defparam ram_block3a30.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004000000;
// synopsys translate_on

// Location: M9K_X64_Y31_N0
cycloneive_ram_block ram_block3a63(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a63_PORTADATAOUT_bus),
	.portbdataout(ram_block3a63_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a63.clk0_core_clock_enable = "ena0";
defparam ram_block3a63.clk1_core_clock_enable = "ena1";
defparam ram_block3a63.data_interleave_offset_in_bits = 1;
defparam ram_block3a63.data_interleave_width_in_bits = 1;
defparam ram_block3a63.init_file = "meminit.hex";
defparam ram_block3a63.init_file_layout = "port_a";
defparam ram_block3a63.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a63.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a63.operation_mode = "bidir_dual_port";
defparam ram_block3a63.port_a_address_clear = "none";
defparam ram_block3a63.port_a_address_width = 13;
defparam ram_block3a63.port_a_byte_enable_clock = "none";
defparam ram_block3a63.port_a_data_out_clear = "none";
defparam ram_block3a63.port_a_data_out_clock = "none";
defparam ram_block3a63.port_a_data_width = 1;
defparam ram_block3a63.port_a_first_address = 0;
defparam ram_block3a63.port_a_first_bit_number = 31;
defparam ram_block3a63.port_a_last_address = 8191;
defparam ram_block3a63.port_a_logical_ram_depth = 16384;
defparam ram_block3a63.port_a_logical_ram_width = 32;
defparam ram_block3a63.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_address_clear = "none";
defparam ram_block3a63.port_b_address_clock = "clock1";
defparam ram_block3a63.port_b_address_width = 13;
defparam ram_block3a63.port_b_data_in_clock = "clock1";
defparam ram_block3a63.port_b_data_out_clear = "none";
defparam ram_block3a63.port_b_data_out_clock = "none";
defparam ram_block3a63.port_b_data_width = 1;
defparam ram_block3a63.port_b_first_address = 0;
defparam ram_block3a63.port_b_first_bit_number = 31;
defparam ram_block3a63.port_b_last_address = 8191;
defparam ram_block3a63.port_b_logical_ram_depth = 16384;
defparam ram_block3a63.port_b_logical_ram_width = 32;
defparam ram_block3a63.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_read_enable_clock = "clock1";
defparam ram_block3a63.port_b_write_enable_clock = "clock1";
defparam ram_block3a63.ram_block_type = "M9K";
defparam ram_block3a63.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y34_N0
cycloneive_ram_block ram_block3a31(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a31_PORTADATAOUT_bus),
	.portbdataout(ram_block3a31_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a31.clk0_core_clock_enable = "ena0";
defparam ram_block3a31.clk1_core_clock_enable = "ena1";
defparam ram_block3a31.data_interleave_offset_in_bits = 1;
defparam ram_block3a31.data_interleave_width_in_bits = 1;
defparam ram_block3a31.init_file = "meminit.hex";
defparam ram_block3a31.init_file_layout = "port_a";
defparam ram_block3a31.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a31.operation_mode = "bidir_dual_port";
defparam ram_block3a31.port_a_address_clear = "none";
defparam ram_block3a31.port_a_address_width = 13;
defparam ram_block3a31.port_a_byte_enable_clock = "none";
defparam ram_block3a31.port_a_data_out_clear = "none";
defparam ram_block3a31.port_a_data_out_clock = "none";
defparam ram_block3a31.port_a_data_width = 1;
defparam ram_block3a31.port_a_first_address = 0;
defparam ram_block3a31.port_a_first_bit_number = 31;
defparam ram_block3a31.port_a_last_address = 8191;
defparam ram_block3a31.port_a_logical_ram_depth = 16384;
defparam ram_block3a31.port_a_logical_ram_width = 32;
defparam ram_block3a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_address_clear = "none";
defparam ram_block3a31.port_b_address_clock = "clock1";
defparam ram_block3a31.port_b_address_width = 13;
defparam ram_block3a31.port_b_data_in_clock = "clock1";
defparam ram_block3a31.port_b_data_out_clear = "none";
defparam ram_block3a31.port_b_data_out_clock = "none";
defparam ram_block3a31.port_b_data_width = 1;
defparam ram_block3a31.port_b_first_address = 0;
defparam ram_block3a31.port_b_first_bit_number = 31;
defparam ram_block3a31.port_b_last_address = 8191;
defparam ram_block3a31.port_b_logical_ram_depth = 16384;
defparam ram_block3a31.port_b_logical_ram_width = 32;
defparam ram_block3a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_read_enable_clock = "clock1";
defparam ram_block3a31.port_b_write_enable_clock = "clock1";
defparam ram_block3a31.ram_block_type = "M9K";
defparam ram_block3a31.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FF8000;
// synopsys translate_on

// Location: FF_X57_Y35_N1
dffeas \address_reg_a[0] (
	.clk(clock0),
	.d(gnd),
	.asdata(ramaddr1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_a_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_a[0] .is_wysiwyg = "true";
defparam \address_reg_a[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N17
dffeas \address_reg_b[0] (
	.clk(clock1),
	.d(\address_reg_b[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_b_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_b[0] .is_wysiwyg = "true";
defparam \address_reg_b[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N16
cycloneive_lcell_comb \address_reg_b[0]~feeder (
// Equation(s):
// \address_reg_b[0]~feeder_combout  = ram_rom_addr_reg_13

	.dataa(gnd),
	.datab(gnd),
	.datac(ram_rom_addr_reg_13),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_reg_b[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \address_reg_b[0]~feeder .lut_mask = 16'hF0F0;
defparam \address_reg_b[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa (
	ramaddr,
	ramWEN,
	always1,
	eq_node_1,
	eq_node_0,
	devpor,
	devclrn,
	devoe);
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	eq_node_1;
output 	eq_node_0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X62_Y32_N8
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (always1 & (!\ramWEN~0_combout  & !\ramaddr~29_combout ))

	.dataa(always1),
	.datab(ramWEN),
	.datac(gnd),
	.datad(ramaddr),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h0022;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N22
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (always1 & (!\ramWEN~0_combout  & \ramaddr~29_combout ))

	.dataa(always1),
	.datab(ramWEN),
	.datac(gnd),
	.datad(ramaddr),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h2200;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa_1 (
	ram_rom_addr_reg_13,
	sdr,
	eq_node_1,
	eq_node_0,
	irf_reg_2_1,
	state_5,
	devpor,
	devclrn,
	devoe);
input 	ram_rom_addr_reg_13;
input 	sdr;
output 	eq_node_1;
output 	eq_node_0;
input 	irf_reg_2_1;
input 	state_5;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X41_Y30_N2
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5] & (ram_rom_addr_reg_13 & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q  & sdr)))

	.dataa(state_5),
	.datab(ram_rom_addr_reg_13),
	.datac(irf_reg_2_1),
	.datad(sdr),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h8000;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y30_N12
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5] & (!ram_rom_addr_reg_13 & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q  & sdr)))

	.dataa(state_5),
	.datab(ram_rom_addr_reg_13),
	.datac(irf_reg_2_1),
	.datad(sdr),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h2000;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_mod_ram_rom (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg1,
	ram_rom_data_reg_0,
	ram_rom_addr_reg_13,
	ram_rom_addr_reg_0,
	ram_rom_addr_reg_1,
	ram_rom_addr_reg_2,
	ram_rom_addr_reg_3,
	ram_rom_addr_reg_4,
	ram_rom_addr_reg_5,
	ram_rom_addr_reg_6,
	ram_rom_addr_reg_7,
	ram_rom_addr_reg_8,
	ram_rom_addr_reg_9,
	ram_rom_addr_reg_10,
	ram_rom_addr_reg_11,
	ram_rom_addr_reg_12,
	ram_rom_data_reg_1,
	ram_rom_data_reg_2,
	ram_rom_data_reg_3,
	ram_rom_data_reg_4,
	ram_rom_data_reg_5,
	ram_rom_data_reg_6,
	ram_rom_data_reg_7,
	ram_rom_data_reg_8,
	ram_rom_data_reg_9,
	ram_rom_data_reg_10,
	ram_rom_data_reg_11,
	ram_rom_data_reg_12,
	ram_rom_data_reg_13,
	ram_rom_data_reg_14,
	ram_rom_data_reg_15,
	ram_rom_data_reg_16,
	ram_rom_data_reg_17,
	ram_rom_data_reg_18,
	ram_rom_data_reg_19,
	ram_rom_data_reg_20,
	ram_rom_data_reg_21,
	ram_rom_data_reg_22,
	ram_rom_data_reg_23,
	ram_rom_data_reg_24,
	ram_rom_data_reg_25,
	ram_rom_data_reg_26,
	ram_rom_data_reg_27,
	ram_rom_data_reg_28,
	ram_rom_data_reg_29,
	ram_rom_data_reg_30,
	ram_rom_data_reg_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	sdr,
	address_reg_b_0,
	altera_internal_jtag,
	state_4,
	ir_in,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_4_1,
	node_ena_1,
	clr,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	raw_tck,
	devpor,
	devclrn,
	devoe);
input 	ram_block3a32;
input 	ram_block3a0;
input 	ram_block3a33;
input 	ram_block3a1;
input 	ram_block3a34;
input 	ram_block3a2;
input 	ram_block3a35;
input 	ram_block3a3;
input 	ram_block3a36;
input 	ram_block3a4;
input 	ram_block3a37;
input 	ram_block3a5;
input 	ram_block3a38;
input 	ram_block3a6;
input 	ram_block3a39;
input 	ram_block3a7;
input 	ram_block3a40;
input 	ram_block3a8;
input 	ram_block3a41;
input 	ram_block3a9;
input 	ram_block3a42;
input 	ram_block3a10;
input 	ram_block3a43;
input 	ram_block3a11;
input 	ram_block3a44;
input 	ram_block3a12;
input 	ram_block3a45;
input 	ram_block3a13;
input 	ram_block3a46;
input 	ram_block3a14;
input 	ram_block3a47;
input 	ram_block3a15;
input 	ram_block3a48;
input 	ram_block3a16;
input 	ram_block3a49;
input 	ram_block3a17;
input 	ram_block3a50;
input 	ram_block3a18;
input 	ram_block3a51;
input 	ram_block3a19;
input 	ram_block3a52;
input 	ram_block3a20;
input 	ram_block3a53;
input 	ram_block3a21;
input 	ram_block3a54;
input 	ram_block3a22;
input 	ram_block3a55;
input 	ram_block3a23;
input 	ram_block3a56;
input 	ram_block3a24;
input 	ram_block3a57;
input 	ram_block3a25;
input 	ram_block3a58;
input 	ram_block3a26;
input 	ram_block3a59;
input 	ram_block3a27;
input 	ram_block3a60;
input 	ram_block3a28;
input 	ram_block3a61;
input 	ram_block3a29;
input 	ram_block3a62;
input 	ram_block3a30;
input 	ram_block3a63;
input 	ram_block3a31;
output 	is_in_use_reg1;
output 	ram_rom_data_reg_0;
output 	ram_rom_addr_reg_13;
output 	ram_rom_addr_reg_0;
output 	ram_rom_addr_reg_1;
output 	ram_rom_addr_reg_2;
output 	ram_rom_addr_reg_3;
output 	ram_rom_addr_reg_4;
output 	ram_rom_addr_reg_5;
output 	ram_rom_addr_reg_6;
output 	ram_rom_addr_reg_7;
output 	ram_rom_addr_reg_8;
output 	ram_rom_addr_reg_9;
output 	ram_rom_addr_reg_10;
output 	ram_rom_addr_reg_11;
output 	ram_rom_addr_reg_12;
output 	ram_rom_data_reg_1;
output 	ram_rom_data_reg_2;
output 	ram_rom_data_reg_3;
output 	ram_rom_data_reg_4;
output 	ram_rom_data_reg_5;
output 	ram_rom_data_reg_6;
output 	ram_rom_data_reg_7;
output 	ram_rom_data_reg_8;
output 	ram_rom_data_reg_9;
output 	ram_rom_data_reg_10;
output 	ram_rom_data_reg_11;
output 	ram_rom_data_reg_12;
output 	ram_rom_data_reg_13;
output 	ram_rom_data_reg_14;
output 	ram_rom_data_reg_15;
output 	ram_rom_data_reg_16;
output 	ram_rom_data_reg_17;
output 	ram_rom_data_reg_18;
output 	ram_rom_data_reg_19;
output 	ram_rom_data_reg_20;
output 	ram_rom_data_reg_21;
output 	ram_rom_data_reg_22;
output 	ram_rom_data_reg_23;
output 	ram_rom_data_reg_24;
output 	ram_rom_data_reg_25;
output 	ram_rom_data_reg_26;
output 	ram_rom_data_reg_27;
output 	ram_rom_data_reg_28;
output 	ram_rom_data_reg_29;
output 	ram_rom_data_reg_30;
output 	ram_rom_data_reg_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
output 	sdr;
input 	address_reg_b_0;
input 	altera_internal_jtag;
input 	state_4;
input 	[4:0] ir_in;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	raw_tck;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~0_combout ;
wire \Add1~4_combout ;
wire \Add1~9 ;
wire \Add1~10_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~10_combout ;
wire \is_in_use_reg~0_combout ;
wire \ram_rom_data_reg[0]~0_combout ;
wire \Add1~1 ;
wire \Add1~2_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~4_combout ;
wire \ram_rom_data_shift_cntr_reg[1]~5_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~11_combout ;
wire \ram_rom_data_shift_cntr_reg[0]~6_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~12_combout ;
wire \ram_rom_data_shift_cntr_reg[2]~9_combout ;
wire \Add1~3 ;
wire \Add1~5 ;
wire \Add1~7 ;
wire \Add1~8_combout ;
wire \ram_rom_data_shift_cntr_reg[4]~7_combout ;
wire \Add1~6_combout ;
wire \ram_rom_data_shift_cntr_reg[3]~8_combout ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \process_0~2_combout ;
wire \ram_rom_data_reg[12]~32_combout ;
wire \ram_rom_addr_reg[0]~15 ;
wire \ram_rom_addr_reg[1]~17 ;
wire \ram_rom_addr_reg[2]~19 ;
wire \ram_rom_addr_reg[3]~21 ;
wire \ram_rom_addr_reg[4]~23 ;
wire \ram_rom_addr_reg[5]~25 ;
wire \ram_rom_addr_reg[6]~27 ;
wire \ram_rom_addr_reg[7]~29 ;
wire \ram_rom_addr_reg[8]~31 ;
wire \ram_rom_addr_reg[9]~33 ;
wire \ram_rom_addr_reg[10]~35 ;
wire \ram_rom_addr_reg[11]~37 ;
wire \ram_rom_addr_reg[12]~39 ;
wire \ram_rom_addr_reg[13]~40_combout ;
wire \process_0~3_combout ;
wire \ram_rom_addr_reg[1]~42_combout ;
wire \ram_rom_addr_reg[1]~43_combout ;
wire \ram_rom_addr_reg[0]~14_combout ;
wire \ram_rom_addr_reg[1]~16_combout ;
wire \ram_rom_addr_reg[2]~18_combout ;
wire \ram_rom_addr_reg[3]~20_combout ;
wire \ram_rom_addr_reg[4]~22_combout ;
wire \ram_rom_addr_reg[5]~24_combout ;
wire \ram_rom_addr_reg[6]~26_combout ;
wire \ram_rom_addr_reg[7]~28_combout ;
wire \ram_rom_addr_reg[8]~30_combout ;
wire \ram_rom_addr_reg[9]~32_combout ;
wire \ram_rom_addr_reg[10]~34_combout ;
wire \ram_rom_addr_reg[11]~36_combout ;
wire \ram_rom_addr_reg[12]~38_combout ;
wire \ram_rom_data_reg[1]~1_combout ;
wire \ram_rom_data_reg[2]~2_combout ;
wire \ram_rom_data_reg[3]~3_combout ;
wire \ram_rom_data_reg[4]~4_combout ;
wire \ram_rom_data_reg[5]~5_combout ;
wire \ram_rom_data_reg[6]~6_combout ;
wire \ram_rom_data_reg[7]~7_combout ;
wire \ram_rom_data_reg[8]~8_combout ;
wire \ram_rom_data_reg[9]~9_combout ;
wire \ram_rom_data_reg[10]~10_combout ;
wire \ram_rom_data_reg[11]~11_combout ;
wire \ram_rom_data_reg[12]~12_combout ;
wire \ram_rom_data_reg[13]~13_combout ;
wire \ram_rom_data_reg[14]~14_combout ;
wire \ram_rom_data_reg[15]~15_combout ;
wire \ram_rom_data_reg[16]~16_combout ;
wire \ram_rom_data_reg[17]~17_combout ;
wire \ram_rom_data_reg[18]~18_combout ;
wire \ram_rom_data_reg[19]~19_combout ;
wire \ram_rom_data_reg[20]~20_combout ;
wire \ram_rom_data_reg[21]~21_combout ;
wire \ram_rom_data_reg[22]~22_combout ;
wire \ram_rom_data_reg[23]~23_combout ;
wire \ram_rom_data_reg[24]~24_combout ;
wire \ram_rom_data_reg[25]~25_combout ;
wire \ram_rom_data_reg[26]~26_combout ;
wire \ram_rom_data_reg[27]~27_combout ;
wire \ram_rom_data_reg[28]~28_combout ;
wire \ram_rom_data_reg[29]~29_combout ;
wire \ram_rom_data_reg[30]~30_combout ;
wire \ram_rom_data_reg[31]~31_combout ;
wire \ir_loaded_address_reg[0]~feeder_combout ;
wire \process_0~0_combout ;
wire \process_0~1_combout ;
wire \ir_loaded_address_reg[1]~feeder_combout ;
wire \ir_loaded_address_reg[3]~feeder_combout ;
wire \bypass_reg_out~0_combout ;
wire \bypass_reg_out~q ;
wire \tdo~0_combout ;
wire [5:0] ram_rom_data_shift_cntr_reg;
wire [3:0] \ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR ;


sld_rom_sr \ram_rom_logic_gen:name_gen:info_rom_sr (
	.WORD_SR_0(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.sdr(sdr),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.TCK(raw_tck),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X42_Y30_N12
cycloneive_lcell_comb \Add1~0 (
	.dataa(ram_rom_data_shift_cntr_reg[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h55AA;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y30_N16
cycloneive_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'hC30C;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X42_Y30_N20
cycloneive_lcell_comb \Add1~8 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'hC30C;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X42_Y30_N22
cycloneive_lcell_comb \Add1~10 (
	.dataa(ram_rom_data_shift_cntr_reg[5]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h5A5A;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X42_Y30_N27
dffeas \ram_rom_data_shift_cntr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[5]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y30_N26
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~10 (
	.dataa(\Add1~10_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[5]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~10 .lut_mask = 16'hC0EA;
defparam \ram_rom_data_shift_cntr_reg[5]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y30_N29
dffeas is_in_use_reg(
	.clk(raw_tck),
	.d(\is_in_use_reg~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(ir_in[0]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(is_in_use_reg1),
	.prn(vcc));
// synopsys translate_off
defparam is_in_use_reg.is_wysiwyg = "true";
defparam is_in_use_reg.power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N1
dffeas \ram_rom_data_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[0]~0_combout ),
	.asdata(ram_rom_data_reg_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y29_N29
dffeas \ram_rom_addr_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[13]~40_combout ),
	.asdata(altera_internal_jtag),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[1]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y29_N3
dffeas \ram_rom_addr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[0]~14_combout ),
	.asdata(ram_rom_addr_reg_1),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[1]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y29_N5
dffeas \ram_rom_addr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[1]~16_combout ),
	.asdata(ram_rom_addr_reg_2),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[1]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y29_N7
dffeas \ram_rom_addr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[2]~18_combout ),
	.asdata(ram_rom_addr_reg_3),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[1]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y29_N9
dffeas \ram_rom_addr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[3]~20_combout ),
	.asdata(ram_rom_addr_reg_4),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[1]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y29_N11
dffeas \ram_rom_addr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[4]~22_combout ),
	.asdata(ram_rom_addr_reg_5),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[1]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y29_N13
dffeas \ram_rom_addr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[5]~24_combout ),
	.asdata(ram_rom_addr_reg_6),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[1]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y29_N15
dffeas \ram_rom_addr_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[6]~26_combout ),
	.asdata(ram_rom_addr_reg_7),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[1]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y29_N17
dffeas \ram_rom_addr_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[7]~28_combout ),
	.asdata(ram_rom_addr_reg_8),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[1]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y29_N19
dffeas \ram_rom_addr_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[8]~30_combout ),
	.asdata(ram_rom_addr_reg_9),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[1]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y29_N21
dffeas \ram_rom_addr_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[9]~32_combout ),
	.asdata(ram_rom_addr_reg_10),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[1]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y29_N23
dffeas \ram_rom_addr_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[10]~34_combout ),
	.asdata(ram_rom_addr_reg_11),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[1]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y29_N25
dffeas \ram_rom_addr_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[11]~36_combout ),
	.asdata(ram_rom_addr_reg_12),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[1]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X40_Y29_N27
dffeas \ram_rom_addr_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[12]~38_combout ),
	.asdata(ram_rom_addr_reg_13),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[1]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N15
dffeas \ram_rom_data_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[1]~1_combout ),
	.asdata(ram_rom_data_reg_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N29
dffeas \ram_rom_data_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[2]~2_combout ),
	.asdata(ram_rom_data_reg_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N27
dffeas \ram_rom_data_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[3]~3_combout ),
	.asdata(ram_rom_data_reg_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N13
dffeas \ram_rom_data_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[4]~4_combout ),
	.asdata(ram_rom_data_reg_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N23
dffeas \ram_rom_data_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[5]~5_combout ),
	.asdata(ram_rom_data_reg_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N9
dffeas \ram_rom_data_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[6]~6_combout ),
	.asdata(ram_rom_data_reg_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N19
dffeas \ram_rom_data_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[7]~7_combout ),
	.asdata(ram_rom_data_reg_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N29
dffeas \ram_rom_data_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[8]~8_combout ),
	.asdata(ram_rom_data_reg_9),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N17
dffeas \ram_rom_data_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[9]~9_combout ),
	.asdata(ram_rom_data_reg_10),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N25
dffeas \ram_rom_data_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[10]~10_combout ),
	.asdata(ram_rom_data_reg_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N31
dffeas \ram_rom_data_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[11]~11_combout ),
	.asdata(ram_rom_data_reg_12),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N13
dffeas \ram_rom_data_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[12]~12_combout ),
	.asdata(ram_rom_data_reg_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N27
dffeas \ram_rom_data_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[13]~13_combout ),
	.asdata(ram_rom_data_reg_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N25
dffeas \ram_rom_data_reg[14] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[14]~14_combout ),
	.asdata(ram_rom_data_reg_15),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_14),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[14] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N21
dffeas \ram_rom_data_reg[15] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[15]~15_combout ),
	.asdata(ram_rom_data_reg_16),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_15),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[15] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N23
dffeas \ram_rom_data_reg[16] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[16]~16_combout ),
	.asdata(ram_rom_data_reg_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_16),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[16] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N1
dffeas \ram_rom_data_reg[17] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[17]~17_combout ),
	.asdata(ram_rom_data_reg_18),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_17),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[17] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N19
dffeas \ram_rom_data_reg[18] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[18]~18_combout ),
	.asdata(ram_rom_data_reg_19),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_18),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[18] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y33_N9
dffeas \ram_rom_data_reg[19] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[19]~19_combout ),
	.asdata(ram_rom_data_reg_20),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_19),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[19] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N1
dffeas \ram_rom_data_reg[20] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[20]~20_combout ),
	.asdata(ram_rom_data_reg_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_20),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[20] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N31
dffeas \ram_rom_data_reg[21] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[21]~21_combout ),
	.asdata(ram_rom_data_reg_22),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_21),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[21] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N31
dffeas \ram_rom_data_reg[22] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[22]~22_combout ),
	.asdata(ram_rom_data_reg_23),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_22),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[22] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N25
dffeas \ram_rom_data_reg[23] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[23]~23_combout ),
	.asdata(ram_rom_data_reg_24),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_23),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[23] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N15
dffeas \ram_rom_data_reg[24] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[24]~24_combout ),
	.asdata(ram_rom_data_reg_25),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_24),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[24] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N9
dffeas \ram_rom_data_reg[25] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[25]~25_combout ),
	.asdata(ram_rom_data_reg_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_25),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[25] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N23
dffeas \ram_rom_data_reg[26] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[26]~26_combout ),
	.asdata(ram_rom_data_reg_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_26),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[26] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N13
dffeas \ram_rom_data_reg[27] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[27]~27_combout ),
	.asdata(ram_rom_data_reg_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_27),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[27] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N27
dffeas \ram_rom_data_reg[28] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[28]~28_combout ),
	.asdata(ram_rom_data_reg_29),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_28),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[28] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N17
dffeas \ram_rom_data_reg[29] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[29]~29_combout ),
	.asdata(ram_rom_data_reg_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_29),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[29] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N19
dffeas \ram_rom_data_reg[30] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[30]~30_combout ),
	.asdata(ram_rom_data_reg_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_30),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[30] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N5
dffeas \ram_rom_data_reg[31] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[31]~31_combout ),
	.asdata(altera_internal_jtag),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[12]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_31),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[31] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y30_N9
dffeas \ir_loaded_address_reg[0] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[0] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y30_N15
dffeas \ir_loaded_address_reg[1] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[1] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y30_N1
dffeas \ir_loaded_address_reg[2] (
	.clk(raw_tck),
	.d(gnd),
	.asdata(ram_rom_addr_reg_2),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[2] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X41_Y30_N23
dffeas \ir_loaded_address_reg[3] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[3] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X40_Y30_N12
cycloneive_lcell_comb \tdo~1 (
	.dataa(ir_in[0]),
	.datab(gnd),
	.datac(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.datad(\tdo~0_combout ),
	.cin(gnd),
	.combout(tdo),
	.cout());
// synopsys translate_off
defparam \tdo~1 .lut_mask = 16'hF5A0;
defparam \tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y30_N4
cycloneive_lcell_comb \sdr~0 (
	.dataa(node_ena_1),
	.datab(gnd),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(sdr),
	.cout());
// synopsys translate_off
defparam \sdr~0 .lut_mask = 16'h00AA;
defparam \sdr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y30_N28
cycloneive_lcell_comb \is_in_use_reg~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(is_in_use_reg1),
	.datad(irf_reg_4_1),
	.cin(gnd),
	.combout(\is_in_use_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \is_in_use_reg~0 .lut_mask = 16'h00F0;
defparam \is_in_use_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N0
cycloneive_lcell_comb \ram_rom_data_reg[0]~0 (
	.dataa(ram_block3a0),
	.datab(ram_block3a32),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[0]~0 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y30_N14
cycloneive_lcell_comb \Add1~2 (
	.dataa(ram_rom_data_shift_cntr_reg[1]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h5A5F;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X41_Y30_N20
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~4 (
	.dataa(irf_reg_1_1),
	.datab(state_4),
	.datac(irf_reg_2_1),
	.datad(sdr),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~4 .lut_mask = 16'hC800;
defparam \ram_rom_data_shift_cntr_reg[5]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y30_N0
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[1]~5 (
	.dataa(\Equal1~1_combout ),
	.datab(\Add1~2_combout ),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1]~5 .lut_mask = 16'h4C50;
defparam \ram_rom_data_shift_cntr_reg[1]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y30_N1
dffeas \ram_rom_data_shift_cntr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[1]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y30_N28
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~11 (
	.dataa(ram_rom_data_shift_cntr_reg[1]),
	.datab(\Equal1~0_combout ),
	.datac(ram_rom_data_shift_cntr_reg[0]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~11 .lut_mask = 16'h007F;
defparam \ram_rom_data_shift_cntr_reg[5]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y30_N30
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[0]~6 (
	.dataa(\Add1~0_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[0]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0]~6 .lut_mask = 16'hC0EA;
defparam \ram_rom_data_shift_cntr_reg[0]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y30_N31
dffeas \ram_rom_data_shift_cntr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[0]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y30_N2
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~12 (
	.dataa(ram_rom_data_shift_cntr_reg[1]),
	.datab(\Equal1~0_combout ),
	.datac(ram_rom_data_shift_cntr_reg[0]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~12 .lut_mask = 16'h80FF;
defparam \ram_rom_data_shift_cntr_reg[5]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y30_N8
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[2]~9 (
	.dataa(\Add1~4_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.datac(ram_rom_data_shift_cntr_reg[2]),
	.datad(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2]~9 .lut_mask = 16'hC0EA;
defparam \ram_rom_data_shift_cntr_reg[2]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y30_N9
dffeas \ram_rom_data_shift_cntr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[2]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y30_N18
cycloneive_lcell_comb \Add1~6 (
	.dataa(ram_rom_data_shift_cntr_reg[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h5A5F;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X42_Y30_N24
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[4]~7 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datac(ram_rom_data_shift_cntr_reg[4]),
	.datad(\Add1~8_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4]~7 .lut_mask = 16'hB3A0;
defparam \ram_rom_data_shift_cntr_reg[4]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y30_N25
dffeas \ram_rom_data_shift_cntr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[4]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y30_N10
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[3]~8 (
	.dataa(\ram_rom_data_shift_cntr_reg[5]~11_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datac(ram_rom_data_shift_cntr_reg[3]),
	.datad(\Add1~6_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3]~8 .lut_mask = 16'hB3A0;
defparam \ram_rom_data_shift_cntr_reg[3]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y30_N11
dffeas \ram_rom_data_shift_cntr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[3]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y30_N4
cycloneive_lcell_comb \Equal1~0 (
	.dataa(ram_rom_data_shift_cntr_reg[5]),
	.datab(ram_rom_data_shift_cntr_reg[4]),
	.datac(ram_rom_data_shift_cntr_reg[2]),
	.datad(ram_rom_data_shift_cntr_reg[3]),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~0 .lut_mask = 16'h4000;
defparam \Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y30_N6
cycloneive_lcell_comb \Equal1~1 (
	.dataa(gnd),
	.datab(\Equal1~0_combout ),
	.datac(ram_rom_data_shift_cntr_reg[0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~1 .lut_mask = 16'hC0C0;
defparam \Equal1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y30_N14
cycloneive_lcell_comb \process_0~2 (
	.dataa(irf_reg_1_1),
	.datab(ir_in[3]),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\process_0~2_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~2 .lut_mask = 16'h1333;
defparam \process_0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N10
cycloneive_lcell_comb \ram_rom_data_reg[12]~32 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datad(\process_0~2_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_reg[12]~32_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[12]~32 .lut_mask = 16'hF0FF;
defparam \ram_rom_data_reg[12]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y29_N2
cycloneive_lcell_comb \ram_rom_addr_reg[0]~14 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[0]~14_combout ),
	.cout(\ram_rom_addr_reg[0]~15 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[0]~14 .lut_mask = 16'h33CC;
defparam \ram_rom_addr_reg[0]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X40_Y29_N4
cycloneive_lcell_comb \ram_rom_addr_reg[1]~16 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[0]~15 ),
	.combout(\ram_rom_addr_reg[1]~16_combout ),
	.cout(\ram_rom_addr_reg[1]~17 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[1]~16 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[1]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X40_Y29_N6
cycloneive_lcell_comb \ram_rom_addr_reg[2]~18 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[1]~17 ),
	.combout(\ram_rom_addr_reg[2]~18_combout ),
	.cout(\ram_rom_addr_reg[2]~19 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[2]~18 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[2]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X40_Y29_N8
cycloneive_lcell_comb \ram_rom_addr_reg[3]~20 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[2]~19 ),
	.combout(\ram_rom_addr_reg[3]~20_combout ),
	.cout(\ram_rom_addr_reg[3]~21 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[3]~20 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[3]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X40_Y29_N10
cycloneive_lcell_comb \ram_rom_addr_reg[4]~22 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[3]~21 ),
	.combout(\ram_rom_addr_reg[4]~22_combout ),
	.cout(\ram_rom_addr_reg[4]~23 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[4]~22 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[4]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X40_Y29_N12
cycloneive_lcell_comb \ram_rom_addr_reg[5]~24 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[4]~23 ),
	.combout(\ram_rom_addr_reg[5]~24_combout ),
	.cout(\ram_rom_addr_reg[5]~25 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[5]~24 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[5]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X40_Y29_N14
cycloneive_lcell_comb \ram_rom_addr_reg[6]~26 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[5]~25 ),
	.combout(\ram_rom_addr_reg[6]~26_combout ),
	.cout(\ram_rom_addr_reg[6]~27 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[6]~26 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[6]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X40_Y29_N16
cycloneive_lcell_comb \ram_rom_addr_reg[7]~28 (
	.dataa(ram_rom_addr_reg_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[6]~27 ),
	.combout(\ram_rom_addr_reg[7]~28_combout ),
	.cout(\ram_rom_addr_reg[7]~29 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[7]~28 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[7]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X40_Y29_N18
cycloneive_lcell_comb \ram_rom_addr_reg[8]~30 (
	.dataa(ram_rom_addr_reg_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[7]~29 ),
	.combout(\ram_rom_addr_reg[8]~30_combout ),
	.cout(\ram_rom_addr_reg[8]~31 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[8]~30 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[8]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X40_Y29_N20
cycloneive_lcell_comb \ram_rom_addr_reg[9]~32 (
	.dataa(ram_rom_addr_reg_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[8]~31 ),
	.combout(\ram_rom_addr_reg[9]~32_combout ),
	.cout(\ram_rom_addr_reg[9]~33 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[9]~32 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[9]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X40_Y29_N22
cycloneive_lcell_comb \ram_rom_addr_reg[10]~34 (
	.dataa(ram_rom_addr_reg_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[9]~33 ),
	.combout(\ram_rom_addr_reg[10]~34_combout ),
	.cout(\ram_rom_addr_reg[10]~35 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[10]~34 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[10]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X40_Y29_N24
cycloneive_lcell_comb \ram_rom_addr_reg[11]~36 (
	.dataa(ram_rom_addr_reg_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[10]~35 ),
	.combout(\ram_rom_addr_reg[11]~36_combout ),
	.cout(\ram_rom_addr_reg[11]~37 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[11]~36 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[11]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X40_Y29_N26
cycloneive_lcell_comb \ram_rom_addr_reg[12]~38 (
	.dataa(ram_rom_addr_reg_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[11]~37 ),
	.combout(\ram_rom_addr_reg[12]~38_combout ),
	.cout(\ram_rom_addr_reg[12]~39 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[12]~38 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[12]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X40_Y29_N28
cycloneive_lcell_comb \ram_rom_addr_reg[13]~40 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_13),
	.datac(gnd),
	.datad(gnd),
	.cin(\ram_rom_addr_reg[12]~39 ),
	.combout(\ram_rom_addr_reg[13]~40_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[13]~40 .lut_mask = 16'h3C3C;
defparam \ram_rom_addr_reg[13]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X41_Y30_N30
cycloneive_lcell_comb \process_0~3 (
	.dataa(node_ena_1),
	.datab(virtual_ir_scan_reg),
	.datac(state_4),
	.datad(ir_in[3]),
	.cin(gnd),
	.combout(\process_0~3_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~3 .lut_mask = 16'h2000;
defparam \process_0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y30_N0
cycloneive_lcell_comb \ram_rom_addr_reg[1]~42 (
	.dataa(irf_reg_1_1),
	.datab(ram_rom_data_shift_cntr_reg[1]),
	.datac(\process_0~3_combout ),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[1]~42_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[1]~42 .lut_mask = 16'hF2F0;
defparam \ram_rom_addr_reg[1]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y30_N18
cycloneive_lcell_comb \ram_rom_addr_reg[1]~43 (
	.dataa(irf_reg_2_1),
	.datab(\ram_rom_addr_reg[1]~42_combout ),
	.datac(state_8),
	.datad(sdr),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[1]~43_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[1]~43 .lut_mask = 16'hECCC;
defparam \ram_rom_addr_reg[1]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N14
cycloneive_lcell_comb \ram_rom_data_reg[1]~1 (
	.dataa(ram_block3a33),
	.datab(ram_block3a1),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[1]~1 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N28
cycloneive_lcell_comb \ram_rom_data_reg[2]~2 (
	.dataa(ram_block3a34),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a2),
	.cin(gnd),
	.combout(\ram_rom_data_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[2]~2 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N26
cycloneive_lcell_comb \ram_rom_data_reg[3]~3 (
	.dataa(ram_block3a35),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a3),
	.cin(gnd),
	.combout(\ram_rom_data_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[3]~3 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N12
cycloneive_lcell_comb \ram_rom_data_reg[4]~4 (
	.dataa(ram_block3a36),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a4),
	.cin(gnd),
	.combout(\ram_rom_data_reg[4]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[4]~4 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N22
cycloneive_lcell_comb \ram_rom_data_reg[5]~5 (
	.dataa(ram_block3a37),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a5),
	.cin(gnd),
	.combout(\ram_rom_data_reg[5]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[5]~5 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[5]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N8
cycloneive_lcell_comb \ram_rom_data_reg[6]~6 (
	.dataa(ram_block3a6),
	.datab(ram_block3a38),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[6]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[6]~6 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[6]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N18
cycloneive_lcell_comb \ram_rom_data_reg[7]~7 (
	.dataa(ram_block3a7),
	.datab(ram_block3a39),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[7]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[7]~7 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[7]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N28
cycloneive_lcell_comb \ram_rom_data_reg[8]~8 (
	.dataa(ram_block3a8),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a40),
	.cin(gnd),
	.combout(\ram_rom_data_reg[8]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[8]~8 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[8]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N16
cycloneive_lcell_comb \ram_rom_data_reg[9]~9 (
	.dataa(ram_block3a9),
	.datab(ram_block3a41),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[9]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[9]~9 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[9]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N24
cycloneive_lcell_comb \ram_rom_data_reg[10]~10 (
	.dataa(ram_block3a10),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a42),
	.cin(gnd),
	.combout(\ram_rom_data_reg[10]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[10]~10 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[10]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N30
cycloneive_lcell_comb \ram_rom_data_reg[11]~11 (
	.dataa(ram_block3a11),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a43),
	.cin(gnd),
	.combout(\ram_rom_data_reg[11]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[11]~11 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[11]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N12
cycloneive_lcell_comb \ram_rom_data_reg[12]~12 (
	.dataa(ram_block3a12),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a44),
	.cin(gnd),
	.combout(\ram_rom_data_reg[12]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[12]~12 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[12]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N26
cycloneive_lcell_comb \ram_rom_data_reg[13]~13 (
	.dataa(ram_block3a13),
	.datab(ram_block3a45),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[13]~13_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[13]~13 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[13]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N24
cycloneive_lcell_comb \ram_rom_data_reg[14]~14 (
	.dataa(ram_block3a14),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a46),
	.cin(gnd),
	.combout(\ram_rom_data_reg[14]~14_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[14]~14 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[14]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N20
cycloneive_lcell_comb \ram_rom_data_reg[15]~15 (
	.dataa(ram_block3a47),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a15),
	.cin(gnd),
	.combout(\ram_rom_data_reg[15]~15_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[15]~15 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[15]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N22
cycloneive_lcell_comb \ram_rom_data_reg[16]~16 (
	.dataa(ram_block3a16),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a48),
	.cin(gnd),
	.combout(\ram_rom_data_reg[16]~16_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[16]~16 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[16]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N0
cycloneive_lcell_comb \ram_rom_data_reg[17]~17 (
	.dataa(ram_block3a49),
	.datab(ram_block3a17),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[17]~17_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[17]~17 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[17]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N18
cycloneive_lcell_comb \ram_rom_data_reg[18]~18 (
	.dataa(ram_block3a50),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a18),
	.cin(gnd),
	.combout(\ram_rom_data_reg[18]~18_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[18]~18 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[18]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N8
cycloneive_lcell_comb \ram_rom_data_reg[19]~19 (
	.dataa(ram_block3a51),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a19),
	.cin(gnd),
	.combout(\ram_rom_data_reg[19]~19_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[19]~19 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[19]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N0
cycloneive_lcell_comb \ram_rom_data_reg[20]~20 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a20),
	.datac(gnd),
	.datad(ram_block3a52),
	.cin(gnd),
	.combout(\ram_rom_data_reg[20]~20_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[20]~20 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[20]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N30
cycloneive_lcell_comb \ram_rom_data_reg[21]~21 (
	.dataa(ram_block3a53),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a21),
	.cin(gnd),
	.combout(\ram_rom_data_reg[21]~21_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[21]~21 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[21]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N30
cycloneive_lcell_comb \ram_rom_data_reg[22]~22 (
	.dataa(ram_block3a22),
	.datab(ram_block3a54),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[22]~22_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[22]~22 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[22]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N24
cycloneive_lcell_comb \ram_rom_data_reg[23]~23 (
	.dataa(ram_block3a55),
	.datab(ram_block3a23),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[23]~23_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[23]~23 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[23]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N14
cycloneive_lcell_comb \ram_rom_data_reg[24]~24 (
	.dataa(ram_block3a56),
	.datab(ram_block3a24),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[24]~24_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[24]~24 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[24]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N8
cycloneive_lcell_comb \ram_rom_data_reg[25]~25 (
	.dataa(ram_block3a25),
	.datab(ram_block3a57),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[25]~25_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[25]~25 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[25]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N22
cycloneive_lcell_comb \ram_rom_data_reg[26]~26 (
	.dataa(ram_block3a58),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a26),
	.cin(gnd),
	.combout(\ram_rom_data_reg[26]~26_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[26]~26 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[26]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N12
cycloneive_lcell_comb \ram_rom_data_reg[27]~27 (
	.dataa(ram_block3a27),
	.datab(ram_block3a59),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[27]~27_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[27]~27 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[27]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N26
cycloneive_lcell_comb \ram_rom_data_reg[28]~28 (
	.dataa(ram_block3a28),
	.datab(ram_block3a60),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[28]~28_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[28]~28 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[28]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N16
cycloneive_lcell_comb \ram_rom_data_reg[29]~29 (
	.dataa(ram_block3a29),
	.datab(ram_block3a61),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[29]~29_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[29]~29 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[29]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N18
cycloneive_lcell_comb \ram_rom_data_reg[30]~30 (
	.dataa(ram_block3a62),
	.datab(ram_block3a30),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[30]~30_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[30]~30 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[30]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N4
cycloneive_lcell_comb \ram_rom_data_reg[31]~31 (
	.dataa(ram_block3a31),
	.datab(ram_block3a63),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[31]~31_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[31]~31 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[31]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y30_N8
cycloneive_lcell_comb \ir_loaded_address_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_0),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y30_N26
cycloneive_lcell_comb \process_0~0 (
	.dataa(irf_reg_4_1),
	.datab(gnd),
	.datac(gnd),
	.datad(ir_in[0]),
	.cin(gnd),
	.combout(\process_0~0_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~0 .lut_mask = 16'hFFAA;
defparam \process_0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y30_N16
cycloneive_lcell_comb \process_0~1 (
	.dataa(node_ena_1),
	.datab(virtual_ir_scan_reg),
	.datac(state_5),
	.datad(ir_in[3]),
	.cin(gnd),
	.combout(\process_0~1_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~1 .lut_mask = 16'h2000;
defparam \process_0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y30_N14
cycloneive_lcell_comb \ir_loaded_address_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_1),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y30_N22
cycloneive_lcell_comb \ir_loaded_address_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_3),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X41_Y30_N24
cycloneive_lcell_comb \bypass_reg_out~0 (
	.dataa(altera_internal_jtag),
	.datab(gnd),
	.datac(\bypass_reg_out~q ),
	.datad(node_ena_1),
	.cin(gnd),
	.combout(\bypass_reg_out~0_combout ),
	.cout());
// synopsys translate_off
defparam \bypass_reg_out~0 .lut_mask = 16'hAAF0;
defparam \bypass_reg_out~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X41_Y30_N25
dffeas bypass_reg_out(
	.clk(raw_tck),
	.d(\bypass_reg_out~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\bypass_reg_out~q ),
	.prn(vcc));
// synopsys translate_off
defparam bypass_reg_out.is_wysiwyg = "true";
defparam bypass_reg_out.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X41_Y30_N6
cycloneive_lcell_comb \tdo~0 (
	.dataa(irf_reg_1_1),
	.datab(ram_rom_data_reg_0),
	.datac(irf_reg_2_1),
	.datad(\bypass_reg_out~q ),
	.cin(gnd),
	.combout(\tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \tdo~0 .lut_mask = 16'hCDC8;
defparam \tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_rom_sr (
	WORD_SR_0,
	sdr,
	altera_internal_jtag,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	TCK,
	devpor,
	devclrn,
	devoe);
output 	WORD_SR_0;
input 	sdr;
input 	altera_internal_jtag;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	TCK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \word_counter[2]~11_combout ;
wire \WORD_SR~2_combout ;
wire \WORD_SR~7_combout ;
wire \WORD_SR~8_combout ;
wire \word_counter[1]~13_combout ;
wire \WORD_SR~10_combout ;
wire \WORD_SR~11_combout ;
wire \clear_signal~combout ;
wire \word_counter[0]~8 ;
wire \word_counter[1]~9_combout ;
wire \word_counter[0]~7_combout ;
wire \word_counter[1]~14_combout ;
wire \word_counter[1]~19_combout ;
wire \word_counter[1]~10 ;
wire \word_counter[2]~12 ;
wire \word_counter[3]~15_combout ;
wire \word_counter[3]~16 ;
wire \word_counter[4]~17_combout ;
wire \WORD_SR~13_combout ;
wire \WORD_SR~14_combout ;
wire \WORD_SR~15_combout ;
wire \WORD_SR[3]~6_combout ;
wire \WORD_SR~12_combout ;
wire \WORD_SR~9_combout ;
wire \WORD_SR~3_combout ;
wire \WORD_SR~4_combout ;
wire \WORD_SR~5_combout ;
wire [4:0] word_counter;
wire [3:0] WORD_SR;


// Location: FF_X33_Y32_N27
dffeas \word_counter[2] (
	.clk(TCK),
	.d(\word_counter[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[1]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[1]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[2]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[2] .is_wysiwyg = "true";
defparam \word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X33_Y32_N26
cycloneive_lcell_comb \word_counter[2]~11 (
	.dataa(word_counter[2]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[1]~10 ),
	.combout(\word_counter[2]~11_combout ),
	.cout(\word_counter[2]~12 ));
// synopsys translate_off
defparam \word_counter[2]~11 .lut_mask = 16'hA50A;
defparam \word_counter[2]~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X32_Y32_N12
cycloneive_lcell_comb \WORD_SR~2 (
	.dataa(word_counter[2]),
	.datab(word_counter[3]),
	.datac(word_counter[4]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~2_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~2 .lut_mask = 16'h0819;
defparam \WORD_SR~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X33_Y32_N12
cycloneive_lcell_comb \WORD_SR~7 (
	.dataa(word_counter[4]),
	.datab(word_counter[1]),
	.datac(word_counter[0]),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~7 .lut_mask = 16'h000D;
defparam \WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X33_Y32_N10
cycloneive_lcell_comb \WORD_SR~8 (
	.dataa(\WORD_SR~7_combout ),
	.datab(gnd),
	.datac(word_counter[2]),
	.datad(word_counter[3]),
	.cin(gnd),
	.combout(\WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~8 .lut_mask = 16'h000A;
defparam \WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X32_Y32_N2
cycloneive_lcell_comb \word_counter[1]~13 (
	.dataa(word_counter[2]),
	.datab(word_counter[3]),
	.datac(word_counter[4]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\word_counter[1]~13_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[1]~13 .lut_mask = 16'hFFDF;
defparam \word_counter[1]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X32_Y32_N0
cycloneive_lcell_comb \WORD_SR~10 (
	.dataa(word_counter[2]),
	.datab(word_counter[0]),
	.datac(word_counter[4]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~10 .lut_mask = 16'hD8F2;
defparam \WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X32_Y32_N14
cycloneive_lcell_comb \WORD_SR~11 (
	.dataa(\WORD_SR~2_combout ),
	.datab(\WORD_SR~10_combout ),
	.datac(gnd),
	.datad(word_counter[0]),
	.cin(gnd),
	.combout(\WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~11 .lut_mask = 16'hCC22;
defparam \WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X33_Y32_N21
dffeas \WORD_SR[0] (
	.clk(TCK),
	.d(\WORD_SR~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[3]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR_0),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[0] .is_wysiwyg = "true";
defparam \WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X33_Y32_N16
cycloneive_lcell_comb clear_signal(
	.dataa(gnd),
	.datab(gnd),
	.datac(state_8),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam clear_signal.lut_mask = 16'hF000;
defparam clear_signal.sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X33_Y32_N22
cycloneive_lcell_comb \word_counter[0]~7 (
	.dataa(word_counter[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\word_counter[0]~7_combout ),
	.cout(\word_counter[0]~8 ));
// synopsys translate_off
defparam \word_counter[0]~7 .lut_mask = 16'h55AA;
defparam \word_counter[0]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X33_Y32_N24
cycloneive_lcell_comb \word_counter[1]~9 (
	.dataa(gnd),
	.datab(word_counter[1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[0]~8 ),
	.combout(\word_counter[1]~9_combout ),
	.cout(\word_counter[1]~10 ));
// synopsys translate_off
defparam \word_counter[1]~9 .lut_mask = 16'h3C3F;
defparam \word_counter[1]~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X33_Y32_N2
cycloneive_lcell_comb \word_counter[1]~14 (
	.dataa(sdr),
	.datab(\clear_signal~combout ),
	.datac(state_3),
	.datad(state_4),
	.cin(gnd),
	.combout(\word_counter[1]~14_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[1]~14 .lut_mask = 16'hCCEC;
defparam \word_counter[1]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X33_Y32_N23
dffeas \word_counter[0] (
	.clk(TCK),
	.d(\word_counter[0]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[1]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[1]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[0]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[0] .is_wysiwyg = "true";
defparam \word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X33_Y32_N4
cycloneive_lcell_comb \word_counter[1]~19 (
	.dataa(\word_counter[1]~13_combout ),
	.datab(state_8),
	.datac(word_counter[0]),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\word_counter[1]~19_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[1]~19 .lut_mask = 16'hCD05;
defparam \word_counter[1]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X33_Y32_N25
dffeas \word_counter[1] (
	.clk(TCK),
	.d(\word_counter[1]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[1]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[1]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[1]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[1] .is_wysiwyg = "true";
defparam \word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X33_Y32_N28
cycloneive_lcell_comb \word_counter[3]~15 (
	.dataa(gnd),
	.datab(word_counter[3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[2]~12 ),
	.combout(\word_counter[3]~15_combout ),
	.cout(\word_counter[3]~16 ));
// synopsys translate_off
defparam \word_counter[3]~15 .lut_mask = 16'h3C3F;
defparam \word_counter[3]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X33_Y32_N29
dffeas \word_counter[3] (
	.clk(TCK),
	.d(\word_counter[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[1]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[1]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[3]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[3] .is_wysiwyg = "true";
defparam \word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X33_Y32_N30
cycloneive_lcell_comb \word_counter[4]~17 (
	.dataa(word_counter[4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\word_counter[3]~16 ),
	.combout(\word_counter[4]~17_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[4]~17 .lut_mask = 16'hA5A5;
defparam \word_counter[4]~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X33_Y32_N31
dffeas \word_counter[4] (
	.clk(TCK),
	.d(\word_counter[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[1]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[1]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[4]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[4] .is_wysiwyg = "true";
defparam \word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X32_Y32_N20
cycloneive_lcell_comb \WORD_SR~13 (
	.dataa(word_counter[2]),
	.datab(word_counter[3]),
	.datac(word_counter[4]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~13 .lut_mask = 16'h0800;
defparam \WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X33_Y32_N14
cycloneive_lcell_comb \WORD_SR~14 (
	.dataa(altera_internal_jtag),
	.datab(\WORD_SR~13_combout ),
	.datac(word_counter[0]),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~14 .lut_mask = 16'hAA0C;
defparam \WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X33_Y32_N0
cycloneive_lcell_comb \WORD_SR~15 (
	.dataa(gnd),
	.datab(state_8),
	.datac(\WORD_SR~14_combout ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\WORD_SR~15_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~15 .lut_mask = 16'h30F0;
defparam \WORD_SR~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X33_Y32_N18
cycloneive_lcell_comb \WORD_SR[3]~6 (
	.dataa(sdr),
	.datab(\clear_signal~combout ),
	.datac(state_3),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR[3]~6_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR[3]~6 .lut_mask = 16'hEEEC;
defparam \WORD_SR[3]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X33_Y32_N1
dffeas \WORD_SR[3] (
	.clk(TCK),
	.d(\WORD_SR~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[3]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[3]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[3] .is_wysiwyg = "true";
defparam \WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X33_Y32_N8
cycloneive_lcell_comb \WORD_SR~12 (
	.dataa(\WORD_SR~11_combout ),
	.datab(\clear_signal~combout ),
	.datac(WORD_SR[3]),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~12 .lut_mask = 16'h3022;
defparam \WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X33_Y32_N9
dffeas \WORD_SR[2] (
	.clk(TCK),
	.d(\WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[3]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[2]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[2] .is_wysiwyg = "true";
defparam \WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X33_Y32_N6
cycloneive_lcell_comb \WORD_SR~9 (
	.dataa(\WORD_SR~8_combout ),
	.datab(\clear_signal~combout ),
	.datac(WORD_SR[2]),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~9 .lut_mask = 16'h3222;
defparam \WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X33_Y32_N7
dffeas \WORD_SR[1] (
	.clk(TCK),
	.d(\WORD_SR~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[3]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[1]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[1] .is_wysiwyg = "true";
defparam \WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X32_Y32_N22
cycloneive_lcell_comb \WORD_SR~3 (
	.dataa(word_counter[2]),
	.datab(word_counter[0]),
	.datac(word_counter[4]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~3_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~3 .lut_mask = 16'hF210;
defparam \WORD_SR~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X32_Y32_N16
cycloneive_lcell_comb \WORD_SR~4 (
	.dataa(\WORD_SR~2_combout ),
	.datab(gnd),
	.datac(\WORD_SR~3_combout ),
	.datad(word_counter[0]),
	.cin(gnd),
	.combout(\WORD_SR~4_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~4 .lut_mask = 16'hF0A0;
defparam \WORD_SR~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X33_Y32_N20
cycloneive_lcell_comb \WORD_SR~5 (
	.dataa(WORD_SR[1]),
	.datab(\clear_signal~combout ),
	.datac(\WORD_SR~4_combout ),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~5_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~5 .lut_mask = 16'h2230;
defparam \WORD_SR~5 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module singlecycle (
	pcifimemaddr_29,
	pcifimemaddr_28,
	pcifimemaddr_31,
	pcifimemaddr_30,
	daddr_1,
	pcifimemaddr_1,
	ruifdmemREN,
	ruifdmemWEN,
	daddr_0,
	pcifimemaddr_0,
	daddr_3,
	pcifimemaddr_3,
	daddr_2,
	pcifimemaddr_2,
	daddr_5,
	pcifimemaddr_5,
	daddr_4,
	pcifimemaddr_4,
	daddr_7,
	pcifimemaddr_7,
	daddr_6,
	pcifimemaddr_6,
	daddr_9,
	pcifimemaddr_9,
	pcifimemaddr_8,
	daddr_8,
	daddr_11,
	pcifimemaddr_11,
	pcifimemaddr_10,
	daddr_10,
	daddr_13,
	pcifimemaddr_13,
	daddr_12,
	pcifimemaddr_12,
	daddr_15,
	pcifimemaddr_15,
	daddr_14,
	pcifimemaddr_14,
	daddr_17,
	pcifimemaddr_17,
	pcifimemaddr_16,
	daddr_16,
	daddr_19,
	pcifimemaddr_19,
	daddr_18,
	pcifimemaddr_18,
	daddr_21,
	pcifimemaddr_21,
	daddr_20,
	pcifimemaddr_20,
	daddr_23,
	pcifimemaddr_23,
	daddr_22,
	pcifimemaddr_22,
	daddr_25,
	pcifimemaddr_25,
	daddr_24,
	pcifimemaddr_24,
	daddr_27,
	pcifimemaddr_27,
	daddr_26,
	pcifimemaddr_26,
	daddr_29,
	daddr_28,
	daddr_31,
	daddr_30,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	Mux63,
	Mux631,
	cuifregT_4,
	Mux32,
	Mux321,
	Mux33,
	Mux331,
	Mux34,
	Mux341,
	Mux35,
	Mux351,
	Mux36,
	Mux361,
	Mux37,
	Mux371,
	Mux38,
	Mux381,
	Mux39,
	Mux391,
	Mux40,
	Mux401,
	Mux41,
	Mux411,
	Mux42,
	Mux421,
	Mux43,
	Mux431,
	Mux58,
	Mux581,
	Mux44,
	Mux441,
	Mux45,
	Mux451,
	Mux46,
	Mux461,
	Mux47,
	Mux471,
	Mux48,
	Mux481,
	Mux49,
	Mux491,
	Mux50,
	Mux501,
	Mux51,
	Mux511,
	Mux52,
	Mux521,
	Mux53,
	Mux531,
	Mux54,
	Mux541,
	Mux55,
	Mux551,
	Mux56,
	Mux561,
	Mux57,
	Mux571,
	Mux62,
	Mux621,
	Mux61,
	Mux611,
	Mux60,
	Mux601,
	Mux59,
	Mux591,
	ramiframload_261,
	ramiframload_271,
	ramiframload_281,
	ramiframload_291,
	ramiframload_301,
	ramiframload_311,
	nRST,
	CLK,
	nRST1,
	dpifhalt,
	devpor,
	devclrn,
	devoe);
output 	pcifimemaddr_29;
output 	pcifimemaddr_28;
output 	pcifimemaddr_31;
output 	pcifimemaddr_30;
output 	daddr_1;
output 	pcifimemaddr_1;
output 	ruifdmemREN;
output 	ruifdmemWEN;
output 	daddr_0;
output 	pcifimemaddr_0;
output 	daddr_3;
output 	pcifimemaddr_3;
output 	daddr_2;
output 	pcifimemaddr_2;
output 	daddr_5;
output 	pcifimemaddr_5;
output 	daddr_4;
output 	pcifimemaddr_4;
output 	daddr_7;
output 	pcifimemaddr_7;
output 	daddr_6;
output 	pcifimemaddr_6;
output 	daddr_9;
output 	pcifimemaddr_9;
output 	pcifimemaddr_8;
output 	daddr_8;
output 	daddr_11;
output 	pcifimemaddr_11;
output 	pcifimemaddr_10;
output 	daddr_10;
output 	daddr_13;
output 	pcifimemaddr_13;
output 	daddr_12;
output 	pcifimemaddr_12;
output 	daddr_15;
output 	pcifimemaddr_15;
output 	daddr_14;
output 	pcifimemaddr_14;
output 	daddr_17;
output 	pcifimemaddr_17;
output 	pcifimemaddr_16;
output 	daddr_16;
output 	daddr_19;
output 	pcifimemaddr_19;
output 	daddr_18;
output 	pcifimemaddr_18;
output 	daddr_21;
output 	pcifimemaddr_21;
output 	daddr_20;
output 	pcifimemaddr_20;
output 	daddr_23;
output 	pcifimemaddr_23;
output 	daddr_22;
output 	pcifimemaddr_22;
output 	daddr_25;
output 	pcifimemaddr_25;
output 	daddr_24;
output 	pcifimemaddr_24;
output 	daddr_27;
output 	pcifimemaddr_27;
output 	daddr_26;
output 	pcifimemaddr_26;
output 	daddr_29;
output 	daddr_28;
output 	daddr_31;
output 	daddr_30;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
output 	Mux63;
output 	Mux631;
output 	cuifregT_4;
output 	Mux32;
output 	Mux321;
output 	Mux33;
output 	Mux331;
output 	Mux34;
output 	Mux341;
output 	Mux35;
output 	Mux351;
output 	Mux36;
output 	Mux361;
output 	Mux37;
output 	Mux371;
output 	Mux38;
output 	Mux381;
output 	Mux39;
output 	Mux391;
output 	Mux40;
output 	Mux401;
output 	Mux41;
output 	Mux411;
output 	Mux42;
output 	Mux421;
output 	Mux43;
output 	Mux431;
output 	Mux58;
output 	Mux581;
output 	Mux44;
output 	Mux441;
output 	Mux45;
output 	Mux451;
output 	Mux46;
output 	Mux461;
output 	Mux47;
output 	Mux471;
output 	Mux48;
output 	Mux481;
output 	Mux49;
output 	Mux491;
output 	Mux50;
output 	Mux501;
output 	Mux51;
output 	Mux511;
output 	Mux52;
output 	Mux521;
output 	Mux53;
output 	Mux531;
output 	Mux54;
output 	Mux541;
output 	Mux55;
output 	Mux551;
output 	Mux56;
output 	Mux561;
output 	Mux57;
output 	Mux571;
output 	Mux62;
output 	Mux621;
output 	Mux61;
output 	Mux611;
output 	Mux60;
output 	Mux601;
output 	Mux59;
output 	Mux591;
input 	ramiframload_261;
input 	ramiframload_271;
input 	ramiframload_281;
input 	ramiframload_291;
input 	ramiframload_301;
input 	ramiframload_311;
input 	nRST;
input 	CLK;
input 	nRST1;
output 	dpifhalt;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \CC|iwait~0_combout ;
wire \CM|dcif.imemload[30]~2_combout ;
wire \CM|dcif.imemload[31]~3_combout ;
wire \CM|dcif.imemload[19]~4_combout ;
wire \CM|dcif.imemload[29]~5_combout ;
wire \CM|dcif.imemload[28]~6_combout ;
wire \CM|dcif.imemload[26]~7_combout ;
wire \CM|dcif.imemload[27]~8_combout ;
wire \CM|dcif.imemload[18]~9_combout ;
wire \CM|dcif.imemload[16]~10_combout ;
wire \CM|dcif.imemload[17]~11_combout ;
wire \CM|dcif.imemload[20]~12_combout ;
wire \CM|dcif.imemload[3]~13_combout ;
wire \CM|dcif.imemload[4]~14_combout ;
wire \CM|dcif.imemload[0]~15_combout ;
wire \CM|dcif.imemload[1]~16_combout ;
wire \CM|dcif.imemload[2]~17_combout ;
wire \CM|dcif.imemload[5]~18_combout ;
wire \CM|dcif.imemload[15]~19_combout ;
wire \CM|dcif.imemload[14]~20_combout ;
wire \CM|dcif.imemload[13]~21_combout ;
wire \CM|dcif.imemload[12]~22_combout ;
wire \CM|dcif.imemload[11]~23_combout ;
wire \CM|dcif.imemload[10]~24_combout ;
wire \CM|dcif.imemload[9]~25_combout ;
wire \CM|dcif.imemload[8]~26_combout ;
wire \CM|dcif.imemload[7]~27_combout ;
wire \CM|dcif.imemload[6]~28_combout ;
wire \CM|dcif.imemload[23]~29_combout ;
wire \CM|dcif.imemload[24]~30_combout ;
wire \CM|dcif.imemload[21]~31_combout ;
wire \CM|dcif.imemload[22]~32_combout ;
wire \CM|dcif.imemload[25]~33_combout ;
wire \DP|rf_dut|Mux31~20_combout ;
wire \DP|alu_dut|Selector30~8_combout ;
wire \DP|alu_dut|ShiftRight0~100_combout ;
wire \DP|alu_dut|Selector31~6_combout ;
wire \DP|alu_dut|Selector31~8_combout ;
wire \DP|alu_dut|Selector28~11_combout ;
wire \CM|dcif.imemload[26]~34_combout ;
wire \DP|alu_dut|ShiftLeft0~60_combout ;
wire \DP|alu_dut|Selector0~38_combout ;
wire \DP|alu_dut|ShiftLeft0~69_combout ;
wire \DP|alu_dut|Selector2~13_combout ;
wire \DP|alu_dut|Selector29~10_combout ;
wire \DP|alu_dut|Selector4~0_combout ;
wire \DP|alu_dut|Selector5~10_combout ;
wire \DP|alu_dut|ShiftLeft0~90_combout ;
wire \DP|alu_dut|Selector3~8_combout ;
wire \DP|alu_dut|ShiftLeft0~94_combout ;
wire \DP|alu_dut|Selector1~11_combout ;
wire \DP|alu_dut|Selector4~9_combout ;
wire \DP|alu_dut|Selector10~9_combout ;
wire \DP|alu_dut|Selector6~8_combout ;
wire \DP|alu_dut|Selector7~7_combout ;
wire \DP|alu_dut|Selector11~9_combout ;
wire \DP|alu_dut|Selector24~7_combout ;
wire \DP|alu_dut|Selector24~8_combout ;
wire \DP|alu_dut|Selector25~6_combout ;
wire \DP|alu_dut|Selector13~8_combout ;
wire \DP|alu_dut|Selector12~8_combout ;
wire \DP|alu_dut|Selector26~6_combout ;
wire \DP|alu_dut|Selector27~7_combout ;
wire \DP|alu_dut|Selector14~8_combout ;
wire \DP|alu_dut|Selector15~8_combout ;
wire \DP|alu_dut|Selector16~11_combout ;
wire \DP|alu_dut|Selector17~7_combout ;
wire \DP|alu_dut|Selector20~9_combout ;
wire \DP|alu_dut|Selector21~8_combout ;
wire \DP|alu_dut|Selector18~7_combout ;
wire \DP|alu_dut|Selector19~7_combout ;
wire \DP|alu_dut|Selector8~2_combout ;
wire \DP|alu_dut|Selector8~3_combout ;
wire \DP|alu_dut|Selector8~10_combout ;
wire \DP|alu_dut|Selector9~9_combout ;
wire \DP|alu_dut|Selector22~8_combout ;
wire \DP|alu_dut|Selector23~8_combout ;
wire \CM|dcif.dhit~2_combout ;
wire \CM|dcif.imemload[26]~35_combout ;
wire [31:0] \CM|instr ;


memory_control CC(
	.ruifdmemREN(ruifdmemREN),
	.ruifdmemWEN(ruifdmemWEN),
	.iwait(\CC|iwait~0_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

caches CM(
	.daddr_1(daddr_1),
	.ruifdmemREN(ruifdmemREN),
	.ruifdmemWEN(ruifdmemWEN),
	.daddr_0(daddr_0),
	.daddr_3(daddr_3),
	.daddr_2(daddr_2),
	.daddr_5(daddr_5),
	.daddr_4(daddr_4),
	.daddr_7(daddr_7),
	.daddr_6(daddr_6),
	.daddr_9(daddr_9),
	.daddr_8(daddr_8),
	.daddr_11(daddr_11),
	.daddr_10(daddr_10),
	.daddr_13(daddr_13),
	.daddr_12(daddr_12),
	.daddr_15(daddr_15),
	.daddr_14(daddr_14),
	.daddr_17(daddr_17),
	.daddr_16(daddr_16),
	.daddr_19(daddr_19),
	.daddr_18(daddr_18),
	.daddr_21(daddr_21),
	.daddr_20(daddr_20),
	.daddr_23(daddr_23),
	.daddr_22(daddr_22),
	.daddr_25(daddr_25),
	.daddr_24(daddr_24),
	.daddr_27(daddr_27),
	.daddr_26(daddr_26),
	.daddr_29(daddr_29),
	.daddr_28(daddr_28),
	.daddr_31(daddr_31),
	.daddr_30(daddr_30),
	.always1(always1),
	.ramiframload_0(ramiframload_0),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.iwait(\CC|iwait~0_combout ),
	.instr_28(\CM|instr [28]),
	.instr_27(\CM|instr [27]),
	.instr_29(\CM|instr [29]),
	.instr_26(\CM|instr [26]),
	.instr_30(\CM|instr [30]),
	.dcifimemload_30(\CM|dcif.imemload[30]~2_combout ),
	.instr_31(\CM|instr [31]),
	.dcifimemload_31(\CM|dcif.imemload[31]~3_combout ),
	.dcifimemload_19(\CM|dcif.imemload[19]~4_combout ),
	.dcifimemload_29(\CM|dcif.imemload[29]~5_combout ),
	.dcifimemload_28(\CM|dcif.imemload[28]~6_combout ),
	.dcifimemload_26(\CM|dcif.imemload[26]~7_combout ),
	.dcifimemload_27(\CM|dcif.imemload[27]~8_combout ),
	.dcifimemload_18(\CM|dcif.imemload[18]~9_combout ),
	.dcifimemload_16(\CM|dcif.imemload[16]~10_combout ),
	.dcifimemload_17(\CM|dcif.imemload[17]~11_combout ),
	.dcifimemload_20(\CM|dcif.imemload[20]~12_combout ),
	.dcifimemload_3(\CM|dcif.imemload[3]~13_combout ),
	.dcifimemload_4(\CM|dcif.imemload[4]~14_combout ),
	.dcifimemload_0(\CM|dcif.imemload[0]~15_combout ),
	.dcifimemload_1(\CM|dcif.imemload[1]~16_combout ),
	.dcifimemload_2(\CM|dcif.imemload[2]~17_combout ),
	.dcifimemload_5(\CM|dcif.imemload[5]~18_combout ),
	.dcifimemload_15(\CM|dcif.imemload[15]~19_combout ),
	.dcifimemload_14(\CM|dcif.imemload[14]~20_combout ),
	.dcifimemload_13(\CM|dcif.imemload[13]~21_combout ),
	.dcifimemload_12(\CM|dcif.imemload[12]~22_combout ),
	.dcifimemload_11(\CM|dcif.imemload[11]~23_combout ),
	.dcifimemload_10(\CM|dcif.imemload[10]~24_combout ),
	.dcifimemload_9(\CM|dcif.imemload[9]~25_combout ),
	.dcifimemload_8(\CM|dcif.imemload[8]~26_combout ),
	.dcifimemload_7(\CM|dcif.imemload[7]~27_combout ),
	.dcifimemload_6(\CM|dcif.imemload[6]~28_combout ),
	.dcifimemload_23(\CM|dcif.imemload[23]~29_combout ),
	.dcifimemload_24(\CM|dcif.imemload[24]~30_combout ),
	.dcifimemload_21(\CM|dcif.imemload[21]~31_combout ),
	.dcifimemload_22(\CM|dcif.imemload[22]~32_combout ),
	.dcifimemload_25(\CM|dcif.imemload[25]~33_combout ),
	.Mux31(\DP|rf_dut|Mux31~20_combout ),
	.Selector30(\DP|alu_dut|Selector30~8_combout ),
	.ShiftRight0(\DP|alu_dut|ShiftRight0~100_combout ),
	.Selector31(\DP|alu_dut|Selector31~6_combout ),
	.Selector311(\DP|alu_dut|Selector31~8_combout ),
	.Selector28(\DP|alu_dut|Selector28~11_combout ),
	.dcifimemload_261(\CM|dcif.imemload[26]~34_combout ),
	.ShiftLeft0(\DP|alu_dut|ShiftLeft0~60_combout ),
	.Selector0(\DP|alu_dut|Selector0~38_combout ),
	.ShiftLeft01(\DP|alu_dut|ShiftLeft0~69_combout ),
	.Selector2(\DP|alu_dut|Selector2~13_combout ),
	.Selector29(\DP|alu_dut|Selector29~10_combout ),
	.Selector4(\DP|alu_dut|Selector4~0_combout ),
	.Selector5(\DP|alu_dut|Selector5~10_combout ),
	.ShiftLeft02(\DP|alu_dut|ShiftLeft0~90_combout ),
	.Selector3(\DP|alu_dut|Selector3~8_combout ),
	.ShiftLeft03(\DP|alu_dut|ShiftLeft0~94_combout ),
	.Selector1(\DP|alu_dut|Selector1~11_combout ),
	.Selector41(\DP|alu_dut|Selector4~9_combout ),
	.Selector10(\DP|alu_dut|Selector10~9_combout ),
	.Selector6(\DP|alu_dut|Selector6~8_combout ),
	.Selector7(\DP|alu_dut|Selector7~7_combout ),
	.Selector11(\DP|alu_dut|Selector11~9_combout ),
	.Selector24(\DP|alu_dut|Selector24~7_combout ),
	.Selector241(\DP|alu_dut|Selector24~8_combout ),
	.Selector25(\DP|alu_dut|Selector25~6_combout ),
	.Selector13(\DP|alu_dut|Selector13~8_combout ),
	.Selector12(\DP|alu_dut|Selector12~8_combout ),
	.Selector26(\DP|alu_dut|Selector26~6_combout ),
	.Selector27(\DP|alu_dut|Selector27~7_combout ),
	.Selector14(\DP|alu_dut|Selector14~8_combout ),
	.Selector15(\DP|alu_dut|Selector15~8_combout ),
	.Selector16(\DP|alu_dut|Selector16~11_combout ),
	.Selector17(\DP|alu_dut|Selector17~7_combout ),
	.Selector20(\DP|alu_dut|Selector20~9_combout ),
	.Selector21(\DP|alu_dut|Selector21~8_combout ),
	.Selector18(\DP|alu_dut|Selector18~7_combout ),
	.Selector19(\DP|alu_dut|Selector19~7_combout ),
	.Selector8(\DP|alu_dut|Selector8~2_combout ),
	.Selector81(\DP|alu_dut|Selector8~3_combout ),
	.Selector82(\DP|alu_dut|Selector8~10_combout ),
	.Selector9(\DP|alu_dut|Selector9~9_combout ),
	.Selector22(\DP|alu_dut|Selector22~8_combout ),
	.Selector23(\DP|alu_dut|Selector23~8_combout ),
	.dcifdhit(\CM|dcif.dhit~2_combout ),
	.dcifimemload_262(\CM|dcif.imemload[26]~35_combout ),
	.nRST(nRST),
	.CLK(CLK),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

datapath DP(
	.pcifimemaddr_29(pcifimemaddr_29),
	.pcifimemaddr_28(pcifimemaddr_28),
	.pcifimemaddr_31(pcifimemaddr_31),
	.pcifimemaddr_30(pcifimemaddr_30),
	.pcifimemaddr_1(pcifimemaddr_1),
	.ruifdmemREN(ruifdmemREN),
	.ruifdmemWEN(ruifdmemWEN),
	.pcifimemaddr_0(pcifimemaddr_0),
	.pcifimemaddr_3(pcifimemaddr_3),
	.pcifimemaddr_2(pcifimemaddr_2),
	.pcifimemaddr_5(pcifimemaddr_5),
	.pcifimemaddr_4(pcifimemaddr_4),
	.pcifimemaddr_7(pcifimemaddr_7),
	.pcifimemaddr_6(pcifimemaddr_6),
	.pcifimemaddr_9(pcifimemaddr_9),
	.pcifimemaddr_8(pcifimemaddr_8),
	.pcifimemaddr_11(pcifimemaddr_11),
	.pcifimemaddr_10(pcifimemaddr_10),
	.pcifimemaddr_13(pcifimemaddr_13),
	.pcifimemaddr_12(pcifimemaddr_12),
	.pcifimemaddr_15(pcifimemaddr_15),
	.pcifimemaddr_14(pcifimemaddr_14),
	.pcifimemaddr_17(pcifimemaddr_17),
	.pcifimemaddr_16(pcifimemaddr_16),
	.pcifimemaddr_19(pcifimemaddr_19),
	.pcifimemaddr_18(pcifimemaddr_18),
	.pcifimemaddr_21(pcifimemaddr_21),
	.pcifimemaddr_20(pcifimemaddr_20),
	.pcifimemaddr_23(pcifimemaddr_23),
	.pcifimemaddr_22(pcifimemaddr_22),
	.pcifimemaddr_25(pcifimemaddr_25),
	.pcifimemaddr_24(pcifimemaddr_24),
	.pcifimemaddr_27(pcifimemaddr_27),
	.pcifimemaddr_26(pcifimemaddr_26),
	.always1(always1),
	.ramiframload_0(ramiframload_0),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.iwait(\CC|iwait~0_combout ),
	.instr_28(\CM|instr [28]),
	.instr_27(\CM|instr [27]),
	.instr_29(\CM|instr [29]),
	.instr_26(\CM|instr [26]),
	.instr_30(\CM|instr [30]),
	.dcifimemload_30(\CM|dcif.imemload[30]~2_combout ),
	.instr_31(\CM|instr [31]),
	.dcifimemload_31(\CM|dcif.imemload[31]~3_combout ),
	.dcifimemload_19(\CM|dcif.imemload[19]~4_combout ),
	.dcifimemload_29(\CM|dcif.imemload[29]~5_combout ),
	.dcifimemload_28(\CM|dcif.imemload[28]~6_combout ),
	.dcifimemload_26(\CM|dcif.imemload[26]~7_combout ),
	.dcifimemload_27(\CM|dcif.imemload[27]~8_combout ),
	.dcifimemload_18(\CM|dcif.imemload[18]~9_combout ),
	.dcifimemload_16(\CM|dcif.imemload[16]~10_combout ),
	.dcifimemload_17(\CM|dcif.imemload[17]~11_combout ),
	.Mux63(Mux63),
	.Mux631(Mux631),
	.dcifimemload_20(\CM|dcif.imemload[20]~12_combout ),
	.cuifregT_4(cuifregT_4),
	.dcifimemload_3(\CM|dcif.imemload[3]~13_combout ),
	.dcifimemload_4(\CM|dcif.imemload[4]~14_combout ),
	.dcifimemload_0(\CM|dcif.imemload[0]~15_combout ),
	.dcifimemload_1(\CM|dcif.imemload[1]~16_combout ),
	.dcifimemload_2(\CM|dcif.imemload[2]~17_combout ),
	.dcifimemload_5(\CM|dcif.imemload[5]~18_combout ),
	.dcifimemload_15(\CM|dcif.imemload[15]~19_combout ),
	.Mux32(Mux32),
	.Mux321(Mux321),
	.Mux33(Mux33),
	.Mux331(Mux331),
	.Mux34(Mux34),
	.Mux341(Mux341),
	.Mux35(Mux35),
	.Mux351(Mux351),
	.Mux36(Mux36),
	.Mux361(Mux361),
	.Mux37(Mux37),
	.Mux371(Mux371),
	.Mux38(Mux38),
	.Mux381(Mux381),
	.Mux39(Mux39),
	.Mux391(Mux391),
	.Mux40(Mux40),
	.Mux401(Mux401),
	.Mux41(Mux41),
	.Mux411(Mux411),
	.Mux42(Mux42),
	.Mux421(Mux421),
	.Mux43(Mux43),
	.Mux431(Mux431),
	.Mux58(Mux58),
	.Mux581(Mux581),
	.Mux44(Mux44),
	.Mux441(Mux441),
	.Mux45(Mux45),
	.Mux451(Mux451),
	.Mux46(Mux46),
	.Mux461(Mux461),
	.Mux47(Mux47),
	.Mux471(Mux471),
	.Mux48(Mux48),
	.Mux481(Mux481),
	.dcifimemload_14(\CM|dcif.imemload[14]~20_combout ),
	.Mux49(Mux49),
	.Mux491(Mux491),
	.dcifimemload_13(\CM|dcif.imemload[13]~21_combout ),
	.Mux50(Mux50),
	.Mux501(Mux501),
	.dcifimemload_12(\CM|dcif.imemload[12]~22_combout ),
	.Mux51(Mux51),
	.Mux511(Mux511),
	.dcifimemload_11(\CM|dcif.imemload[11]~23_combout ),
	.Mux52(Mux52),
	.Mux521(Mux521),
	.dcifimemload_10(\CM|dcif.imemload[10]~24_combout ),
	.Mux53(Mux53),
	.Mux531(Mux531),
	.dcifimemload_9(\CM|dcif.imemload[9]~25_combout ),
	.Mux54(Mux54),
	.Mux541(Mux541),
	.dcifimemload_8(\CM|dcif.imemload[8]~26_combout ),
	.Mux55(Mux55),
	.Mux551(Mux551),
	.dcifimemload_7(\CM|dcif.imemload[7]~27_combout ),
	.Mux56(Mux56),
	.Mux561(Mux561),
	.dcifimemload_6(\CM|dcif.imemload[6]~28_combout ),
	.Mux57(Mux57),
	.Mux571(Mux571),
	.dcifimemload_23(\CM|dcif.imemload[23]~29_combout ),
	.dcifimemload_24(\CM|dcif.imemload[24]~30_combout ),
	.dcifimemload_21(\CM|dcif.imemload[21]~31_combout ),
	.dcifimemload_22(\CM|dcif.imemload[22]~32_combout ),
	.dcifimemload_25(\CM|dcif.imemload[25]~33_combout ),
	.Mux62(Mux62),
	.Mux621(Mux621),
	.Mux61(Mux61),
	.Mux611(Mux611),
	.Mux60(Mux60),
	.Mux601(Mux601),
	.Mux59(Mux59),
	.Mux591(Mux591),
	.Mux31(\DP|rf_dut|Mux31~20_combout ),
	.Selector30(\DP|alu_dut|Selector30~8_combout ),
	.ShiftRight0(\DP|alu_dut|ShiftRight0~100_combout ),
	.Selector31(\DP|alu_dut|Selector31~6_combout ),
	.Selector311(\DP|alu_dut|Selector31~8_combout ),
	.Selector28(\DP|alu_dut|Selector28~11_combout ),
	.dcifimemload_261(\CM|dcif.imemload[26]~34_combout ),
	.ShiftLeft0(\DP|alu_dut|ShiftLeft0~60_combout ),
	.Selector0(\DP|alu_dut|Selector0~38_combout ),
	.ShiftLeft01(\DP|alu_dut|ShiftLeft0~69_combout ),
	.Selector2(\DP|alu_dut|Selector2~13_combout ),
	.Selector29(\DP|alu_dut|Selector29~10_combout ),
	.Selector4(\DP|alu_dut|Selector4~0_combout ),
	.Selector5(\DP|alu_dut|Selector5~10_combout ),
	.ShiftLeft02(\DP|alu_dut|ShiftLeft0~90_combout ),
	.Selector3(\DP|alu_dut|Selector3~8_combout ),
	.ShiftLeft03(\DP|alu_dut|ShiftLeft0~94_combout ),
	.Selector1(\DP|alu_dut|Selector1~11_combout ),
	.Selector41(\DP|alu_dut|Selector4~9_combout ),
	.Selector10(\DP|alu_dut|Selector10~9_combout ),
	.Selector6(\DP|alu_dut|Selector6~8_combout ),
	.Selector7(\DP|alu_dut|Selector7~7_combout ),
	.Selector11(\DP|alu_dut|Selector11~9_combout ),
	.Selector24(\DP|alu_dut|Selector24~7_combout ),
	.Selector241(\DP|alu_dut|Selector24~8_combout ),
	.Selector25(\DP|alu_dut|Selector25~6_combout ),
	.Selector13(\DP|alu_dut|Selector13~8_combout ),
	.Selector12(\DP|alu_dut|Selector12~8_combout ),
	.Selector26(\DP|alu_dut|Selector26~6_combout ),
	.Selector27(\DP|alu_dut|Selector27~7_combout ),
	.Selector14(\DP|alu_dut|Selector14~8_combout ),
	.Selector15(\DP|alu_dut|Selector15~8_combout ),
	.Selector16(\DP|alu_dut|Selector16~11_combout ),
	.Selector17(\DP|alu_dut|Selector17~7_combout ),
	.Selector20(\DP|alu_dut|Selector20~9_combout ),
	.Selector21(\DP|alu_dut|Selector21~8_combout ),
	.Selector18(\DP|alu_dut|Selector18~7_combout ),
	.Selector19(\DP|alu_dut|Selector19~7_combout ),
	.Selector8(\DP|alu_dut|Selector8~2_combout ),
	.Selector81(\DP|alu_dut|Selector8~3_combout ),
	.Selector82(\DP|alu_dut|Selector8~10_combout ),
	.Selector9(\DP|alu_dut|Selector9~9_combout ),
	.Selector22(\DP|alu_dut|Selector22~8_combout ),
	.Selector23(\DP|alu_dut|Selector23~8_combout ),
	.ramiframload_261(ramiframload_261),
	.ramiframload_271(ramiframload_271),
	.ramiframload_281(ramiframload_281),
	.ramiframload_291(ramiframload_291),
	.ramiframload_301(ramiframload_301),
	.ramiframload_311(ramiframload_311),
	.dcifdhit(\CM|dcif.dhit~2_combout ),
	.dcifimemload_262(\CM|dcif.imemload[26]~35_combout ),
	.CLK(CLK),
	.nRST(nRST1),
	.dpifhalt(dpifhalt),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module caches (
	daddr_1,
	ruifdmemREN,
	ruifdmemWEN,
	daddr_0,
	daddr_3,
	daddr_2,
	daddr_5,
	daddr_4,
	daddr_7,
	daddr_6,
	daddr_9,
	daddr_8,
	daddr_11,
	daddr_10,
	daddr_13,
	daddr_12,
	daddr_15,
	daddr_14,
	daddr_17,
	daddr_16,
	daddr_19,
	daddr_18,
	daddr_21,
	daddr_20,
	daddr_23,
	daddr_22,
	daddr_25,
	daddr_24,
	daddr_27,
	daddr_26,
	daddr_29,
	daddr_28,
	daddr_31,
	daddr_30,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	iwait,
	instr_28,
	instr_27,
	instr_29,
	instr_26,
	instr_30,
	dcifimemload_30,
	instr_31,
	dcifimemload_31,
	dcifimemload_19,
	dcifimemload_29,
	dcifimemload_28,
	dcifimemload_26,
	dcifimemload_27,
	dcifimemload_18,
	dcifimemload_16,
	dcifimemload_17,
	dcifimemload_20,
	dcifimemload_3,
	dcifimemload_4,
	dcifimemload_0,
	dcifimemload_1,
	dcifimemload_2,
	dcifimemload_5,
	dcifimemload_15,
	dcifimemload_14,
	dcifimemload_13,
	dcifimemload_12,
	dcifimemload_11,
	dcifimemload_10,
	dcifimemload_9,
	dcifimemload_8,
	dcifimemload_7,
	dcifimemload_6,
	dcifimemload_23,
	dcifimemload_24,
	dcifimemload_21,
	dcifimemload_22,
	dcifimemload_25,
	Mux31,
	Selector30,
	ShiftRight0,
	Selector31,
	Selector311,
	Selector28,
	dcifimemload_261,
	ShiftLeft0,
	Selector0,
	ShiftLeft01,
	Selector2,
	Selector29,
	Selector4,
	Selector5,
	ShiftLeft02,
	Selector3,
	ShiftLeft03,
	Selector1,
	Selector41,
	Selector10,
	Selector6,
	Selector7,
	Selector11,
	Selector24,
	Selector241,
	Selector25,
	Selector13,
	Selector12,
	Selector26,
	Selector27,
	Selector14,
	Selector15,
	Selector16,
	Selector17,
	Selector20,
	Selector21,
	Selector18,
	Selector19,
	Selector8,
	Selector81,
	Selector82,
	Selector9,
	Selector22,
	Selector23,
	dcifdhit,
	dcifimemload_262,
	nRST,
	CLK,
	devpor,
	devclrn,
	devoe);
output 	daddr_1;
input 	ruifdmemREN;
input 	ruifdmemWEN;
output 	daddr_0;
output 	daddr_3;
output 	daddr_2;
output 	daddr_5;
output 	daddr_4;
output 	daddr_7;
output 	daddr_6;
output 	daddr_9;
output 	daddr_8;
output 	daddr_11;
output 	daddr_10;
output 	daddr_13;
output 	daddr_12;
output 	daddr_15;
output 	daddr_14;
output 	daddr_17;
output 	daddr_16;
output 	daddr_19;
output 	daddr_18;
output 	daddr_21;
output 	daddr_20;
output 	daddr_23;
output 	daddr_22;
output 	daddr_25;
output 	daddr_24;
output 	daddr_27;
output 	daddr_26;
output 	daddr_29;
output 	daddr_28;
output 	daddr_31;
output 	daddr_30;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
input 	iwait;
output 	instr_28;
output 	instr_27;
output 	instr_29;
output 	instr_26;
output 	instr_30;
output 	dcifimemload_30;
output 	instr_31;
output 	dcifimemload_31;
output 	dcifimemload_19;
output 	dcifimemload_29;
output 	dcifimemload_28;
output 	dcifimemload_26;
output 	dcifimemload_27;
output 	dcifimemload_18;
output 	dcifimemload_16;
output 	dcifimemload_17;
output 	dcifimemload_20;
output 	dcifimemload_3;
output 	dcifimemload_4;
output 	dcifimemload_0;
output 	dcifimemload_1;
output 	dcifimemload_2;
output 	dcifimemload_5;
output 	dcifimemload_15;
output 	dcifimemload_14;
output 	dcifimemload_13;
output 	dcifimemload_12;
output 	dcifimemload_11;
output 	dcifimemload_10;
output 	dcifimemload_9;
output 	dcifimemload_8;
output 	dcifimemload_7;
output 	dcifimemload_6;
output 	dcifimemload_23;
output 	dcifimemload_24;
output 	dcifimemload_21;
output 	dcifimemload_22;
output 	dcifimemload_25;
input 	Mux31;
input 	Selector30;
input 	ShiftRight0;
input 	Selector31;
input 	Selector311;
input 	Selector28;
output 	dcifimemload_261;
input 	ShiftLeft0;
input 	Selector0;
input 	ShiftLeft01;
input 	Selector2;
input 	Selector29;
input 	Selector4;
input 	Selector5;
input 	ShiftLeft02;
input 	Selector3;
input 	ShiftLeft03;
input 	Selector1;
input 	Selector41;
input 	Selector10;
input 	Selector6;
input 	Selector7;
input 	Selector11;
input 	Selector24;
input 	Selector241;
input 	Selector25;
input 	Selector13;
input 	Selector12;
input 	Selector26;
input 	Selector27;
input 	Selector14;
input 	Selector15;
input 	Selector16;
input 	Selector17;
input 	Selector20;
input 	Selector21;
input 	Selector18;
input 	Selector19;
input 	Selector8;
input 	Selector81;
input 	Selector82;
input 	Selector9;
input 	Selector22;
input 	Selector23;
output 	dcifdhit;
output 	dcifimemload_262;
input 	nRST;
input 	CLK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \daddr~2_combout ;
wire \daddr[31]~34_combout ;
wire \daddr~3_combout ;
wire \daddr~4_combout ;
wire \daddr~5_combout ;
wire \daddr~6_combout ;
wire \daddr~7_combout ;
wire \daddr~8_combout ;
wire \daddr~9_combout ;
wire \daddr~10_combout ;
wire \daddr~11_combout ;
wire \daddr~12_combout ;
wire \daddr~13_combout ;
wire \daddr~14_combout ;
wire \daddr~15_combout ;
wire \daddr~16_combout ;
wire \daddr~17_combout ;
wire \daddr~18_combout ;
wire \daddr~19_combout ;
wire \daddr~20_combout ;
wire \daddr~21_combout ;
wire \daddr~22_combout ;
wire \daddr~23_combout ;
wire \daddr~24_combout ;
wire \daddr~25_combout ;
wire \daddr~26_combout ;
wire \daddr~27_combout ;
wire \daddr~28_combout ;
wire \daddr~29_combout ;
wire \daddr~30_combout ;
wire \daddr~31_combout ;
wire \daddr~32_combout ;
wire \daddr~33_combout ;
wire \instr~52_combout ;
wire \instr~53_combout ;
wire \instr~54_combout ;
wire \instr~55_combout ;
wire \instr~56_combout ;
wire \instr~57_combout ;
wire \instr~58_combout ;
wire \instr~59_combout ;
wire \instr~60_combout ;
wire \instr~61_combout ;
wire \instr~62_combout ;
wire \instr~63_combout ;
wire \instr~64_combout ;
wire \instr~65_combout ;
wire \instr~66_combout ;
wire \instr~67_combout ;
wire \instr~68_combout ;
wire \instr~69_combout ;
wire \instr~70_combout ;
wire \instr~71_combout ;
wire \instr~72_combout ;
wire \instr~73_combout ;
wire \instr~74_combout ;
wire \instr~75_combout ;
wire \instr~76_combout ;
wire \instr~77_combout ;
wire \instr~78_combout ;
wire \instr~79_combout ;
wire \instr~80_combout ;
wire \instr~81_combout ;
wire \instr~82_combout ;
wire \instr~83_combout ;
wire [31:0] instr;


// Location: FF_X55_Y36_N13
dffeas \daddr[1] (
	.clk(CLK),
	.d(\daddr~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_1),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[1] .is_wysiwyg = "true";
defparam \daddr[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y36_N27
dffeas \daddr[0] (
	.clk(CLK),
	.d(\daddr~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_0),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[0] .is_wysiwyg = "true";
defparam \daddr[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N9
dffeas \daddr[3] (
	.clk(CLK),
	.d(\daddr~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_3),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[3] .is_wysiwyg = "true";
defparam \daddr[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N29
dffeas \daddr[2] (
	.clk(CLK),
	.d(\daddr~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_2),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[2] .is_wysiwyg = "true";
defparam \daddr[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N21
dffeas \daddr[5] (
	.clk(CLK),
	.d(\daddr~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_5),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[5] .is_wysiwyg = "true";
defparam \daddr[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N1
dffeas \daddr[4] (
	.clk(CLK),
	.d(\daddr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_4),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[4] .is_wysiwyg = "true";
defparam \daddr[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N13
dffeas \daddr[7] (
	.clk(CLK),
	.d(\daddr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_7),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[7] .is_wysiwyg = "true";
defparam \daddr[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N3
dffeas \daddr[6] (
	.clk(CLK),
	.d(\daddr~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_6),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[6] .is_wysiwyg = "true";
defparam \daddr[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N29
dffeas \daddr[9] (
	.clk(CLK),
	.d(\daddr~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_9),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[9] .is_wysiwyg = "true";
defparam \daddr[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N5
dffeas \daddr[8] (
	.clk(CLK),
	.d(\daddr~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_8),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[8] .is_wysiwyg = "true";
defparam \daddr[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N5
dffeas \daddr[11] (
	.clk(CLK),
	.d(\daddr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_11),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[11] .is_wysiwyg = "true";
defparam \daddr[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y36_N1
dffeas \daddr[10] (
	.clk(CLK),
	.d(\daddr~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_10),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[10] .is_wysiwyg = "true";
defparam \daddr[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N23
dffeas \daddr[13] (
	.clk(CLK),
	.d(\daddr~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_13),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[13] .is_wysiwyg = "true";
defparam \daddr[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N25
dffeas \daddr[12] (
	.clk(CLK),
	.d(\daddr~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_12),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[12] .is_wysiwyg = "true";
defparam \daddr[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N25
dffeas \daddr[15] (
	.clk(CLK),
	.d(\daddr~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_15),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[15] .is_wysiwyg = "true";
defparam \daddr[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N13
dffeas \daddr[14] (
	.clk(CLK),
	.d(\daddr~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_14),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[14] .is_wysiwyg = "true";
defparam \daddr[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N7
dffeas \daddr[17] (
	.clk(CLK),
	.d(\daddr~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_17),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[17] .is_wysiwyg = "true";
defparam \daddr[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y37_N25
dffeas \daddr[16] (
	.clk(CLK),
	.d(\daddr~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_16),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[16] .is_wysiwyg = "true";
defparam \daddr[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N9
dffeas \daddr[19] (
	.clk(CLK),
	.d(\daddr~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_19),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[19] .is_wysiwyg = "true";
defparam \daddr[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y38_N11
dffeas \daddr[18] (
	.clk(CLK),
	.d(\daddr~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_18),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[18] .is_wysiwyg = "true";
defparam \daddr[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N27
dffeas \daddr[21] (
	.clk(CLK),
	.d(\daddr~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_21),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[21] .is_wysiwyg = "true";
defparam \daddr[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y38_N17
dffeas \daddr[20] (
	.clk(CLK),
	.d(\daddr~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_20),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[20] .is_wysiwyg = "true";
defparam \daddr[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N7
dffeas \daddr[23] (
	.clk(CLK),
	.d(\daddr~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_23),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[23] .is_wysiwyg = "true";
defparam \daddr[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y39_N5
dffeas \daddr[22] (
	.clk(CLK),
	.d(\daddr~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_22),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[22] .is_wysiwyg = "true";
defparam \daddr[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N27
dffeas \daddr[25] (
	.clk(CLK),
	.d(\daddr~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_25),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[25] .is_wysiwyg = "true";
defparam \daddr[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y33_N15
dffeas \daddr[24] (
	.clk(CLK),
	.d(\daddr~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_24),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[24] .is_wysiwyg = "true";
defparam \daddr[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N1
dffeas \daddr[27] (
	.clk(CLK),
	.d(\daddr~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_27),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[27] .is_wysiwyg = "true";
defparam \daddr[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y38_N31
dffeas \daddr[26] (
	.clk(CLK),
	.d(\daddr~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_26),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[26] .is_wysiwyg = "true";
defparam \daddr[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N5
dffeas \daddr[29] (
	.clk(CLK),
	.d(\daddr~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_29),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[29] .is_wysiwyg = "true";
defparam \daddr[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N19
dffeas \daddr[28] (
	.clk(CLK),
	.d(\daddr~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_28),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[28] .is_wysiwyg = "true";
defparam \daddr[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N31
dffeas \daddr[31] (
	.clk(CLK),
	.d(\daddr~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_31),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[31] .is_wysiwyg = "true";
defparam \daddr[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y37_N5
dffeas \daddr[30] (
	.clk(CLK),
	.d(\daddr~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(daddr_30),
	.prn(vcc));
// synopsys translate_off
defparam \daddr[30] .is_wysiwyg = "true";
defparam \daddr[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N23
dffeas \instr[28] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~52_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_28),
	.prn(vcc));
// synopsys translate_off
defparam \instr[28] .is_wysiwyg = "true";
defparam \instr[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N13
dffeas \instr[27] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~53_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_27),
	.prn(vcc));
// synopsys translate_off
defparam \instr[27] .is_wysiwyg = "true";
defparam \instr[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N11
dffeas \instr[29] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~54_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_29),
	.prn(vcc));
// synopsys translate_off
defparam \instr[29] .is_wysiwyg = "true";
defparam \instr[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y35_N5
dffeas \instr[26] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~55_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_26),
	.prn(vcc));
// synopsys translate_off
defparam \instr[26] .is_wysiwyg = "true";
defparam \instr[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y35_N3
dffeas \instr[30] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~56_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_30),
	.prn(vcc));
// synopsys translate_off
defparam \instr[30] .is_wysiwyg = "true";
defparam \instr[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N22
cycloneive_lcell_comb \dcif.imemload[30]~2 (
// Equation(s):
// dcifimemload_30 = (always1 & ((iwait & ((instr_30))) # (!iwait & (ramiframload_30)))) # (!always1 & (((instr_30))))

	.dataa(ramiframload_30),
	.datab(always1),
	.datac(instr_30),
	.datad(iwait),
	.cin(gnd),
	.combout(dcifimemload_30),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[30]~2 .lut_mask = 16'hF0B8;
defparam \dcif.imemload[30]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y35_N1
dffeas \instr[31] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~57_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr_31),
	.prn(vcc));
// synopsys translate_off
defparam \instr[31] .is_wysiwyg = "true";
defparam \instr[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N26
cycloneive_lcell_comb \dcif.imemload[31]~3 (
// Equation(s):
// dcifimemload_31 = (always1 & ((iwait & (instr_31)) # (!iwait & ((ramiframload_31))))) # (!always1 & (instr_31))

	.dataa(instr_31),
	.datab(always1),
	.datac(ramiframload_31),
	.datad(iwait),
	.cin(gnd),
	.combout(dcifimemload_31),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[31]~3 .lut_mask = 16'hAAE2;
defparam \dcif.imemload[31]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N8
cycloneive_lcell_comb \dcif.imemload[19]~4 (
// Equation(s):
// dcifimemload_19 = (always1 & ((iwait & (instr[19])) # (!iwait & ((ramiframload_19))))) # (!always1 & (((instr[19]))))

	.dataa(always1),
	.datab(iwait),
	.datac(instr[19]),
	.datad(ramiframload_19),
	.cin(gnd),
	.combout(dcifimemload_19),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[19]~4 .lut_mask = 16'hF2D0;
defparam \dcif.imemload[19]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N10
cycloneive_lcell_comb \dcif.imemload[29]~5 (
// Equation(s):
// dcifimemload_29 = (iwait & (((instr_29)))) # (!iwait & ((always1 & ((ramiframload_29))) # (!always1 & (instr_29))))

	.dataa(iwait),
	.datab(always1),
	.datac(instr_29),
	.datad(ramiframload_29),
	.cin(gnd),
	.combout(dcifimemload_29),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[29]~5 .lut_mask = 16'hF4B0;
defparam \dcif.imemload[29]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N14
cycloneive_lcell_comb \dcif.imemload[28]~6 (
// Equation(s):
// dcifimemload_28 = (iwait & (((instr_28)))) # (!iwait & ((always1 & (ramiframload_28)) # (!always1 & ((instr_28)))))

	.dataa(ramiframload_28),
	.datab(iwait),
	.datac(always1),
	.datad(instr_28),
	.cin(gnd),
	.combout(dcifimemload_28),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[28]~6 .lut_mask = 16'hEF20;
defparam \dcif.imemload[28]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N28
cycloneive_lcell_comb \dcif.imemload[26]~7 (
// Equation(s):
// dcifimemload_26 = (iwait & (instr_26)) # (!iwait & ((always1 & ((ramiframload_26))) # (!always1 & (instr_26))))

	.dataa(instr_26),
	.datab(iwait),
	.datac(ramiframload_26),
	.datad(always1),
	.cin(gnd),
	.combout(dcifimemload_26),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[26]~7 .lut_mask = 16'hB8AA;
defparam \dcif.imemload[26]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N12
cycloneive_lcell_comb \dcif.imemload[27]~8 (
// Equation(s):
// dcifimemload_27 = (iwait & (((instr_27)))) # (!iwait & ((always1 & (ramiframload_27)) # (!always1 & ((instr_27)))))

	.dataa(iwait),
	.datab(ramiframload_27),
	.datac(instr_27),
	.datad(always1),
	.cin(gnd),
	.combout(dcifimemload_27),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[27]~8 .lut_mask = 16'hE4F0;
defparam \dcif.imemload[27]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N6
cycloneive_lcell_comb \dcif.imemload[18]~9 (
// Equation(s):
// dcifimemload_18 = (iwait & (((instr[18])))) # (!iwait & ((always1 & ((ramiframload_18))) # (!always1 & (instr[18]))))

	.dataa(iwait),
	.datab(always1),
	.datac(instr[18]),
	.datad(ramiframload_18),
	.cin(gnd),
	.combout(dcifimemload_18),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[18]~9 .lut_mask = 16'hF4B0;
defparam \dcif.imemload[18]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N0
cycloneive_lcell_comb \dcif.imemload[16]~10 (
// Equation(s):
// dcifimemload_16 = (always1 & ((iwait & (instr[16])) # (!iwait & ((ramiframload_16))))) # (!always1 & (((instr[16]))))

	.dataa(always1),
	.datab(iwait),
	.datac(instr[16]),
	.datad(ramiframload_16),
	.cin(gnd),
	.combout(dcifimemload_16),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[16]~10 .lut_mask = 16'hF2D0;
defparam \dcif.imemload[16]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N4
cycloneive_lcell_comb \dcif.imemload[17]~11 (
// Equation(s):
// dcifimemload_17 = (iwait & (((instr[17])))) # (!iwait & ((always1 & ((ramiframload_17))) # (!always1 & (instr[17]))))

	.dataa(iwait),
	.datab(always1),
	.datac(instr[17]),
	.datad(ramiframload_17),
	.cin(gnd),
	.combout(dcifimemload_17),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[17]~11 .lut_mask = 16'hF4B0;
defparam \dcif.imemload[17]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N20
cycloneive_lcell_comb \dcif.imemload[20]~12 (
// Equation(s):
// dcifimemload_20 = (iwait & (((instr[20])))) # (!iwait & ((always1 & (ramiframload_20)) # (!always1 & ((instr[20])))))

	.dataa(iwait),
	.datab(ramiframload_20),
	.datac(instr[20]),
	.datad(always1),
	.cin(gnd),
	.combout(dcifimemload_20),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[20]~12 .lut_mask = 16'hE4F0;
defparam \dcif.imemload[20]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N30
cycloneive_lcell_comb \dcif.imemload[3]~13 (
// Equation(s):
// dcifimemload_3 = (always1 & ((iwait & (instr[3])) # (!iwait & ((ramiframload_3))))) # (!always1 & (((instr[3]))))

	.dataa(always1),
	.datab(iwait),
	.datac(instr[3]),
	.datad(ramiframload_3),
	.cin(gnd),
	.combout(dcifimemload_3),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[3]~13 .lut_mask = 16'hF2D0;
defparam \dcif.imemload[3]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N0
cycloneive_lcell_comb \dcif.imemload[4]~14 (
// Equation(s):
// dcifimemload_4 = (always1 & ((iwait & ((instr[4]))) # (!iwait & (ramiframload_4)))) # (!always1 & (((instr[4]))))

	.dataa(always1),
	.datab(ramiframload_4),
	.datac(instr[4]),
	.datad(iwait),
	.cin(gnd),
	.combout(dcifimemload_4),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[4]~14 .lut_mask = 16'hF0D8;
defparam \dcif.imemload[4]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N16
cycloneive_lcell_comb \dcif.imemload[0]~15 (
// Equation(s):
// dcifimemload_0 = (iwait & (((instr[0])))) # (!iwait & ((always1 & (ramiframload_0)) # (!always1 & ((instr[0])))))

	.dataa(ramiframload_0),
	.datab(iwait),
	.datac(instr[0]),
	.datad(always1),
	.cin(gnd),
	.combout(dcifimemload_0),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[0]~15 .lut_mask = 16'hE2F0;
defparam \dcif.imemload[0]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N14
cycloneive_lcell_comb \dcif.imemload[1]~16 (
// Equation(s):
// dcifimemload_1 = (always1 & ((iwait & (instr[1])) # (!iwait & ((ramiframload_1))))) # (!always1 & (((instr[1]))))

	.dataa(always1),
	.datab(iwait),
	.datac(instr[1]),
	.datad(ramiframload_1),
	.cin(gnd),
	.combout(dcifimemload_1),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[1]~16 .lut_mask = 16'hF2D0;
defparam \dcif.imemload[1]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N14
cycloneive_lcell_comb \dcif.imemload[2]~17 (
// Equation(s):
// dcifimemload_2 = (always1 & ((iwait & (instr[2])) # (!iwait & ((ramiframload_2))))) # (!always1 & (((instr[2]))))

	.dataa(always1),
	.datab(iwait),
	.datac(instr[2]),
	.datad(ramiframload_2),
	.cin(gnd),
	.combout(dcifimemload_2),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[2]~17 .lut_mask = 16'hF2D0;
defparam \dcif.imemload[2]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N18
cycloneive_lcell_comb \dcif.imemload[5]~18 (
// Equation(s):
// dcifimemload_5 = (iwait & (((instr[5])))) # (!iwait & ((always1 & (ramiframload_5)) # (!always1 & ((instr[5])))))

	.dataa(ramiframload_5),
	.datab(iwait),
	.datac(instr[5]),
	.datad(always1),
	.cin(gnd),
	.combout(dcifimemload_5),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[5]~18 .lut_mask = 16'hE2F0;
defparam \dcif.imemload[5]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N20
cycloneive_lcell_comb \dcif.imemload[15]~19 (
// Equation(s):
// dcifimemload_15 = (always1 & ((iwait & (instr[15])) # (!iwait & ((ramiframload_15))))) # (!always1 & (((instr[15]))))

	.dataa(always1),
	.datab(iwait),
	.datac(instr[15]),
	.datad(ramiframload_15),
	.cin(gnd),
	.combout(dcifimemload_15),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[15]~19 .lut_mask = 16'hF2D0;
defparam \dcif.imemload[15]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N6
cycloneive_lcell_comb \dcif.imemload[14]~20 (
// Equation(s):
// dcifimemload_14 = (always1 & ((iwait & (instr[14])) # (!iwait & ((ramiframload_14))))) # (!always1 & (((instr[14]))))

	.dataa(always1),
	.datab(iwait),
	.datac(instr[14]),
	.datad(ramiframload_14),
	.cin(gnd),
	.combout(dcifimemload_14),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[14]~20 .lut_mask = 16'hF2D0;
defparam \dcif.imemload[14]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N28
cycloneive_lcell_comb \dcif.imemload[13]~21 (
// Equation(s):
// dcifimemload_13 = (iwait & (((instr[13])))) # (!iwait & ((always1 & (ramiframload_13)) # (!always1 & ((instr[13])))))

	.dataa(ramiframload_13),
	.datab(iwait),
	.datac(instr[13]),
	.datad(always1),
	.cin(gnd),
	.combout(dcifimemload_13),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[13]~21 .lut_mask = 16'hE2F0;
defparam \dcif.imemload[13]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N2
cycloneive_lcell_comb \dcif.imemload[12]~22 (
// Equation(s):
// dcifimemload_12 = (iwait & (((instr[12])))) # (!iwait & ((always1 & ((ramiframload_12))) # (!always1 & (instr[12]))))

	.dataa(iwait),
	.datab(always1),
	.datac(instr[12]),
	.datad(ramiframload_12),
	.cin(gnd),
	.combout(dcifimemload_12),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[12]~22 .lut_mask = 16'hF4B0;
defparam \dcif.imemload[12]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N30
cycloneive_lcell_comb \dcif.imemload[11]~23 (
// Equation(s):
// dcifimemload_11 = (always1 & ((iwait & ((instr[11]))) # (!iwait & (ramiframload_11)))) # (!always1 & (((instr[11]))))

	.dataa(always1),
	.datab(ramiframload_11),
	.datac(instr[11]),
	.datad(iwait),
	.cin(gnd),
	.combout(dcifimemload_11),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[11]~23 .lut_mask = 16'hF0D8;
defparam \dcif.imemload[11]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N8
cycloneive_lcell_comb \dcif.imemload[10]~24 (
// Equation(s):
// dcifimemload_10 = (iwait & (((instr[10])))) # (!iwait & ((always1 & (ramiframload_10)) # (!always1 & ((instr[10])))))

	.dataa(ramiframload_10),
	.datab(iwait),
	.datac(instr[10]),
	.datad(always1),
	.cin(gnd),
	.combout(dcifimemload_10),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[10]~24 .lut_mask = 16'hE2F0;
defparam \dcif.imemload[10]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N30
cycloneive_lcell_comb \dcif.imemload[9]~25 (
// Equation(s):
// dcifimemload_9 = (always1 & ((iwait & (instr[9])) # (!iwait & ((ramiframload_9))))) # (!always1 & (((instr[9]))))

	.dataa(always1),
	.datab(iwait),
	.datac(instr[9]),
	.datad(ramiframload_9),
	.cin(gnd),
	.combout(dcifimemload_9),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[9]~25 .lut_mask = 16'hF2D0;
defparam \dcif.imemload[9]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N30
cycloneive_lcell_comb \dcif.imemload[8]~26 (
// Equation(s):
// dcifimemload_8 = (iwait & (((instr[8])))) # (!iwait & ((always1 & ((ramiframload_8))) # (!always1 & (instr[8]))))

	.dataa(iwait),
	.datab(always1),
	.datac(instr[8]),
	.datad(ramiframload_8),
	.cin(gnd),
	.combout(dcifimemload_8),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[8]~26 .lut_mask = 16'hF4B0;
defparam \dcif.imemload[8]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N14
cycloneive_lcell_comb \dcif.imemload[7]~27 (
// Equation(s):
// dcifimemload_7 = (iwait & (((instr[7])))) # (!iwait & ((always1 & (ramiframload_7)) # (!always1 & ((instr[7])))))

	.dataa(iwait),
	.datab(ramiframload_7),
	.datac(instr[7]),
	.datad(always1),
	.cin(gnd),
	.combout(dcifimemload_7),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[7]~27 .lut_mask = 16'hE4F0;
defparam \dcif.imemload[7]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N16
cycloneive_lcell_comb \dcif.imemload[6]~28 (
// Equation(s):
// dcifimemload_6 = (iwait & (((instr[6])))) # (!iwait & ((always1 & (ramiframload_6)) # (!always1 & ((instr[6])))))

	.dataa(ramiframload_6),
	.datab(iwait),
	.datac(instr[6]),
	.datad(always1),
	.cin(gnd),
	.combout(dcifimemload_6),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[6]~28 .lut_mask = 16'hE2F0;
defparam \dcif.imemload[6]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N24
cycloneive_lcell_comb \dcif.imemload[23]~29 (
// Equation(s):
// dcifimemload_23 = (always1 & ((iwait & ((instr[23]))) # (!iwait & (ramiframload_23)))) # (!always1 & (((instr[23]))))

	.dataa(always1),
	.datab(ramiframload_23),
	.datac(instr[23]),
	.datad(iwait),
	.cin(gnd),
	.combout(dcifimemload_23),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[23]~29 .lut_mask = 16'hF0D8;
defparam \dcif.imemload[23]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N12
cycloneive_lcell_comb \dcif.imemload[24]~30 (
// Equation(s):
// dcifimemload_24 = (always1 & ((iwait & (instr[24])) # (!iwait & ((ramiframload_24))))) # (!always1 & (((instr[24]))))

	.dataa(always1),
	.datab(iwait),
	.datac(instr[24]),
	.datad(ramiframload_24),
	.cin(gnd),
	.combout(dcifimemload_24),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[24]~30 .lut_mask = 16'hF2D0;
defparam \dcif.imemload[24]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N16
cycloneive_lcell_comb \dcif.imemload[21]~31 (
// Equation(s):
// dcifimemload_21 = (always1 & ((iwait & (instr[21])) # (!iwait & ((ramiframload_21))))) # (!always1 & (((instr[21]))))

	.dataa(always1),
	.datab(iwait),
	.datac(instr[21]),
	.datad(ramiframload_21),
	.cin(gnd),
	.combout(dcifimemload_21),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[21]~31 .lut_mask = 16'hF2D0;
defparam \dcif.imemload[21]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N8
cycloneive_lcell_comb \dcif.imemload[22]~32 (
// Equation(s):
// dcifimemload_22 = (always1 & ((iwait & (instr[22])) # (!iwait & ((ramiframload_22))))) # (!always1 & (((instr[22]))))

	.dataa(always1),
	.datab(iwait),
	.datac(instr[22]),
	.datad(ramiframload_22),
	.cin(gnd),
	.combout(dcifimemload_22),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[22]~32 .lut_mask = 16'hF2D0;
defparam \dcif.imemload[22]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N24
cycloneive_lcell_comb \dcif.imemload[25]~33 (
// Equation(s):
// dcifimemload_25 = (always1 & ((iwait & (instr[25])) # (!iwait & ((ramiframload_25))))) # (!always1 & (((instr[25]))))

	.dataa(always1),
	.datab(iwait),
	.datac(instr[25]),
	.datad(ramiframload_25),
	.cin(gnd),
	.combout(dcifimemload_25),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[25]~33 .lut_mask = 16'hF2D0;
defparam \dcif.imemload[25]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N12
cycloneive_lcell_comb \dcif.imemload[26]~34 (
// Equation(s):
// dcifimemload_261 = (instr_26 & ((ruifdmemREN) # ((ruifdmemWEN) # (!always1))))

	.dataa(ruifdmemREN),
	.datab(always1),
	.datac(instr_26),
	.datad(ruifdmemWEN),
	.cin(gnd),
	.combout(dcifimemload_261),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[26]~34 .lut_mask = 16'hF0B0;
defparam \dcif.imemload[26]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N6
cycloneive_lcell_comb \dcif.dhit~2 (
// Equation(s):
// dcifdhit = ((!ruifdmemWEN & !ruifdmemREN)) # (!always1)

	.dataa(always1),
	.datab(ruifdmemWEN),
	.datac(gnd),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(dcifdhit),
	.cout());
// synopsys translate_off
defparam \dcif.dhit~2 .lut_mask = 16'h5577;
defparam \dcif.dhit~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N10
cycloneive_lcell_comb \dcif.imemload[26]~35 (
// Equation(s):
// dcifimemload_262 = (!ruifdmemWEN & (ramiframload_26 & (!ruifdmemREN & always1)))

	.dataa(ruifdmemWEN),
	.datab(ramiframload_26),
	.datac(ruifdmemREN),
	.datad(always1),
	.cin(gnd),
	.combout(dcifimemload_262),
	.cout());
// synopsys translate_off
defparam \dcif.imemload[26]~35 .lut_mask = 16'h0400;
defparam \dcif.imemload[26]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N12
cycloneive_lcell_comb \daddr~2 (
// Equation(s):
// \daddr~2_combout  = (Selector30 & \nRST~input_o )

	.dataa(gnd),
	.datab(Selector30),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~2_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~2 .lut_mask = 16'hCC00;
defparam \daddr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N24
cycloneive_lcell_comb \daddr[31]~34 (
// Equation(s):
// \daddr[31]~34_combout  = ((!ruifdmemWEN & (always1 & !ruifdmemREN))) # (!\nRST~input_o )

	.dataa(ruifdmemWEN),
	.datab(nRST),
	.datac(always1),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(\daddr[31]~34_combout ),
	.cout());
// synopsys translate_off
defparam \daddr[31]~34 .lut_mask = 16'h3373;
defparam \daddr[31]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N26
cycloneive_lcell_comb \daddr~3 (
// Equation(s):
// \daddr~3_combout  = (\nRST~input_o  & ((Selector31) # ((Mux31 & Selector311))))

	.dataa(Mux31),
	.datab(Selector311),
	.datac(Selector31),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~3_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~3 .lut_mask = 16'hF800;
defparam \daddr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N8
cycloneive_lcell_comb \daddr~4 (
// Equation(s):
// \daddr~4_combout  = (\nRST~input_o  & Selector28)

	.dataa(gnd),
	.datab(nRST),
	.datac(Selector28),
	.datad(gnd),
	.cin(gnd),
	.combout(\daddr~4_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~4 .lut_mask = 16'hC0C0;
defparam \daddr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N28
cycloneive_lcell_comb \daddr~5 (
// Equation(s):
// \daddr~5_combout  = (Selector29 & \nRST~input_o )

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector29),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~5_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~5 .lut_mask = 16'hF000;
defparam \daddr~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N20
cycloneive_lcell_comb \daddr~6 (
// Equation(s):
// \daddr~6_combout  = (\nRST~input_o  & ((Selector26) # ((ShiftLeft01 & Selector241))))

	.dataa(ShiftLeft01),
	.datab(nRST),
	.datac(Selector241),
	.datad(Selector26),
	.cin(gnd),
	.combout(\daddr~6_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~6 .lut_mask = 16'hCC80;
defparam \daddr~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N0
cycloneive_lcell_comb \daddr~7 (
// Equation(s):
// \daddr~7_combout  = (\nRST~input_o  & ((Selector27) # ((ShiftLeft02 & Selector241))))

	.dataa(Selector27),
	.datab(ShiftLeft02),
	.datac(Selector241),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~7_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~7 .lut_mask = 16'hEA00;
defparam \daddr~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N12
cycloneive_lcell_comb \daddr~8 (
// Equation(s):
// \daddr~8_combout  = (\nRST~input_o  & ((Selector24) # ((ShiftLeft0 & Selector241))))

	.dataa(nRST),
	.datab(ShiftLeft0),
	.datac(Selector241),
	.datad(Selector24),
	.cin(gnd),
	.combout(\daddr~8_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~8 .lut_mask = 16'hAA80;
defparam \daddr~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N2
cycloneive_lcell_comb \daddr~9 (
// Equation(s):
// \daddr~9_combout  = (\nRST~input_o  & ((Selector25) # ((Selector241 & ShiftLeft03))))

	.dataa(Selector25),
	.datab(nRST),
	.datac(Selector241),
	.datad(ShiftLeft03),
	.cin(gnd),
	.combout(\daddr~9_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~9 .lut_mask = 16'hC888;
defparam \daddr~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N28
cycloneive_lcell_comb \daddr~10 (
// Equation(s):
// \daddr~10_combout  = (\nRST~input_o  & Selector22)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(Selector22),
	.cin(gnd),
	.combout(\daddr~10_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~10 .lut_mask = 16'hF000;
defparam \daddr~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N4
cycloneive_lcell_comb \daddr~11 (
// Equation(s):
// \daddr~11_combout  = (Selector23 & \nRST~input_o )

	.dataa(Selector23),
	.datab(gnd),
	.datac(nRST),
	.datad(gnd),
	.cin(gnd),
	.combout(\daddr~11_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~11 .lut_mask = 16'hA0A0;
defparam \daddr~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N4
cycloneive_lcell_comb \daddr~12 (
// Equation(s):
// \daddr~12_combout  = (\nRST~input_o  & Selector20)

	.dataa(gnd),
	.datab(nRST),
	.datac(Selector20),
	.datad(gnd),
	.cin(gnd),
	.combout(\daddr~12_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~12 .lut_mask = 16'hC0C0;
defparam \daddr~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N0
cycloneive_lcell_comb \daddr~13 (
// Equation(s):
// \daddr~13_combout  = (\nRST~input_o  & Selector21)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(Selector21),
	.cin(gnd),
	.combout(\daddr~13_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~13 .lut_mask = 16'hF000;
defparam \daddr~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N22
cycloneive_lcell_comb \daddr~14 (
// Equation(s):
// \daddr~14_combout  = (\nRST~input_o  & Selector18)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(Selector18),
	.cin(gnd),
	.combout(\daddr~14_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~14 .lut_mask = 16'hF000;
defparam \daddr~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N24
cycloneive_lcell_comb \daddr~15 (
// Equation(s):
// \daddr~15_combout  = (\nRST~input_o  & Selector19)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(Selector19),
	.cin(gnd),
	.combout(\daddr~15_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~15 .lut_mask = 16'hCC00;
defparam \daddr~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N24
cycloneive_lcell_comb \daddr~16 (
// Equation(s):
// \daddr~16_combout  = (\nRST~input_o  & Selector16)

	.dataa(gnd),
	.datab(nRST),
	.datac(Selector16),
	.datad(gnd),
	.cin(gnd),
	.combout(\daddr~16_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~16 .lut_mask = 16'hC0C0;
defparam \daddr~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N12
cycloneive_lcell_comb \daddr~17 (
// Equation(s):
// \daddr~17_combout  = (\nRST~input_o  & Selector17)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(Selector17),
	.cin(gnd),
	.combout(\daddr~17_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~17 .lut_mask = 16'hCC00;
defparam \daddr~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N6
cycloneive_lcell_comb \daddr~18 (
// Equation(s):
// \daddr~18_combout  = (Selector14 & \nRST~input_o )

	.dataa(gnd),
	.datab(gnd),
	.datac(Selector14),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~18_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~18 .lut_mask = 16'hF000;
defparam \daddr~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N24
cycloneive_lcell_comb \daddr~19 (
// Equation(s):
// \daddr~19_combout  = (\nRST~input_o  & Selector15)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(Selector15),
	.cin(gnd),
	.combout(\daddr~19_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~19 .lut_mask = 16'hCC00;
defparam \daddr~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N8
cycloneive_lcell_comb \daddr~20 (
// Equation(s):
// \daddr~20_combout  = (\nRST~input_o  & Selector12)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(Selector12),
	.cin(gnd),
	.combout(\daddr~20_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~20 .lut_mask = 16'hF000;
defparam \daddr~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N10
cycloneive_lcell_comb \daddr~21 (
// Equation(s):
// \daddr~21_combout  = (\nRST~input_o  & Selector13)

	.dataa(gnd),
	.datab(nRST),
	.datac(Selector13),
	.datad(gnd),
	.cin(gnd),
	.combout(\daddr~21_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~21 .lut_mask = 16'hC0C0;
defparam \daddr~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N26
cycloneive_lcell_comb \daddr~22 (
// Equation(s):
// \daddr~22_combout  = (\nRST~input_o  & Selector10)

	.dataa(nRST),
	.datab(gnd),
	.datac(Selector10),
	.datad(gnd),
	.cin(gnd),
	.combout(\daddr~22_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~22 .lut_mask = 16'hA0A0;
defparam \daddr~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N16
cycloneive_lcell_comb \daddr~23 (
// Equation(s):
// \daddr~23_combout  = (Selector11 & \nRST~input_o )

	.dataa(gnd),
	.datab(Selector11),
	.datac(gnd),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~23_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~23 .lut_mask = 16'hCC00;
defparam \daddr~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N6
cycloneive_lcell_comb \daddr~24 (
// Equation(s):
// \daddr~24_combout  = (\nRST~input_o  & ((Selector81) # ((Selector8) # (Selector82))))

	.dataa(Selector81),
	.datab(Selector8),
	.datac(Selector82),
	.datad(nRST),
	.cin(gnd),
	.combout(\daddr~24_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~24 .lut_mask = 16'hFE00;
defparam \daddr~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N4
cycloneive_lcell_comb \daddr~25 (
// Equation(s):
// \daddr~25_combout  = (\nRST~input_o  & Selector9)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(Selector9),
	.cin(gnd),
	.combout(\daddr~25_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~25 .lut_mask = 16'hCC00;
defparam \daddr~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N26
cycloneive_lcell_comb \daddr~26 (
// Equation(s):
// \daddr~26_combout  = (\nRST~input_o  & Selector6)

	.dataa(gnd),
	.datab(nRST),
	.datac(gnd),
	.datad(Selector6),
	.cin(gnd),
	.combout(\daddr~26_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~26 .lut_mask = 16'hCC00;
defparam \daddr~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y33_N14
cycloneive_lcell_comb \daddr~27 (
// Equation(s):
// \daddr~27_combout  = (\nRST~input_o  & ((Selector7) # ((ShiftRight0 & Selector4))))

	.dataa(nRST),
	.datab(ShiftRight0),
	.datac(Selector4),
	.datad(Selector7),
	.cin(gnd),
	.combout(\daddr~27_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~27 .lut_mask = 16'hAA80;
defparam \daddr~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N0
cycloneive_lcell_comb \daddr~28 (
// Equation(s):
// \daddr~28_combout  = (\nRST~input_o  & Selector41)

	.dataa(gnd),
	.datab(nRST),
	.datac(Selector41),
	.datad(gnd),
	.cin(gnd),
	.combout(\daddr~28_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~28 .lut_mask = 16'hC0C0;
defparam \daddr~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y38_N30
cycloneive_lcell_comb \daddr~29 (
// Equation(s):
// \daddr~29_combout  = (\nRST~input_o  & Selector5)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(Selector5),
	.cin(gnd),
	.combout(\daddr~29_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~29 .lut_mask = 16'hF000;
defparam \daddr~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N4
cycloneive_lcell_comb \daddr~30 (
// Equation(s):
// \daddr~30_combout  = (\nRST~input_o  & Selector2)

	.dataa(gnd),
	.datab(nRST),
	.datac(Selector2),
	.datad(gnd),
	.cin(gnd),
	.combout(\daddr~30_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~30 .lut_mask = 16'hC0C0;
defparam \daddr~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N18
cycloneive_lcell_comb \daddr~31 (
// Equation(s):
// \daddr~31_combout  = (\nRST~input_o  & Selector3)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(Selector3),
	.cin(gnd),
	.combout(\daddr~31_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~31 .lut_mask = 16'hF000;
defparam \daddr~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N30
cycloneive_lcell_comb \daddr~32 (
// Equation(s):
// \daddr~32_combout  = (\nRST~input_o  & Selector0)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(Selector0),
	.cin(gnd),
	.combout(\daddr~32_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~32 .lut_mask = 16'hF000;
defparam \daddr~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N4
cycloneive_lcell_comb \daddr~33 (
// Equation(s):
// \daddr~33_combout  = (\nRST~input_o  & Selector1)

	.dataa(gnd),
	.datab(gnd),
	.datac(nRST),
	.datad(Selector1),
	.cin(gnd),
	.combout(\daddr~33_combout ),
	.cout());
// synopsys translate_off
defparam \daddr~33 .lut_mask = 16'hF000;
defparam \daddr~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N10
cycloneive_lcell_comb \instr~52 (
// Equation(s):
// \instr~52_combout  = (\nRST~input_o  & (!iwait & ((ramiframload_28) # (!always1))))

	.dataa(ramiframload_28),
	.datab(nRST),
	.datac(iwait),
	.datad(always1),
	.cin(gnd),
	.combout(\instr~52_combout ),
	.cout());
// synopsys translate_off
defparam \instr~52 .lut_mask = 16'h080C;
defparam \instr~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N30
cycloneive_lcell_comb \instr~53 (
// Equation(s):
// \instr~53_combout  = (\nRST~input_o  & (!iwait & ((ramiframload_27) # (!always1))))

	.dataa(nRST),
	.datab(ramiframload_27),
	.datac(iwait),
	.datad(always1),
	.cin(gnd),
	.combout(\instr~53_combout ),
	.cout());
// synopsys translate_off
defparam \instr~53 .lut_mask = 16'h080A;
defparam \instr~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N18
cycloneive_lcell_comb \instr~54 (
// Equation(s):
// \instr~54_combout  = (!iwait & (\nRST~input_o  & ((ramiframload_29) # (!always1))))

	.dataa(always1),
	.datab(ramiframload_29),
	.datac(iwait),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~54_combout ),
	.cout());
// synopsys translate_off
defparam \instr~54 .lut_mask = 16'h0D00;
defparam \instr~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N20
cycloneive_lcell_comb \instr~55 (
// Equation(s):
// \instr~55_combout  = (ramiframload_26 & (!iwait & (\nRST~input_o  & always1)))

	.dataa(ramiframload_26),
	.datab(iwait),
	.datac(nRST),
	.datad(always1),
	.cin(gnd),
	.combout(\instr~55_combout ),
	.cout());
// synopsys translate_off
defparam \instr~55 .lut_mask = 16'h2000;
defparam \instr~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N4
cycloneive_lcell_comb \instr~56 (
// Equation(s):
// \instr~56_combout  = (\nRST~input_o  & (always1 & (!iwait & ramiframload_30)))

	.dataa(nRST),
	.datab(always1),
	.datac(iwait),
	.datad(ramiframload_30),
	.cin(gnd),
	.combout(\instr~56_combout ),
	.cout());
// synopsys translate_off
defparam \instr~56 .lut_mask = 16'h0800;
defparam \instr~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N14
cycloneive_lcell_comb \instr~57 (
// Equation(s):
// \instr~57_combout  = (!iwait & (\nRST~input_o  & ((ramiframload_31) # (!always1))))

	.dataa(always1),
	.datab(ramiframload_31),
	.datac(iwait),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~57_combout ),
	.cout());
// synopsys translate_off
defparam \instr~57 .lut_mask = 16'h0D00;
defparam \instr~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N28
cycloneive_lcell_comb \instr~58 (
// Equation(s):
// \instr~58_combout  = (ramiframload_19 & (\nRST~input_o  & (!ruifdmemWEN & !ruifdmemREN)))

	.dataa(ramiframload_19),
	.datab(nRST),
	.datac(ruifdmemWEN),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(\instr~58_combout ),
	.cout());
// synopsys translate_off
defparam \instr~58 .lut_mask = 16'h0008;
defparam \instr~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N9
dffeas \instr[19] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~58_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[19]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[19] .is_wysiwyg = "true";
defparam \instr[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N20
cycloneive_lcell_comb \instr~59 (
// Equation(s):
// \instr~59_combout  = (ramiframload_18 & (!ruifdmemREN & (!ruifdmemWEN & \nRST~input_o )))

	.dataa(ramiframload_18),
	.datab(ruifdmemREN),
	.datac(ruifdmemWEN),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~59_combout ),
	.cout());
// synopsys translate_off
defparam \instr~59 .lut_mask = 16'h0200;
defparam \instr~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y32_N7
dffeas \instr[18] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~59_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[18]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[18] .is_wysiwyg = "true";
defparam \instr[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N20
cycloneive_lcell_comb \instr~60 (
// Equation(s):
// \instr~60_combout  = (ramiframload_16 & (!ruifdmemWEN & (\nRST~input_o  & !ruifdmemREN)))

	.dataa(ramiframload_16),
	.datab(ruifdmemWEN),
	.datac(nRST),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(\instr~60_combout ),
	.cout());
// synopsys translate_off
defparam \instr~60 .lut_mask = 16'h0020;
defparam \instr~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N1
dffeas \instr[16] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~60_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[16]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[16] .is_wysiwyg = "true";
defparam \instr[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N26
cycloneive_lcell_comb \instr~61 (
// Equation(s):
// \instr~61_combout  = (\nRST~input_o  & (!ruifdmemWEN & (ramiframload_17 & !ruifdmemREN)))

	.dataa(nRST),
	.datab(ruifdmemWEN),
	.datac(ramiframload_17),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(\instr~61_combout ),
	.cout());
// synopsys translate_off
defparam \instr~61 .lut_mask = 16'h0020;
defparam \instr~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y37_N5
dffeas \instr[17] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~61_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[17]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[17] .is_wysiwyg = "true";
defparam \instr[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N2
cycloneive_lcell_comb \instr~62 (
// Equation(s):
// \instr~62_combout  = (!ruifdmemREN & (ramiframload_20 & (!ruifdmemWEN & \nRST~input_o )))

	.dataa(ruifdmemREN),
	.datab(ramiframload_20),
	.datac(ruifdmemWEN),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~62_combout ),
	.cout());
// synopsys translate_off
defparam \instr~62 .lut_mask = 16'h0400;
defparam \instr~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y33_N21
dffeas \instr[20] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~62_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[20]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[20] .is_wysiwyg = "true";
defparam \instr[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N16
cycloneive_lcell_comb \instr~63 (
// Equation(s):
// \instr~63_combout  = (!ruifdmemREN & (\nRST~input_o  & (!ruifdmemWEN & ramiframload_3)))

	.dataa(ruifdmemREN),
	.datab(nRST),
	.datac(ruifdmemWEN),
	.datad(ramiframload_3),
	.cin(gnd),
	.combout(\instr~63_combout ),
	.cout());
// synopsys translate_off
defparam \instr~63 .lut_mask = 16'h0400;
defparam \instr~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N31
dffeas \instr[3] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~63_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[3]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[3] .is_wysiwyg = "true";
defparam \instr[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N20
cycloneive_lcell_comb \instr~64 (
// Equation(s):
// \instr~64_combout  = (!ruifdmemWEN & (ramiframload_4 & (!ruifdmemREN & \nRST~input_o )))

	.dataa(ruifdmemWEN),
	.datab(ramiframload_4),
	.datac(ruifdmemREN),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~64_combout ),
	.cout());
// synopsys translate_off
defparam \instr~64 .lut_mask = 16'h0400;
defparam \instr~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N1
dffeas \instr[4] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~64_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[4]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[4] .is_wysiwyg = "true";
defparam \instr[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N22
cycloneive_lcell_comb \instr~65 (
// Equation(s):
// \instr~65_combout  = (\nRST~input_o  & (!ruifdmemWEN & (ramiframload_0 & !ruifdmemREN)))

	.dataa(nRST),
	.datab(ruifdmemWEN),
	.datac(ramiframload_0),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(\instr~65_combout ),
	.cout());
// synopsys translate_off
defparam \instr~65 .lut_mask = 16'h0020;
defparam \instr~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y32_N17
dffeas \instr[0] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~65_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[0]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[0] .is_wysiwyg = "true";
defparam \instr[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N2
cycloneive_lcell_comb \instr~66 (
// Equation(s):
// \instr~66_combout  = (ramiframload_1 & (!ruifdmemWEN & (!ruifdmemREN & \nRST~input_o )))

	.dataa(ramiframload_1),
	.datab(ruifdmemWEN),
	.datac(ruifdmemREN),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~66_combout ),
	.cout());
// synopsys translate_off
defparam \instr~66 .lut_mask = 16'h0200;
defparam \instr~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N15
dffeas \instr[1] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~66_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[1]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[1] .is_wysiwyg = "true";
defparam \instr[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N18
cycloneive_lcell_comb \instr~67 (
// Equation(s):
// \instr~67_combout  = (ramiframload_2 & (!ruifdmemWEN & (\nRST~input_o  & !ruifdmemREN)))

	.dataa(ramiframload_2),
	.datab(ruifdmemWEN),
	.datac(nRST),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(\instr~67_combout ),
	.cout());
// synopsys translate_off
defparam \instr~67 .lut_mask = 16'h0020;
defparam \instr~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N15
dffeas \instr[2] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~67_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[2]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[2] .is_wysiwyg = "true";
defparam \instr[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N30
cycloneive_lcell_comb \instr~68 (
// Equation(s):
// \instr~68_combout  = (ramiframload_5 & (!ruifdmemWEN & (!ruifdmemREN & \nRST~input_o )))

	.dataa(ramiframload_5),
	.datab(ruifdmemWEN),
	.datac(ruifdmemREN),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~68_combout ),
	.cout());
// synopsys translate_off
defparam \instr~68 .lut_mask = 16'h0200;
defparam \instr~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y35_N19
dffeas \instr[5] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~68_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[5]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[5] .is_wysiwyg = "true";
defparam \instr[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N22
cycloneive_lcell_comb \instr~69 (
// Equation(s):
// \instr~69_combout  = (!ruifdmemREN & (\nRST~input_o  & (ramiframload_15 & !ruifdmemWEN)))

	.dataa(ruifdmemREN),
	.datab(nRST),
	.datac(ramiframload_15),
	.datad(ruifdmemWEN),
	.cin(gnd),
	.combout(\instr~69_combout ),
	.cout());
// synopsys translate_off
defparam \instr~69 .lut_mask = 16'h0040;
defparam \instr~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y35_N21
dffeas \instr[15] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~69_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[15]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[15] .is_wysiwyg = "true";
defparam \instr[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N26
cycloneive_lcell_comb \instr~70 (
// Equation(s):
// \instr~70_combout  = (!ruifdmemREN & (!ruifdmemWEN & (\nRST~input_o  & ramiframload_14)))

	.dataa(ruifdmemREN),
	.datab(ruifdmemWEN),
	.datac(nRST),
	.datad(ramiframload_14),
	.cin(gnd),
	.combout(\instr~70_combout ),
	.cout());
// synopsys translate_off
defparam \instr~70 .lut_mask = 16'h1000;
defparam \instr~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y35_N7
dffeas \instr[14] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~70_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[14]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[14] .is_wysiwyg = "true";
defparam \instr[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N8
cycloneive_lcell_comb \instr~71 (
// Equation(s):
// \instr~71_combout  = (!ruifdmemREN & (ramiframload_13 & (!ruifdmemWEN & \nRST~input_o )))

	.dataa(ruifdmemREN),
	.datab(ramiframload_13),
	.datac(ruifdmemWEN),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~71_combout ),
	.cout());
// synopsys translate_off
defparam \instr~71 .lut_mask = 16'h0400;
defparam \instr~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y32_N29
dffeas \instr[13] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~71_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[13]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[13] .is_wysiwyg = "true";
defparam \instr[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N22
cycloneive_lcell_comb \instr~72 (
// Equation(s):
// \instr~72_combout  = (!ruifdmemWEN & (!ruifdmemREN & (ramiframload_12 & \nRST~input_o )))

	.dataa(ruifdmemWEN),
	.datab(ruifdmemREN),
	.datac(ramiframload_12),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~72_combout ),
	.cout());
// synopsys translate_off
defparam \instr~72 .lut_mask = 16'h1000;
defparam \instr~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y33_N3
dffeas \instr[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~72_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[12]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[12] .is_wysiwyg = "true";
defparam \instr[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N0
cycloneive_lcell_comb \instr~73 (
// Equation(s):
// \instr~73_combout  = (\nRST~input_o  & (!ruifdmemWEN & (ramiframload_11 & !ruifdmemREN)))

	.dataa(nRST),
	.datab(ruifdmemWEN),
	.datac(ramiframload_11),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(\instr~73_combout ),
	.cout());
// synopsys translate_off
defparam \instr~73 .lut_mask = 16'h0020;
defparam \instr~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y33_N31
dffeas \instr[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~73_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[11]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[11] .is_wysiwyg = "true";
defparam \instr[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N10
cycloneive_lcell_comb \instr~74 (
// Equation(s):
// \instr~74_combout  = (\nRST~input_o  & (ramiframload_10 & (!ruifdmemWEN & !ruifdmemREN)))

	.dataa(nRST),
	.datab(ramiframload_10),
	.datac(ruifdmemWEN),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(\instr~74_combout ),
	.cout());
// synopsys translate_off
defparam \instr~74 .lut_mask = 16'h0008;
defparam \instr~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y35_N9
dffeas \instr[10] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~74_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[10]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[10] .is_wysiwyg = "true";
defparam \instr[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N4
cycloneive_lcell_comb \instr~75 (
// Equation(s):
// \instr~75_combout  = (ramiframload_9 & (!ruifdmemWEN & (\nRST~input_o  & !ruifdmemREN)))

	.dataa(ramiframload_9),
	.datab(ruifdmemWEN),
	.datac(nRST),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(\instr~75_combout ),
	.cout());
// synopsys translate_off
defparam \instr~75 .lut_mask = 16'h0020;
defparam \instr~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y35_N31
dffeas \instr[9] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~75_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[9]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[9] .is_wysiwyg = "true";
defparam \instr[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N8
cycloneive_lcell_comb \instr~76 (
// Equation(s):
// \instr~76_combout  = (ramiframload_8 & (!ruifdmemWEN & (!ruifdmemREN & \nRST~input_o )))

	.dataa(ramiframload_8),
	.datab(ruifdmemWEN),
	.datac(ruifdmemREN),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~76_combout ),
	.cout());
// synopsys translate_off
defparam \instr~76 .lut_mask = 16'h0200;
defparam \instr~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y33_N31
dffeas \instr[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~76_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[8]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[8] .is_wysiwyg = "true";
defparam \instr[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N26
cycloneive_lcell_comb \instr~77 (
// Equation(s):
// \instr~77_combout  = (!ruifdmemREN & (ramiframload_7 & (!ruifdmemWEN & \nRST~input_o )))

	.dataa(ruifdmemREN),
	.datab(ramiframload_7),
	.datac(ruifdmemWEN),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~77_combout ),
	.cout());
// synopsys translate_off
defparam \instr~77 .lut_mask = 16'h0400;
defparam \instr~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y33_N15
dffeas \instr[7] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~77_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[7]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[7] .is_wysiwyg = "true";
defparam \instr[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N28
cycloneive_lcell_comb \instr~78 (
// Equation(s):
// \instr~78_combout  = (!ruifdmemWEN & (\nRST~input_o  & (ramiframload_6 & !ruifdmemREN)))

	.dataa(ruifdmemWEN),
	.datab(nRST),
	.datac(ramiframload_6),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(\instr~78_combout ),
	.cout());
// synopsys translate_off
defparam \instr~78 .lut_mask = 16'h0040;
defparam \instr~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y35_N17
dffeas \instr[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~78_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[6]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[6] .is_wysiwyg = "true";
defparam \instr[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y35_N22
cycloneive_lcell_comb \instr~79 (
// Equation(s):
// \instr~79_combout  = (ramiframload_23 & (!ruifdmemWEN & (\nRST~input_o  & !ruifdmemREN)))

	.dataa(ramiframload_23),
	.datab(ruifdmemWEN),
	.datac(nRST),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(\instr~79_combout ),
	.cout());
// synopsys translate_off
defparam \instr~79 .lut_mask = 16'h0020;
defparam \instr~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N25
dffeas \instr[23] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~79_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[23]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[23] .is_wysiwyg = "true";
defparam \instr[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N26
cycloneive_lcell_comb \instr~80 (
// Equation(s):
// \instr~80_combout  = (\nRST~input_o  & (!ruifdmemWEN & (ramiframload_24 & !ruifdmemREN)))

	.dataa(nRST),
	.datab(ruifdmemWEN),
	.datac(ramiframload_24),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(\instr~80_combout ),
	.cout());
// synopsys translate_off
defparam \instr~80 .lut_mask = 16'h0020;
defparam \instr~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N13
dffeas \instr[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~80_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[24]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[24] .is_wysiwyg = "true";
defparam \instr[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N30
cycloneive_lcell_comb \instr~81 (
// Equation(s):
// \instr~81_combout  = (!ruifdmemREN & (ramiframload_21 & (!ruifdmemWEN & \nRST~input_o )))

	.dataa(ruifdmemREN),
	.datab(ramiframload_21),
	.datac(ruifdmemWEN),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~81_combout ),
	.cout());
// synopsys translate_off
defparam \instr~81 .lut_mask = 16'h0400;
defparam \instr~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N17
dffeas \instr[21] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~81_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[21]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[21] .is_wysiwyg = "true";
defparam \instr[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N30
cycloneive_lcell_comb \instr~82 (
// Equation(s):
// \instr~82_combout  = (ramiframload_22 & (\nRST~input_o  & (!ruifdmemWEN & !ruifdmemREN)))

	.dataa(ramiframload_22),
	.datab(nRST),
	.datac(ruifdmemWEN),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(\instr~82_combout ),
	.cout());
// synopsys translate_off
defparam \instr~82 .lut_mask = 16'h0008;
defparam \instr~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y35_N9
dffeas \instr[22] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~82_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[22]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[22] .is_wysiwyg = "true";
defparam \instr[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N12
cycloneive_lcell_comb \instr~83 (
// Equation(s):
// \instr~83_combout  = (ramiframload_25 & (!ruifdmemWEN & (!ruifdmemREN & \nRST~input_o )))

	.dataa(ramiframload_25),
	.datab(ruifdmemWEN),
	.datac(ruifdmemREN),
	.datad(nRST),
	.cin(gnd),
	.combout(\instr~83_combout ),
	.cout());
// synopsys translate_off
defparam \instr~83 .lut_mask = 16'h0200;
defparam \instr~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y36_N25
dffeas \instr[25] (
	.clk(CLK),
	.d(gnd),
	.asdata(\instr~83_combout ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\daddr[31]~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(instr[25]),
	.prn(vcc));
// synopsys translate_off
defparam \instr[25] .is_wysiwyg = "true";
defparam \instr[25] .power_up = "low";
// synopsys translate_on

endmodule

module datapath (
	pcifimemaddr_29,
	pcifimemaddr_28,
	pcifimemaddr_31,
	pcifimemaddr_30,
	pcifimemaddr_1,
	ruifdmemREN,
	ruifdmemWEN,
	pcifimemaddr_0,
	pcifimemaddr_3,
	pcifimemaddr_2,
	pcifimemaddr_5,
	pcifimemaddr_4,
	pcifimemaddr_7,
	pcifimemaddr_6,
	pcifimemaddr_9,
	pcifimemaddr_8,
	pcifimemaddr_11,
	pcifimemaddr_10,
	pcifimemaddr_13,
	pcifimemaddr_12,
	pcifimemaddr_15,
	pcifimemaddr_14,
	pcifimemaddr_17,
	pcifimemaddr_16,
	pcifimemaddr_19,
	pcifimemaddr_18,
	pcifimemaddr_21,
	pcifimemaddr_20,
	pcifimemaddr_23,
	pcifimemaddr_22,
	pcifimemaddr_25,
	pcifimemaddr_24,
	pcifimemaddr_27,
	pcifimemaddr_26,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	iwait,
	instr_28,
	instr_27,
	instr_29,
	instr_26,
	instr_30,
	dcifimemload_30,
	instr_31,
	dcifimemload_31,
	dcifimemload_19,
	dcifimemload_29,
	dcifimemload_28,
	dcifimemload_26,
	dcifimemload_27,
	dcifimemload_18,
	dcifimemload_16,
	dcifimemload_17,
	Mux63,
	Mux631,
	dcifimemload_20,
	cuifregT_4,
	dcifimemload_3,
	dcifimemload_4,
	dcifimemload_0,
	dcifimemload_1,
	dcifimemload_2,
	dcifimemload_5,
	dcifimemload_15,
	Mux32,
	Mux321,
	Mux33,
	Mux331,
	Mux34,
	Mux341,
	Mux35,
	Mux351,
	Mux36,
	Mux361,
	Mux37,
	Mux371,
	Mux38,
	Mux381,
	Mux39,
	Mux391,
	Mux40,
	Mux401,
	Mux41,
	Mux411,
	Mux42,
	Mux421,
	Mux43,
	Mux431,
	Mux58,
	Mux581,
	Mux44,
	Mux441,
	Mux45,
	Mux451,
	Mux46,
	Mux461,
	Mux47,
	Mux471,
	Mux48,
	Mux481,
	dcifimemload_14,
	Mux49,
	Mux491,
	dcifimemload_13,
	Mux50,
	Mux501,
	dcifimemload_12,
	Mux51,
	Mux511,
	dcifimemload_11,
	Mux52,
	Mux521,
	dcifimemload_10,
	Mux53,
	Mux531,
	dcifimemload_9,
	Mux54,
	Mux541,
	dcifimemload_8,
	Mux55,
	Mux551,
	dcifimemload_7,
	Mux56,
	Mux561,
	dcifimemload_6,
	Mux57,
	Mux571,
	dcifimemload_23,
	dcifimemload_24,
	dcifimemload_21,
	dcifimemload_22,
	dcifimemload_25,
	Mux62,
	Mux621,
	Mux61,
	Mux611,
	Mux60,
	Mux601,
	Mux59,
	Mux591,
	Mux31,
	Selector30,
	ShiftRight0,
	Selector31,
	Selector311,
	Selector28,
	dcifimemload_261,
	ShiftLeft0,
	Selector0,
	ShiftLeft01,
	Selector2,
	Selector29,
	Selector4,
	Selector5,
	ShiftLeft02,
	Selector3,
	ShiftLeft03,
	Selector1,
	Selector41,
	Selector10,
	Selector6,
	Selector7,
	Selector11,
	Selector24,
	Selector241,
	Selector25,
	Selector13,
	Selector12,
	Selector26,
	Selector27,
	Selector14,
	Selector15,
	Selector16,
	Selector17,
	Selector20,
	Selector21,
	Selector18,
	Selector19,
	Selector8,
	Selector81,
	Selector82,
	Selector9,
	Selector22,
	Selector23,
	ramiframload_261,
	ramiframload_271,
	ramiframload_281,
	ramiframload_291,
	ramiframload_301,
	ramiframload_311,
	dcifdhit,
	dcifimemload_262,
	CLK,
	nRST,
	dpifhalt,
	devpor,
	devclrn,
	devoe);
output 	pcifimemaddr_29;
output 	pcifimemaddr_28;
output 	pcifimemaddr_31;
output 	pcifimemaddr_30;
output 	pcifimemaddr_1;
output 	ruifdmemREN;
output 	ruifdmemWEN;
output 	pcifimemaddr_0;
output 	pcifimemaddr_3;
output 	pcifimemaddr_2;
output 	pcifimemaddr_5;
output 	pcifimemaddr_4;
output 	pcifimemaddr_7;
output 	pcifimemaddr_6;
output 	pcifimemaddr_9;
output 	pcifimemaddr_8;
output 	pcifimemaddr_11;
output 	pcifimemaddr_10;
output 	pcifimemaddr_13;
output 	pcifimemaddr_12;
output 	pcifimemaddr_15;
output 	pcifimemaddr_14;
output 	pcifimemaddr_17;
output 	pcifimemaddr_16;
output 	pcifimemaddr_19;
output 	pcifimemaddr_18;
output 	pcifimemaddr_21;
output 	pcifimemaddr_20;
output 	pcifimemaddr_23;
output 	pcifimemaddr_22;
output 	pcifimemaddr_25;
output 	pcifimemaddr_24;
output 	pcifimemaddr_27;
output 	pcifimemaddr_26;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
input 	iwait;
input 	instr_28;
input 	instr_27;
input 	instr_29;
input 	instr_26;
input 	instr_30;
input 	dcifimemload_30;
input 	instr_31;
input 	dcifimemload_31;
input 	dcifimemload_19;
input 	dcifimemload_29;
input 	dcifimemload_28;
input 	dcifimemload_26;
input 	dcifimemload_27;
input 	dcifimemload_18;
input 	dcifimemload_16;
input 	dcifimemload_17;
output 	Mux63;
output 	Mux631;
input 	dcifimemload_20;
output 	cuifregT_4;
input 	dcifimemload_3;
input 	dcifimemload_4;
input 	dcifimemload_0;
input 	dcifimemload_1;
input 	dcifimemload_2;
input 	dcifimemload_5;
input 	dcifimemload_15;
output 	Mux32;
output 	Mux321;
output 	Mux33;
output 	Mux331;
output 	Mux34;
output 	Mux341;
output 	Mux35;
output 	Mux351;
output 	Mux36;
output 	Mux361;
output 	Mux37;
output 	Mux371;
output 	Mux38;
output 	Mux381;
output 	Mux39;
output 	Mux391;
output 	Mux40;
output 	Mux401;
output 	Mux41;
output 	Mux411;
output 	Mux42;
output 	Mux421;
output 	Mux43;
output 	Mux431;
output 	Mux58;
output 	Mux581;
output 	Mux44;
output 	Mux441;
output 	Mux45;
output 	Mux451;
output 	Mux46;
output 	Mux461;
output 	Mux47;
output 	Mux471;
output 	Mux48;
output 	Mux481;
input 	dcifimemload_14;
output 	Mux49;
output 	Mux491;
input 	dcifimemload_13;
output 	Mux50;
output 	Mux501;
input 	dcifimemload_12;
output 	Mux51;
output 	Mux511;
input 	dcifimemload_11;
output 	Mux52;
output 	Mux521;
input 	dcifimemload_10;
output 	Mux53;
output 	Mux531;
input 	dcifimemload_9;
output 	Mux54;
output 	Mux541;
input 	dcifimemload_8;
output 	Mux55;
output 	Mux551;
input 	dcifimemload_7;
output 	Mux56;
output 	Mux561;
input 	dcifimemload_6;
output 	Mux57;
output 	Mux571;
input 	dcifimemload_23;
input 	dcifimemload_24;
input 	dcifimemload_21;
input 	dcifimemload_22;
input 	dcifimemload_25;
output 	Mux62;
output 	Mux621;
output 	Mux61;
output 	Mux611;
output 	Mux60;
output 	Mux601;
output 	Mux59;
output 	Mux591;
output 	Mux31;
output 	Selector30;
output 	ShiftRight0;
output 	Selector31;
output 	Selector311;
output 	Selector28;
input 	dcifimemload_261;
output 	ShiftLeft0;
output 	Selector0;
output 	ShiftLeft01;
output 	Selector2;
output 	Selector29;
output 	Selector4;
output 	Selector5;
output 	ShiftLeft02;
output 	Selector3;
output 	ShiftLeft03;
output 	Selector1;
output 	Selector41;
output 	Selector10;
output 	Selector6;
output 	Selector7;
output 	Selector11;
output 	Selector24;
output 	Selector241;
output 	Selector25;
output 	Selector13;
output 	Selector12;
output 	Selector26;
output 	Selector27;
output 	Selector14;
output 	Selector15;
output 	Selector16;
output 	Selector17;
output 	Selector20;
output 	Selector21;
output 	Selector18;
output 	Selector19;
output 	Selector8;
output 	Selector81;
output 	Selector82;
output 	Selector9;
output 	Selector22;
output 	Selector23;
input 	ramiframload_261;
input 	ramiframload_271;
input 	ramiframload_281;
input 	ramiframload_291;
input 	ramiframload_301;
input 	ramiframload_311;
input 	dcifdhit;
input 	dcifimemload_262;
input 	CLK;
input 	nRST;
output 	dpifhalt;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add0~1 ;
wire \Add0~0_combout ;
wire \Add0~3 ;
wire \Add0~2_combout ;
wire \Add0~5 ;
wire \Add0~4_combout ;
wire \Add0~7 ;
wire \Add0~6_combout ;
wire \Add0~9 ;
wire \Add0~8_combout ;
wire \Add0~11 ;
wire \Add0~10_combout ;
wire \Add0~13 ;
wire \Add0~12_combout ;
wire \Add0~15 ;
wire \Add0~14_combout ;
wire \Add0~17 ;
wire \Add0~16_combout ;
wire \Add0~19 ;
wire \Add0~18_combout ;
wire \Add0~21 ;
wire \Add0~20_combout ;
wire \Add0~23 ;
wire \Add0~22_combout ;
wire \Add0~25 ;
wire \Add0~24_combout ;
wire \Add0~27 ;
wire \Add0~26_combout ;
wire \Add0~29 ;
wire \Add0~28_combout ;
wire \Add0~31 ;
wire \Add0~30_combout ;
wire \Add0~33 ;
wire \Add0~32_combout ;
wire \Add0~35 ;
wire \Add0~34_combout ;
wire \Add0~37 ;
wire \Add0~36_combout ;
wire \Add0~39 ;
wire \Add0~38_combout ;
wire \Add0~41 ;
wire \Add0~40_combout ;
wire \Add0~43 ;
wire \Add0~42_combout ;
wire \Add0~45 ;
wire \Add0~44_combout ;
wire \Add0~47 ;
wire \Add0~46_combout ;
wire \Add0~49 ;
wire \Add0~48_combout ;
wire \Add0~51 ;
wire \Add0~50_combout ;
wire \Add0~53 ;
wire \Add0~52_combout ;
wire \Add0~55 ;
wire \Add0~54_combout ;
wire \Add0~57 ;
wire \Add0~56_combout ;
wire \Add0~58_combout ;
wire \cu_dut|Equal12~2_combout ;
wire \cu_dut|Equal2~4_combout ;
wire \cu_dut|Equal2~7_combout ;
wire \cu_dut|cuif.regT[0]~1_combout ;
wire \cu_dut|cuif.regT[3]~2_combout ;
wire \cu_dut|cuif.regT[2]~3_combout ;
wire \cu_dut|cuif.regT[0]~4_combout ;
wire \cu_dut|cuif.regT[1]~5_combout ;
wire \cu_dut|cuif.aluOp[3]~1_combout ;
wire \cu_dut|cuif.aluOp[3]~3_combout ;
wire \cu_dut|cuif.aluOp[2]~8_combout ;
wire \cu_dut|cuif.aluOp[1]~13_combout ;
wire \cu_dut|cuif.aluOp[0]~17_combout ;
wire \cu_dut|cuif.aluSrc[0]~0_combout ;
wire \WideOr0~0_combout ;
wire \Mux5~0_combout ;
wire \cu_dut|WideOr4~2_combout ;
wire \cu_dut|Equal2~8_combout ;
wire \cu_dut|Equal0~0_combout ;
wire \cu_dut|cuif.aluSrc[1]~1_combout ;
wire \Mux5~1_combout ;
wire \Mux5~2_combout ;
wire \Mux5~3_combout ;
wire \Mux5~4_combout ;
wire \Mux6~0_combout ;
wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \Mux8~0_combout ;
wire \Mux9~0_combout ;
wire \Mux10~0_combout ;
wire \Mux11~0_combout ;
wire \Mux12~0_combout ;
wire \Mux12~1_combout ;
wire \Mux13~0_combout ;
wire \Mux14~0_combout ;
wire \Mux14~1_combout ;
wire \Mux15~0_combout ;
wire \Mux15~1_combout ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \Mux36~0_combout ;
wire \Mux31~0_combout ;
wire \Mux36~1_combout ;
wire \Mux31~1_combout ;
wire \Mux17~0_combout ;
wire \Mux18~0_combout ;
wire \Mux19~0_combout ;
wire \Mux20~0_combout ;
wire \Mux20~1_combout ;
wire \Mux5~5_combout ;
wire \Mux21~0_combout ;
wire \Mux21~1_combout ;
wire \Mux22~0_combout ;
wire \Mux22~1_combout ;
wire \Mux23~0_combout ;
wire \Mux23~1_combout ;
wire \Mux24~0_combout ;
wire \Mux24~1_combout ;
wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \Mux26~0_combout ;
wire \Mux26~1_combout ;
wire \Mux27~0_combout ;
wire \Mux27~1_combout ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \Mux29~0_combout ;
wire \Mux29~1_combout ;
wire \Mux30~0_combout ;
wire \Mux30~1_combout ;
wire \cu_dut|cuif.regS[2]~0_combout ;
wire \cu_dut|cuif.regS[3]~1_combout ;
wire \cu_dut|cuif.regS[0]~2_combout ;
wire \cu_dut|cuif.regS[1]~3_combout ;
wire \cu_dut|cuif.regS[4]~4_combout ;
wire \rf_dut|Mux29~20_combout ;
wire \rf_dut|Mux30~20_combout ;
wire \Mux36~2_combout ;
wire \Mux32~2_combout ;
wire \Mux36~3_combout ;
wire \Mux36~4_combout ;
wire \Mux35~2_combout ;
wire \Mux35~3_combout ;
wire \Mux35~4_combout ;
wire \rf_dut|Mux27~20_combout ;
wire \rf_dut|Mux28~20_combout ;
wire \Mux34~2_combout ;
wire \Mux34~3_combout ;
wire \rf_dut|Mux23~20_combout ;
wire \rf_dut|Mux24~20_combout ;
wire \rf_dut|Mux25~20_combout ;
wire \rf_dut|Mux26~20_combout ;
wire \Mux33~2_combout ;
wire \Mux33~3_combout ;
wire \rf_dut|Mux15~20_combout ;
wire \rf_dut|Mux16~20_combout ;
wire \rf_dut|Mux17~20_combout ;
wire \rf_dut|Mux18~20_combout ;
wire \rf_dut|Mux19~20_combout ;
wire \rf_dut|Mux20~20_combout ;
wire \rf_dut|Mux21~20_combout ;
wire \rf_dut|Mux22~20_combout ;
wire \Mux32~3_combout ;
wire \Mux32~4_combout ;
wire \rf_dut|Mux0~20_combout ;
wire \rf_dut|Mux2~20_combout ;
wire \rf_dut|Mux1~20_combout ;
wire \rf_dut|Mux3~20_combout ;
wire \rf_dut|Mux4~20_combout ;
wire \rf_dut|Mux5~20_combout ;
wire \rf_dut|Mux6~20_combout ;
wire \rf_dut|Mux7~20_combout ;
wire \rf_dut|Mux8~20_combout ;
wire \rf_dut|Mux9~20_combout ;
wire \rf_dut|Mux10~20_combout ;
wire \rf_dut|Mux11~20_combout ;
wire \rf_dut|Mux12~20_combout ;
wire \rf_dut|Mux13~20_combout ;
wire \rf_dut|Mux14~20_combout ;
wire \cu_dut|cuif.JmpSel[1]~1_combout ;
wire \cu_dut|cuif.JmpSel[0]~2_combout ;
wire \Mux5~6_combout ;
wire \Mux6~1_combout ;
wire \Mux8~1_combout ;
wire \Mux9~1_combout ;
wire \Mux10~1_combout ;
wire \Mux11~1_combout ;
wire \Mux13~1_combout ;
wire \Mux17~1_combout ;
wire \Mux18~1_combout ;
wire \Mux19~1_combout ;
wire \pc_dut|Equal0~0_combout ;
wire \alu_dut|Selector7~8_combout ;
wire \alu_dut|Selector24~9_combout ;
wire \alu_dut|Selector25~7_combout ;
wire \alu_dut|Selector26~7_combout ;
wire \alu_dut|Selector27~8_combout ;
wire \alu_dut|Equal10~6_combout ;
wire \alu_dut|Equal10~7_combout ;
wire \alu_dut|Selector31~9_combout ;
wire \alu_dut|Equal10~9_combout ;
wire \cu_dut|cuif.MemtoReg[1]~2_combout ;
wire \Mux68~0_combout ;
wire \cu_dut|cuif.MemtoReg[0]~4_combout ;
wire \Mux68~1_combout ;
wire \Mux0~0_combout ;
wire \Mux4~0_combout ;
wire \cu_dut|cuif.RegDst[0]~0_combout ;
wire \Mux4~1_combout ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \Mux0~1_combout ;
wire \Mux0~2_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \WEN~2_combout ;
wire \WEN~3_combout ;
wire \WEN~4_combout ;
wire \WEN~5_combout ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \Mux37~0_combout ;
wire \Mux37~1_combout ;
wire \Mux38~0_combout ;
wire \Mux38~1_combout ;
wire \Mux39~0_combout ;
wire \Mux39~1_combout ;
wire \Mux40~0_combout ;
wire \Mux40~1_combout ;
wire \Mux41~0_combout ;
wire \Mux41~1_combout ;
wire \Mux42~0_combout ;
wire \Mux42~1_combout ;
wire \Mux43~0_combout ;
wire \Mux43~1_combout ;
wire \Mux44~0_combout ;
wire \Mux44~1_combout ;
wire \alu_dut|Selector8~11_combout ;
wire \Mux45~0_combout ;
wire \Mux45~1_combout ;
wire \Mux46~0_combout ;
wire \Mux46~1_combout ;
wire \Mux47~0_combout ;
wire \Mux47~1_combout ;
wire \Mux48~0_combout ;
wire \Mux48~1_combout ;
wire \Mux63~0_combout ;
wire \Mux63~1_combout ;
wire \Mux49~0_combout ;
wire \Mux49~1_combout ;
wire \Mux50~0_combout ;
wire \Mux50~1_combout ;
wire \Mux51~0_combout ;
wire \Mux51~1_combout ;
wire \Mux52~0_combout ;
wire \Mux52~1_combout ;
wire \Mux53~0_combout ;
wire \Mux53~1_combout ;
wire \Mux54~0_combout ;
wire \Mux54~1_combout ;
wire \Mux55~0_combout ;
wire \Mux55~1_combout ;
wire \Mux56~0_combout ;
wire \Mux56~1_combout ;
wire \Mux57~0_combout ;
wire \Mux57~1_combout ;
wire \Mux58~0_combout ;
wire \Mux58~1_combout ;
wire \Mux59~0_combout ;
wire \Mux59~1_combout ;
wire \Mux60~0_combout ;
wire \Mux60~1_combout ;
wire \Mux61~0_combout ;
wire \Mux61~1_combout ;
wire \Mux62~0_combout ;
wire \Mux62~1_combout ;
wire \Mux66~0_combout ;
wire \Mux66~1_combout ;
wire \Mux67~0_combout ;
wire \Mux67~1_combout ;
wire \Mux64~0_combout ;
wire \Mux64~1_combout ;
wire \Mux65~0_combout ;
wire \Mux65~1_combout ;
wire \Mux35~5_combout ;
wire \Mux34~4_combout ;
wire \Mux33~4_combout ;
wire \Mux32~5_combout ;
wire \cu_dut|Equal2~9_combout ;
wire \WEN~6_combout ;
wire \dpif.halt~_Duplicate_1feeder_combout ;
wire \dpif.halt~_Duplicate_1_q ;
wire \dpif.halt~0_combout ;


register_file rf_dut(
	.always1(always1),
	.cuifregT_3(\cu_dut|cuif.regT[3]~2_combout ),
	.cuifregT_2(\cu_dut|cuif.regT[2]~3_combout ),
	.cuifregT_0(\cu_dut|cuif.regT[0]~4_combout ),
	.cuifregT_1(\cu_dut|cuif.regT[1]~5_combout ),
	.Mux63(Mux63),
	.Mux631(Mux631),
	.Mux32(Mux32),
	.Mux321(Mux321),
	.Mux33(Mux33),
	.Mux331(Mux331),
	.Mux34(Mux34),
	.Mux341(Mux341),
	.Mux35(Mux35),
	.Mux351(Mux351),
	.Mux36(Mux36),
	.Mux361(Mux361),
	.Mux37(Mux37),
	.Mux371(Mux371),
	.Mux38(Mux38),
	.Mux381(Mux381),
	.Mux39(Mux39),
	.Mux391(Mux391),
	.Mux40(Mux40),
	.Mux401(Mux401),
	.Mux41(Mux41),
	.Mux411(Mux411),
	.Mux42(Mux42),
	.Mux421(Mux421),
	.Mux43(Mux43),
	.Mux431(Mux431),
	.Mux58(Mux58),
	.Mux581(Mux581),
	.Mux44(Mux44),
	.Mux441(Mux441),
	.Mux45(Mux45),
	.Mux451(Mux451),
	.Mux46(Mux46),
	.Mux461(Mux461),
	.Mux47(Mux47),
	.Mux471(Mux471),
	.Mux48(Mux48),
	.Mux481(Mux481),
	.Mux49(Mux49),
	.Mux491(Mux491),
	.Mux50(Mux50),
	.Mux501(Mux501),
	.Mux51(Mux51),
	.Mux511(Mux511),
	.Mux52(Mux52),
	.Mux521(Mux521),
	.Mux53(Mux53),
	.Mux531(Mux531),
	.Mux54(Mux54),
	.Mux541(Mux541),
	.Mux55(Mux55),
	.Mux551(Mux551),
	.Mux56(Mux56),
	.Mux561(Mux561),
	.Mux57(Mux57),
	.Mux571(Mux571),
	.cuifregS_2(\cu_dut|cuif.regS[2]~0_combout ),
	.cuifregS_3(\cu_dut|cuif.regS[3]~1_combout ),
	.cuifregS_0(\cu_dut|cuif.regS[0]~2_combout ),
	.cuifregS_1(\cu_dut|cuif.regS[1]~3_combout ),
	.cuifregS_4(\cu_dut|cuif.regS[4]~4_combout ),
	.Mux29(\rf_dut|Mux29~20_combout ),
	.Mux30(\rf_dut|Mux30~20_combout ),
	.Mux62(Mux62),
	.Mux621(Mux621),
	.Mux27(\rf_dut|Mux27~20_combout ),
	.Mux28(\rf_dut|Mux28~20_combout ),
	.Mux61(Mux61),
	.Mux611(Mux611),
	.Mux23(\rf_dut|Mux23~20_combout ),
	.Mux24(\rf_dut|Mux24~20_combout ),
	.Mux25(\rf_dut|Mux25~20_combout ),
	.Mux26(\rf_dut|Mux26~20_combout ),
	.Mux60(Mux60),
	.Mux601(Mux601),
	.Mux15(\rf_dut|Mux15~20_combout ),
	.Mux16(\rf_dut|Mux16~20_combout ),
	.Mux17(\rf_dut|Mux17~20_combout ),
	.Mux18(\rf_dut|Mux18~20_combout ),
	.Mux19(\rf_dut|Mux19~20_combout ),
	.Mux20(\rf_dut|Mux20~20_combout ),
	.Mux21(\rf_dut|Mux21~20_combout ),
	.Mux22(\rf_dut|Mux22~20_combout ),
	.Mux59(Mux59),
	.Mux591(Mux591),
	.Mux0(\rf_dut|Mux0~20_combout ),
	.Mux2(\rf_dut|Mux2~20_combout ),
	.Mux1(\rf_dut|Mux1~20_combout ),
	.Mux3(\rf_dut|Mux3~20_combout ),
	.Mux4(\rf_dut|Mux4~20_combout ),
	.Mux5(\rf_dut|Mux5~20_combout ),
	.Mux6(\rf_dut|Mux6~20_combout ),
	.Mux7(\rf_dut|Mux7~20_combout ),
	.Mux8(\rf_dut|Mux8~20_combout ),
	.Mux9(\rf_dut|Mux9~20_combout ),
	.Mux10(\rf_dut|Mux10~20_combout ),
	.Mux11(\rf_dut|Mux11~20_combout ),
	.Mux12(\rf_dut|Mux12~20_combout ),
	.Mux13(\rf_dut|Mux13~20_combout ),
	.Mux14(\rf_dut|Mux14~20_combout ),
	.Mux31(Mux31),
	.Mux68(\Mux68~1_combout ),
	.Mux410(\Mux4~1_combout ),
	.Mux210(\Mux2~1_combout ),
	.Mux01(\Mux0~2_combout ),
	.Mux110(\Mux1~1_combout ),
	.WEN(\WEN~5_combout ),
	.Mux310(\Mux3~1_combout ),
	.Mux372(\Mux37~1_combout ),
	.Mux382(\Mux38~1_combout ),
	.Mux392(\Mux39~1_combout ),
	.Mux402(\Mux40~1_combout ),
	.Mux412(\Mux41~1_combout ),
	.Mux422(\Mux42~1_combout ),
	.Mux432(\Mux43~1_combout ),
	.Mux442(\Mux44~1_combout ),
	.Mux452(\Mux45~1_combout ),
	.Mux462(\Mux46~1_combout ),
	.Mux472(\Mux47~1_combout ),
	.Mux482(\Mux48~1_combout ),
	.Mux632(\Mux63~1_combout ),
	.Mux492(\Mux49~1_combout ),
	.Mux502(\Mux50~1_combout ),
	.Mux512(\Mux51~1_combout ),
	.Mux522(\Mux52~1_combout ),
	.Mux532(\Mux53~1_combout ),
	.Mux542(\Mux54~1_combout ),
	.Mux552(\Mux55~1_combout ),
	.Mux562(\Mux56~1_combout ),
	.Mux572(\Mux57~1_combout ),
	.Mux582(\Mux58~1_combout ),
	.Mux592(\Mux59~1_combout ),
	.Mux602(\Mux60~1_combout ),
	.Mux612(\Mux61~1_combout ),
	.Mux622(\Mux62~1_combout ),
	.Mux66(\Mux66~1_combout ),
	.Mux67(\Mux67~1_combout ),
	.Mux64(\Mux64~1_combout ),
	.Mux65(\Mux65~1_combout ),
	.clk(CLK),
	.n_rst(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

alu alu_dut(
	.cuifaluOp_3(\cu_dut|cuif.aluOp[3]~3_combout ),
	.cuifaluOp_2(\cu_dut|cuif.aluOp[2]~8_combout ),
	.cuifaluOp_1(\cu_dut|cuif.aluOp[1]~13_combout ),
	.cuifaluOp_0(\cu_dut|cuif.aluOp[0]~17_combout ),
	.Mux5(\Mux5~1_combout ),
	.Mux51(\Mux5~4_combout ),
	.Mux6(\Mux6~0_combout ),
	.Mux7(\Mux7~1_combout ),
	.Mux8(\Mux8~0_combout ),
	.Mux9(\Mux9~0_combout ),
	.Mux10(\Mux10~0_combout ),
	.Mux11(\Mux11~0_combout ),
	.Mux12(\Mux12~1_combout ),
	.Mux13(\Mux13~0_combout ),
	.Mux14(\Mux14~1_combout ),
	.Mux15(\Mux15~0_combout ),
	.Mux151(\Mux15~1_combout ),
	.Mux16(\Mux16~1_combout ),
	.Mux31(\Mux31~1_combout ),
	.Mux17(\Mux17~0_combout ),
	.Mux18(\Mux18~0_combout ),
	.Mux19(\Mux19~0_combout ),
	.Mux20(\Mux20~1_combout ),
	.Mux21(\Mux21~1_combout ),
	.Mux22(\Mux22~1_combout ),
	.Mux23(\Mux23~1_combout ),
	.Mux24(\Mux24~1_combout ),
	.Mux25(\Mux25~1_combout ),
	.Mux26(\Mux26~1_combout ),
	.Mux27(\Mux27~1_combout ),
	.Mux28(\Mux28~1_combout ),
	.Mux29(\Mux29~1_combout ),
	.Mux30(\Mux30~1_combout ),
	.Mux291(\rf_dut|Mux29~20_combout ),
	.Mux301(\rf_dut|Mux30~20_combout ),
	.Mux36(\Mux36~4_combout ),
	.Mux35(\Mux35~2_combout ),
	.Mux351(\Mux35~3_combout ),
	.Mux352(\Mux35~4_combout ),
	.Mux271(\rf_dut|Mux27~20_combout ),
	.Mux281(\rf_dut|Mux28~20_combout ),
	.Mux34(\Mux34~3_combout ),
	.Mux231(\rf_dut|Mux23~20_combout ),
	.Mux241(\rf_dut|Mux24~20_combout ),
	.Mux251(\rf_dut|Mux25~20_combout ),
	.Mux261(\rf_dut|Mux26~20_combout ),
	.Mux33(\Mux33~3_combout ),
	.Mux152(\rf_dut|Mux15~20_combout ),
	.Mux161(\rf_dut|Mux16~20_combout ),
	.Mux171(\rf_dut|Mux17~20_combout ),
	.Mux181(\rf_dut|Mux18~20_combout ),
	.Mux191(\rf_dut|Mux19~20_combout ),
	.Mux201(\rf_dut|Mux20~20_combout ),
	.Mux211(\rf_dut|Mux21~20_combout ),
	.Mux221(\rf_dut|Mux22~20_combout ),
	.Mux32(\Mux32~4_combout ),
	.Mux0(\rf_dut|Mux0~20_combout ),
	.Mux2(\rf_dut|Mux2~20_combout ),
	.Mux1(\rf_dut|Mux1~20_combout ),
	.Mux3(\rf_dut|Mux3~20_combout ),
	.Mux4(\rf_dut|Mux4~20_combout ),
	.Mux52(\rf_dut|Mux5~20_combout ),
	.Mux61(\rf_dut|Mux6~20_combout ),
	.Mux71(\rf_dut|Mux7~20_combout ),
	.Mux81(\rf_dut|Mux8~20_combout ),
	.Mux91(\rf_dut|Mux9~20_combout ),
	.Mux101(\rf_dut|Mux10~20_combout ),
	.Mux111(\rf_dut|Mux11~20_combout ),
	.Mux121(\rf_dut|Mux12~20_combout ),
	.Mux131(\rf_dut|Mux13~20_combout ),
	.Mux141(\rf_dut|Mux14~20_combout ),
	.Mux311(Mux31),
	.Selector30(Selector30),
	.ShiftRight0(ShiftRight0),
	.Mux53(\Mux5~6_combout ),
	.Mux62(\Mux6~1_combout ),
	.Mux82(\Mux8~1_combout ),
	.Mux92(\Mux9~1_combout ),
	.Mux102(\Mux10~1_combout ),
	.Mux112(\Mux11~1_combout ),
	.Mux132(\Mux13~1_combout ),
	.Mux172(\Mux17~1_combout ),
	.Mux182(\Mux18~1_combout ),
	.Mux192(\Mux19~1_combout ),
	.Selector31(Selector31),
	.Selector311(Selector311),
	.Selector28(Selector28),
	.ShiftLeft0(ShiftLeft0),
	.Selector0(Selector0),
	.ShiftLeft01(ShiftLeft01),
	.Selector2(Selector2),
	.Selector29(Selector29),
	.Selector4(Selector4),
	.Selector5(Selector5),
	.ShiftLeft02(ShiftLeft02),
	.Selector3(Selector3),
	.ShiftLeft03(ShiftLeft03),
	.Selector1(Selector1),
	.Selector41(Selector41),
	.Selector10(Selector10),
	.Selector6(Selector6),
	.Selector7(Selector7),
	.Selector71(\alu_dut|Selector7~8_combout ),
	.Selector11(Selector11),
	.Selector24(Selector24),
	.Selector241(Selector241),
	.Selector242(\alu_dut|Selector24~9_combout ),
	.Selector25(Selector25),
	.Selector251(\alu_dut|Selector25~7_combout ),
	.Selector13(Selector13),
	.Selector12(Selector12),
	.Selector26(Selector26),
	.Selector261(\alu_dut|Selector26~7_combout ),
	.Selector27(Selector27),
	.Selector271(\alu_dut|Selector27~8_combout ),
	.Equal10(\alu_dut|Equal10~6_combout ),
	.Selector14(Selector14),
	.Selector15(Selector15),
	.Selector16(Selector16),
	.Selector17(Selector17),
	.Equal101(\alu_dut|Equal10~7_combout ),
	.Selector20(Selector20),
	.Selector21(Selector21),
	.Selector18(Selector18),
	.Selector19(Selector19),
	.Selector8(Selector8),
	.Selector81(Selector81),
	.Selector82(Selector82),
	.Selector9(Selector9),
	.Selector312(\alu_dut|Selector31~9_combout ),
	.Selector22(Selector22),
	.Selector23(Selector23),
	.Equal102(\alu_dut|Equal10~9_combout ),
	.Selector83(\alu_dut|Selector8~11_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

pc_logic pc_dut(
	.pcifimemaddr_29(pcifimemaddr_29),
	.pcifimemaddr_28(pcifimemaddr_28),
	.pcifimemaddr_31(pcifimemaddr_31),
	.pcifimemaddr_30(pcifimemaddr_30),
	.dpifhalt(\dpif.halt~_Duplicate_1_q ),
	.pcifimemaddr_1(pcifimemaddr_1),
	.ruifdmemREN(ruifdmemREN),
	.ruifdmemWEN(ruifdmemWEN),
	.pcifimemaddr_0(pcifimemaddr_0),
	.pcifimemaddr_3(pcifimemaddr_3),
	.pcifimemaddr_2(pcifimemaddr_2),
	.pcifimemaddr_5(pcifimemaddr_5),
	.pcifimemaddr_4(pcifimemaddr_4),
	.pcifimemaddr_7(pcifimemaddr_7),
	.pcifimemaddr_6(pcifimemaddr_6),
	.pcifimemaddr_9(pcifimemaddr_9),
	.pcifimemaddr_8(pcifimemaddr_8),
	.pcifimemaddr_11(pcifimemaddr_11),
	.pcifimemaddr_10(pcifimemaddr_10),
	.pcifimemaddr_13(pcifimemaddr_13),
	.pcifimemaddr_12(pcifimemaddr_12),
	.pcifimemaddr_15(pcifimemaddr_15),
	.pcifimemaddr_14(pcifimemaddr_14),
	.pcifimemaddr_17(pcifimemaddr_17),
	.pcifimemaddr_16(pcifimemaddr_16),
	.pcifimemaddr_19(pcifimemaddr_19),
	.pcifimemaddr_18(pcifimemaddr_18),
	.pcifimemaddr_21(pcifimemaddr_21),
	.pcifimemaddr_20(pcifimemaddr_20),
	.pcifimemaddr_23(pcifimemaddr_23),
	.pcifimemaddr_22(pcifimemaddr_22),
	.pcifimemaddr_25(pcifimemaddr_25),
	.pcifimemaddr_24(pcifimemaddr_24),
	.pcifimemaddr_27(pcifimemaddr_27),
	.pcifimemaddr_26(pcifimemaddr_26),
	.always1(always1),
	.dcifimemload_19(dcifimemload_19),
	.dcifimemload_28(dcifimemload_28),
	.dcifimemload_27(dcifimemload_27),
	.dcifimemload_18(dcifimemload_18),
	.dcifimemload_16(dcifimemload_16),
	.dcifimemload_17(dcifimemload_17),
	.dcifimemload_20(dcifimemload_20),
	.dcifimemload_3(dcifimemload_3),
	.dcifimemload_4(dcifimemload_4),
	.dcifimemload_0(dcifimemload_0),
	.dcifimemload_1(dcifimemload_1),
	.dcifimemload_2(dcifimemload_2),
	.dcifimemload_5(dcifimemload_5),
	.dcifimemload_15(dcifimemload_15),
	.Equal2(\cu_dut|Equal2~8_combout ),
	.dcifimemload_14(dcifimemload_14),
	.dcifimemload_13(dcifimemload_13),
	.dcifimemload_12(dcifimemload_12),
	.dcifimemload_11(dcifimemload_11),
	.dcifimemload_10(dcifimemload_10),
	.dcifimemload_9(dcifimemload_9),
	.dcifimemload_8(dcifimemload_8),
	.dcifimemload_7(dcifimemload_7),
	.dcifimemload_6(dcifimemload_6),
	.dcifimemload_23(dcifimemload_23),
	.dcifimemload_24(dcifimemload_24),
	.dcifimemload_21(dcifimemload_21),
	.dcifimemload_22(dcifimemload_22),
	.dcifimemload_25(dcifimemload_25),
	.Mux29(\rf_dut|Mux29~20_combout ),
	.Mux30(\rf_dut|Mux30~20_combout ),
	.Mux27(\rf_dut|Mux27~20_combout ),
	.Mux28(\rf_dut|Mux28~20_combout ),
	.Mux23(\rf_dut|Mux23~20_combout ),
	.Mux24(\rf_dut|Mux24~20_combout ),
	.Mux25(\rf_dut|Mux25~20_combout ),
	.Mux26(\rf_dut|Mux26~20_combout ),
	.Mux15(\rf_dut|Mux15~20_combout ),
	.Mux16(\rf_dut|Mux16~20_combout ),
	.Mux17(\rf_dut|Mux17~20_combout ),
	.Mux18(\rf_dut|Mux18~20_combout ),
	.Mux19(\rf_dut|Mux19~20_combout ),
	.Mux20(\rf_dut|Mux20~20_combout ),
	.Mux21(\rf_dut|Mux21~20_combout ),
	.Mux22(\rf_dut|Mux22~20_combout ),
	.Mux0(\rf_dut|Mux0~20_combout ),
	.Mux2(\rf_dut|Mux2~20_combout ),
	.Mux1(\rf_dut|Mux1~20_combout ),
	.Mux3(\rf_dut|Mux3~20_combout ),
	.Mux4(\rf_dut|Mux4~20_combout ),
	.Mux5(\rf_dut|Mux5~20_combout ),
	.Mux6(\rf_dut|Mux6~20_combout ),
	.Mux7(\rf_dut|Mux7~20_combout ),
	.Mux8(\rf_dut|Mux8~20_combout ),
	.Mux9(\rf_dut|Mux9~20_combout ),
	.Mux10(\rf_dut|Mux10~20_combout ),
	.Mux11(\rf_dut|Mux11~20_combout ),
	.Mux12(\rf_dut|Mux12~20_combout ),
	.Mux13(\rf_dut|Mux13~20_combout ),
	.Mux14(\rf_dut|Mux14~20_combout ),
	.Mux31(Mux31),
	.cuifJmpSel_1(\cu_dut|cuif.JmpSel[1]~1_combout ),
	.cuifJmpSel_0(\cu_dut|cuif.JmpSel[0]~2_combout ),
	.Equal0(\pc_dut|Equal0~0_combout ),
	.dcifimemload_26(dcifimemload_261),
	.Equal10(\alu_dut|Equal10~6_combout ),
	.Equal101(\alu_dut|Equal10~7_combout ),
	.Selector20(Selector20),
	.Selector21(Selector21),
	.Selector18(Selector18),
	.Selector19(Selector19),
	.Equal102(\alu_dut|Equal10~9_combout ),
	.dcifimemload_261(dcifimemload_262),
	.CPUCLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

control_unit cu_dut(
	.always1(always1),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.iwait(iwait),
	.instr_28(instr_28),
	.instr_27(instr_27),
	.instr_29(instr_29),
	.instr_26(instr_26),
	.Equal12(\cu_dut|Equal12~2_combout ),
	.instr_30(instr_30),
	.dcifimemload_30(dcifimemload_30),
	.instr_31(instr_31),
	.dcifimemload_31(dcifimemload_31),
	.dcifimemload_19(dcifimemload_19),
	.dcifimemload_29(dcifimemload_29),
	.dcifimemload_28(dcifimemload_28),
	.dcifimemload_26(dcifimemload_26),
	.dcifimemload_27(dcifimemload_27),
	.Equal2(\cu_dut|Equal2~4_combout ),
	.Equal21(\cu_dut|Equal2~7_combout ),
	.cuifregT_0(\cu_dut|cuif.regT[0]~1_combout ),
	.cuifregT_3(\cu_dut|cuif.regT[3]~2_combout ),
	.dcifimemload_18(dcifimemload_18),
	.cuifregT_2(\cu_dut|cuif.regT[2]~3_combout ),
	.dcifimemload_16(dcifimemload_16),
	.cuifregT_01(\cu_dut|cuif.regT[0]~4_combout ),
	.dcifimemload_17(dcifimemload_17),
	.cuifregT_1(\cu_dut|cuif.regT[1]~5_combout ),
	.dcifimemload_20(dcifimemload_20),
	.cuifregT_4(cuifregT_4),
	.dcifimemload_3(dcifimemload_3),
	.dcifimemload_4(dcifimemload_4),
	.cuifaluOp_3(\cu_dut|cuif.aluOp[3]~1_combout ),
	.dcifimemload_0(dcifimemload_0),
	.dcifimemload_1(dcifimemload_1),
	.dcifimemload_2(dcifimemload_2),
	.dcifimemload_5(dcifimemload_5),
	.cuifaluOp_31(\cu_dut|cuif.aluOp[3]~3_combout ),
	.cuifaluOp_2(\cu_dut|cuif.aluOp[2]~8_combout ),
	.cuifaluOp_1(\cu_dut|cuif.aluOp[1]~13_combout ),
	.cuifaluOp_0(\cu_dut|cuif.aluOp[0]~17_combout ),
	.cuifaluSrc_0(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.WideOr4(\cu_dut|WideOr4~2_combout ),
	.Equal22(\cu_dut|Equal2~8_combout ),
	.Equal0(\cu_dut|Equal0~0_combout ),
	.cuifaluSrc_1(\cu_dut|cuif.aluSrc[1]~1_combout ),
	.dcifimemload_23(dcifimemload_23),
	.cuifregS_2(\cu_dut|cuif.regS[2]~0_combout ),
	.dcifimemload_24(dcifimemload_24),
	.cuifregS_3(\cu_dut|cuif.regS[3]~1_combout ),
	.dcifimemload_21(dcifimemload_21),
	.cuifregS_0(\cu_dut|cuif.regS[0]~2_combout ),
	.dcifimemload_22(dcifimemload_22),
	.cuifregS_1(\cu_dut|cuif.regS[1]~3_combout ),
	.dcifimemload_25(dcifimemload_25),
	.cuifregS_4(\cu_dut|cuif.regS[4]~4_combout ),
	.cuifJmpSel_1(\cu_dut|cuif.JmpSel[1]~1_combout ),
	.cuifJmpSel_0(\cu_dut|cuif.JmpSel[0]~2_combout ),
	.Equal01(\pc_dut|Equal0~0_combout ),
	.cuifMemtoReg_1(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.cuifMemtoReg_0(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.cuifRegDst_0(\cu_dut|cuif.RegDst[0]~0_combout ),
	.Equal23(\cu_dut|Equal2~9_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

request_unit ru_dut(
	.ruifdmemREN(ruifdmemREN),
	.ruifdmemWEN(ruifdmemWEN),
	.always1(always1),
	.dcifimemload_30(dcifimemload_30),
	.dcifimemload_31(dcifimemload_31),
	.dcifimemload_29(dcifimemload_29),
	.Equal2(\cu_dut|Equal2~7_combout ),
	.dcifdhit(dcifdhit),
	.CPUCLK(CLK),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X50_Y39_N2
cycloneive_lcell_comb \Add0~0 (
// Equation(s):
// \Add0~0_combout  = pcifimemaddr_2 $ (VCC)
// \Add0~1  = CARRY(pcifimemaddr_2)

	.dataa(pcifimemaddr_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
// synopsys translate_off
defparam \Add0~0 .lut_mask = 16'h55AA;
defparam \Add0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N4
cycloneive_lcell_comb \Add0~2 (
// Equation(s):
// \Add0~2_combout  = (pcifimemaddr_3 & (!\Add0~1 )) # (!pcifimemaddr_3 & ((\Add0~1 ) # (GND)))
// \Add0~3  = CARRY((!\Add0~1 ) # (!pcifimemaddr_3))

	.dataa(gnd),
	.datab(pcifimemaddr_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
// synopsys translate_off
defparam \Add0~2 .lut_mask = 16'h3C3F;
defparam \Add0~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N6
cycloneive_lcell_comb \Add0~4 (
// Equation(s):
// \Add0~4_combout  = (pcifimemaddr_4 & (\Add0~3  $ (GND))) # (!pcifimemaddr_4 & (!\Add0~3  & VCC))
// \Add0~5  = CARRY((pcifimemaddr_4 & !\Add0~3 ))

	.dataa(pcifimemaddr_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
// synopsys translate_off
defparam \Add0~4 .lut_mask = 16'hA50A;
defparam \Add0~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N8
cycloneive_lcell_comb \Add0~6 (
// Equation(s):
// \Add0~6_combout  = (pcifimemaddr_5 & (!\Add0~5 )) # (!pcifimemaddr_5 & ((\Add0~5 ) # (GND)))
// \Add0~7  = CARRY((!\Add0~5 ) # (!pcifimemaddr_5))

	.dataa(gnd),
	.datab(pcifimemaddr_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
// synopsys translate_off
defparam \Add0~6 .lut_mask = 16'h3C3F;
defparam \Add0~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N10
cycloneive_lcell_comb \Add0~8 (
// Equation(s):
// \Add0~8_combout  = (pcifimemaddr_6 & (\Add0~7  $ (GND))) # (!pcifimemaddr_6 & (!\Add0~7  & VCC))
// \Add0~9  = CARRY((pcifimemaddr_6 & !\Add0~7 ))

	.dataa(gnd),
	.datab(pcifimemaddr_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
// synopsys translate_off
defparam \Add0~8 .lut_mask = 16'hC30C;
defparam \Add0~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N12
cycloneive_lcell_comb \Add0~10 (
// Equation(s):
// \Add0~10_combout  = (pcifimemaddr_7 & (!\Add0~9 )) # (!pcifimemaddr_7 & ((\Add0~9 ) # (GND)))
// \Add0~11  = CARRY((!\Add0~9 ) # (!pcifimemaddr_7))

	.dataa(pcifimemaddr_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
// synopsys translate_off
defparam \Add0~10 .lut_mask = 16'h5A5F;
defparam \Add0~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N14
cycloneive_lcell_comb \Add0~12 (
// Equation(s):
// \Add0~12_combout  = (pcifimemaddr_8 & (\Add0~11  $ (GND))) # (!pcifimemaddr_8 & (!\Add0~11  & VCC))
// \Add0~13  = CARRY((pcifimemaddr_8 & !\Add0~11 ))

	.dataa(gnd),
	.datab(pcifimemaddr_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
// synopsys translate_off
defparam \Add0~12 .lut_mask = 16'hC30C;
defparam \Add0~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N16
cycloneive_lcell_comb \Add0~14 (
// Equation(s):
// \Add0~14_combout  = (pcifimemaddr_9 & (!\Add0~13 )) # (!pcifimemaddr_9 & ((\Add0~13 ) # (GND)))
// \Add0~15  = CARRY((!\Add0~13 ) # (!pcifimemaddr_9))

	.dataa(pcifimemaddr_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
// synopsys translate_off
defparam \Add0~14 .lut_mask = 16'h5A5F;
defparam \Add0~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N18
cycloneive_lcell_comb \Add0~16 (
// Equation(s):
// \Add0~16_combout  = (pcifimemaddr_10 & (\Add0~15  $ (GND))) # (!pcifimemaddr_10 & (!\Add0~15  & VCC))
// \Add0~17  = CARRY((pcifimemaddr_10 & !\Add0~15 ))

	.dataa(gnd),
	.datab(pcifimemaddr_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
// synopsys translate_off
defparam \Add0~16 .lut_mask = 16'hC30C;
defparam \Add0~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N20
cycloneive_lcell_comb \Add0~18 (
// Equation(s):
// \Add0~18_combout  = (pcifimemaddr_11 & (!\Add0~17 )) # (!pcifimemaddr_11 & ((\Add0~17 ) # (GND)))
// \Add0~19  = CARRY((!\Add0~17 ) # (!pcifimemaddr_11))

	.dataa(pcifimemaddr_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
// synopsys translate_off
defparam \Add0~18 .lut_mask = 16'h5A5F;
defparam \Add0~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N22
cycloneive_lcell_comb \Add0~20 (
// Equation(s):
// \Add0~20_combout  = (pcifimemaddr_12 & (\Add0~19  $ (GND))) # (!pcifimemaddr_12 & (!\Add0~19  & VCC))
// \Add0~21  = CARRY((pcifimemaddr_12 & !\Add0~19 ))

	.dataa(gnd),
	.datab(pcifimemaddr_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
// synopsys translate_off
defparam \Add0~20 .lut_mask = 16'hC30C;
defparam \Add0~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N24
cycloneive_lcell_comb \Add0~22 (
// Equation(s):
// \Add0~22_combout  = (pcifimemaddr_13 & (!\Add0~21 )) # (!pcifimemaddr_13 & ((\Add0~21 ) # (GND)))
// \Add0~23  = CARRY((!\Add0~21 ) # (!pcifimemaddr_13))

	.dataa(pcifimemaddr_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
// synopsys translate_off
defparam \Add0~22 .lut_mask = 16'h5A5F;
defparam \Add0~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N26
cycloneive_lcell_comb \Add0~24 (
// Equation(s):
// \Add0~24_combout  = (pcifimemaddr_14 & (\Add0~23  $ (GND))) # (!pcifimemaddr_14 & (!\Add0~23  & VCC))
// \Add0~25  = CARRY((pcifimemaddr_14 & !\Add0~23 ))

	.dataa(gnd),
	.datab(pcifimemaddr_14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
// synopsys translate_off
defparam \Add0~24 .lut_mask = 16'hC30C;
defparam \Add0~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N28
cycloneive_lcell_comb \Add0~26 (
// Equation(s):
// \Add0~26_combout  = (pcifimemaddr_15 & (!\Add0~25 )) # (!pcifimemaddr_15 & ((\Add0~25 ) # (GND)))
// \Add0~27  = CARRY((!\Add0~25 ) # (!pcifimemaddr_15))

	.dataa(pcifimemaddr_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout(\Add0~27 ));
// synopsys translate_off
defparam \Add0~26 .lut_mask = 16'h5A5F;
defparam \Add0~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y39_N30
cycloneive_lcell_comb \Add0~28 (
// Equation(s):
// \Add0~28_combout  = (pcifimemaddr_16 & (\Add0~27  $ (GND))) # (!pcifimemaddr_16 & (!\Add0~27  & VCC))
// \Add0~29  = CARRY((pcifimemaddr_16 & !\Add0~27 ))

	.dataa(gnd),
	.datab(pcifimemaddr_16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~27 ),
	.combout(\Add0~28_combout ),
	.cout(\Add0~29 ));
// synopsys translate_off
defparam \Add0~28 .lut_mask = 16'hC30C;
defparam \Add0~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N0
cycloneive_lcell_comb \Add0~30 (
// Equation(s):
// \Add0~30_combout  = (pcifimemaddr_17 & (!\Add0~29 )) # (!pcifimemaddr_17 & ((\Add0~29 ) # (GND)))
// \Add0~31  = CARRY((!\Add0~29 ) # (!pcifimemaddr_17))

	.dataa(gnd),
	.datab(pcifimemaddr_17),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~29 ),
	.combout(\Add0~30_combout ),
	.cout(\Add0~31 ));
// synopsys translate_off
defparam \Add0~30 .lut_mask = 16'h3C3F;
defparam \Add0~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N2
cycloneive_lcell_comb \Add0~32 (
// Equation(s):
// \Add0~32_combout  = (pcifimemaddr_18 & (\Add0~31  $ (GND))) # (!pcifimemaddr_18 & (!\Add0~31  & VCC))
// \Add0~33  = CARRY((pcifimemaddr_18 & !\Add0~31 ))

	.dataa(gnd),
	.datab(pcifimemaddr_18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~31 ),
	.combout(\Add0~32_combout ),
	.cout(\Add0~33 ));
// synopsys translate_off
defparam \Add0~32 .lut_mask = 16'hC30C;
defparam \Add0~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N4
cycloneive_lcell_comb \Add0~34 (
// Equation(s):
// \Add0~34_combout  = (pcifimemaddr_19 & (!\Add0~33 )) # (!pcifimemaddr_19 & ((\Add0~33 ) # (GND)))
// \Add0~35  = CARRY((!\Add0~33 ) # (!pcifimemaddr_19))

	.dataa(gnd),
	.datab(pcifimemaddr_19),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~33 ),
	.combout(\Add0~34_combout ),
	.cout(\Add0~35 ));
// synopsys translate_off
defparam \Add0~34 .lut_mask = 16'h3C3F;
defparam \Add0~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N6
cycloneive_lcell_comb \Add0~36 (
// Equation(s):
// \Add0~36_combout  = (pcifimemaddr_20 & (\Add0~35  $ (GND))) # (!pcifimemaddr_20 & (!\Add0~35  & VCC))
// \Add0~37  = CARRY((pcifimemaddr_20 & !\Add0~35 ))

	.dataa(pcifimemaddr_20),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~35 ),
	.combout(\Add0~36_combout ),
	.cout(\Add0~37 ));
// synopsys translate_off
defparam \Add0~36 .lut_mask = 16'hA50A;
defparam \Add0~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N8
cycloneive_lcell_comb \Add0~38 (
// Equation(s):
// \Add0~38_combout  = (pcifimemaddr_21 & (!\Add0~37 )) # (!pcifimemaddr_21 & ((\Add0~37 ) # (GND)))
// \Add0~39  = CARRY((!\Add0~37 ) # (!pcifimemaddr_21))

	.dataa(gnd),
	.datab(pcifimemaddr_21),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~37 ),
	.combout(\Add0~38_combout ),
	.cout(\Add0~39 ));
// synopsys translate_off
defparam \Add0~38 .lut_mask = 16'h3C3F;
defparam \Add0~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N10
cycloneive_lcell_comb \Add0~40 (
// Equation(s):
// \Add0~40_combout  = (pcifimemaddr_22 & (\Add0~39  $ (GND))) # (!pcifimemaddr_22 & (!\Add0~39  & VCC))
// \Add0~41  = CARRY((pcifimemaddr_22 & !\Add0~39 ))

	.dataa(pcifimemaddr_22),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~39 ),
	.combout(\Add0~40_combout ),
	.cout(\Add0~41 ));
// synopsys translate_off
defparam \Add0~40 .lut_mask = 16'hA50A;
defparam \Add0~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N12
cycloneive_lcell_comb \Add0~42 (
// Equation(s):
// \Add0~42_combout  = (pcifimemaddr_23 & (!\Add0~41 )) # (!pcifimemaddr_23 & ((\Add0~41 ) # (GND)))
// \Add0~43  = CARRY((!\Add0~41 ) # (!pcifimemaddr_23))

	.dataa(pcifimemaddr_23),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~41 ),
	.combout(\Add0~42_combout ),
	.cout(\Add0~43 ));
// synopsys translate_off
defparam \Add0~42 .lut_mask = 16'h5A5F;
defparam \Add0~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N14
cycloneive_lcell_comb \Add0~44 (
// Equation(s):
// \Add0~44_combout  = (pcifimemaddr_24 & (\Add0~43  $ (GND))) # (!pcifimemaddr_24 & (!\Add0~43  & VCC))
// \Add0~45  = CARRY((pcifimemaddr_24 & !\Add0~43 ))

	.dataa(pcifimemaddr_24),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~43 ),
	.combout(\Add0~44_combout ),
	.cout(\Add0~45 ));
// synopsys translate_off
defparam \Add0~44 .lut_mask = 16'hA50A;
defparam \Add0~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N16
cycloneive_lcell_comb \Add0~46 (
// Equation(s):
// \Add0~46_combout  = (pcifimemaddr_25 & (!\Add0~45 )) # (!pcifimemaddr_25 & ((\Add0~45 ) # (GND)))
// \Add0~47  = CARRY((!\Add0~45 ) # (!pcifimemaddr_25))

	.dataa(gnd),
	.datab(pcifimemaddr_25),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~45 ),
	.combout(\Add0~46_combout ),
	.cout(\Add0~47 ));
// synopsys translate_off
defparam \Add0~46 .lut_mask = 16'h3C3F;
defparam \Add0~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N18
cycloneive_lcell_comb \Add0~48 (
// Equation(s):
// \Add0~48_combout  = (pcifimemaddr_26 & (\Add0~47  $ (GND))) # (!pcifimemaddr_26 & (!\Add0~47  & VCC))
// \Add0~49  = CARRY((pcifimemaddr_26 & !\Add0~47 ))

	.dataa(pcifimemaddr_26),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~47 ),
	.combout(\Add0~48_combout ),
	.cout(\Add0~49 ));
// synopsys translate_off
defparam \Add0~48 .lut_mask = 16'hA50A;
defparam \Add0~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N20
cycloneive_lcell_comb \Add0~50 (
// Equation(s):
// \Add0~50_combout  = (pcifimemaddr_27 & (!\Add0~49 )) # (!pcifimemaddr_27 & ((\Add0~49 ) # (GND)))
// \Add0~51  = CARRY((!\Add0~49 ) # (!pcifimemaddr_27))

	.dataa(pcifimemaddr_27),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~49 ),
	.combout(\Add0~50_combout ),
	.cout(\Add0~51 ));
// synopsys translate_off
defparam \Add0~50 .lut_mask = 16'h5A5F;
defparam \Add0~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N22
cycloneive_lcell_comb \Add0~52 (
// Equation(s):
// \Add0~52_combout  = (pcifimemaddr_28 & (\Add0~51  $ (GND))) # (!pcifimemaddr_28 & (!\Add0~51  & VCC))
// \Add0~53  = CARRY((pcifimemaddr_28 & !\Add0~51 ))

	.dataa(pcifimemaddr_28),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~51 ),
	.combout(\Add0~52_combout ),
	.cout(\Add0~53 ));
// synopsys translate_off
defparam \Add0~52 .lut_mask = 16'hA50A;
defparam \Add0~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N24
cycloneive_lcell_comb \Add0~54 (
// Equation(s):
// \Add0~54_combout  = (pcifimemaddr_29 & (!\Add0~53 )) # (!pcifimemaddr_29 & ((\Add0~53 ) # (GND)))
// \Add0~55  = CARRY((!\Add0~53 ) # (!pcifimemaddr_29))

	.dataa(pcifimemaddr_29),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~53 ),
	.combout(\Add0~54_combout ),
	.cout(\Add0~55 ));
// synopsys translate_off
defparam \Add0~54 .lut_mask = 16'h5A5F;
defparam \Add0~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N26
cycloneive_lcell_comb \Add0~56 (
// Equation(s):
// \Add0~56_combout  = (pcifimemaddr_30 & (\Add0~55  $ (GND))) # (!pcifimemaddr_30 & (!\Add0~55  & VCC))
// \Add0~57  = CARRY((pcifimemaddr_30 & !\Add0~55 ))

	.dataa(gnd),
	.datab(pcifimemaddr_30),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~55 ),
	.combout(\Add0~56_combout ),
	.cout(\Add0~57 ));
// synopsys translate_off
defparam \Add0~56 .lut_mask = 16'hC30C;
defparam \Add0~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y38_N28
cycloneive_lcell_comb \Add0~58 (
// Equation(s):
// \Add0~58_combout  = pcifimemaddr_31 $ (\Add0~57 )

	.dataa(gnd),
	.datab(pcifimemaddr_31),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~57 ),
	.combout(\Add0~58_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~58 .lut_mask = 16'h3C3C;
defparam \Add0~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N8
cycloneive_lcell_comb \WideOr0~0 (
// Equation(s):
// \WideOr0~0_combout  = (dcifimemload_31 & (dcifimemload_27 & (dcifimemload_26))) # (!dcifimemload_31 & (((dcifimemload_29))))

	.dataa(dcifimemload_27),
	.datab(dcifimemload_26),
	.datac(dcifimemload_31),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(\WideOr0~0_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr0~0 .lut_mask = 16'h8F80;
defparam \WideOr0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N30
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// \Mux5~0_combout  = ((\WideOr0~0_combout  & (!dcifimemload_30 & !dcifimemload_28))) # (!cuifaluSrc_0)

	.dataa(\WideOr0~0_combout ),
	.datab(dcifimemload_30),
	.datac(dcifimemload_28),
	.datad(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'h02FF;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N20
cycloneive_lcell_comb \Mux5~1 (
// Equation(s):
// \Mux5~1_combout  = (dcifimemload_15 & (!cuifaluSrc_1 & (\Mux5~0_combout  & cuifaluSrc_0)))

	.dataa(dcifimemload_15),
	.datab(\cu_dut|cuif.aluSrc[1]~1_combout ),
	.datac(\Mux5~0_combout ),
	.datad(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~1 .lut_mask = 16'h2000;
defparam \Mux5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N14
cycloneive_lcell_comb \Mux5~2 (
// Equation(s):
// \Mux5~2_combout  = (!cuifaluSrc_1 & (\Mux5~0_combout  & (!cuifregT_4 & !cuifaluSrc_0)))

	.dataa(\cu_dut|cuif.aluSrc[1]~1_combout ),
	.datab(\Mux5~0_combout ),
	.datac(cuifregT_4),
	.datad(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~2 .lut_mask = 16'h0004;
defparam \Mux5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N26
cycloneive_lcell_comb \Mux5~3 (
// Equation(s):
// \Mux5~3_combout  = (\Mux5~0_combout  & (cuifregT_4 & (!cuifaluSrc_1 & !cuifaluSrc_0)))

	.dataa(\Mux5~0_combout ),
	.datab(cuifregT_4),
	.datac(\cu_dut|cuif.aluSrc[1]~1_combout ),
	.datad(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~3 .lut_mask = 16'h0008;
defparam \Mux5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N12
cycloneive_lcell_comb \Mux5~4 (
// Equation(s):
// \Mux5~4_combout  = (\Mux5~2_combout  & ((Mux321) # ((\Mux5~3_combout  & Mux32)))) # (!\Mux5~2_combout  & (\Mux5~3_combout  & (Mux32)))

	.dataa(\Mux5~2_combout ),
	.datab(\Mux5~3_combout ),
	.datac(Mux32),
	.datad(Mux321),
	.cin(gnd),
	.combout(\Mux5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~4 .lut_mask = 16'hEAC0;
defparam \Mux5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N28
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// \Mux6~0_combout  = (\Mux5~2_combout  & ((Mux33) # ((\Mux5~3_combout  & Mux331)))) # (!\Mux5~2_combout  & (\Mux5~3_combout  & ((Mux331))))

	.dataa(\Mux5~2_combout ),
	.datab(\Mux5~3_combout ),
	.datac(Mux33),
	.datad(Mux331),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'hECA0;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N24
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (Mux34 & \Mux5~3_combout )

	.dataa(Mux34),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux5~3_combout ),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hAA00;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N4
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// \Mux7~1_combout  = (\Mux5~1_combout ) # ((\Mux7~0_combout ) # ((\Mux5~2_combout  & Mux341)))

	.dataa(\Mux5~1_combout ),
	.datab(\Mux7~0_combout ),
	.datac(\Mux5~2_combout ),
	.datad(Mux341),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hFEEE;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N2
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// \Mux8~0_combout  = (\Mux5~2_combout  & ((Mux35) # ((\Mux5~3_combout  & Mux351)))) # (!\Mux5~2_combout  & (\Mux5~3_combout  & (Mux351)))

	.dataa(\Mux5~2_combout ),
	.datab(\Mux5~3_combout ),
	.datac(Mux351),
	.datad(Mux35),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hEAC0;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N6
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// \Mux9~0_combout  = (\Mux5~2_combout  & ((Mux36) # ((\Mux5~3_combout  & Mux361)))) # (!\Mux5~2_combout  & (\Mux5~3_combout  & (Mux361)))

	.dataa(\Mux5~2_combout ),
	.datab(\Mux5~3_combout ),
	.datac(Mux361),
	.datad(Mux36),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hEAC0;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N18
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// \Mux10~0_combout  = (\Mux5~2_combout  & ((Mux37) # ((\Mux5~3_combout  & Mux371)))) # (!\Mux5~2_combout  & (\Mux5~3_combout  & ((Mux371))))

	.dataa(\Mux5~2_combout ),
	.datab(\Mux5~3_combout ),
	.datac(Mux37),
	.datad(Mux371),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hECA0;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N2
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// \Mux11~0_combout  = (\Mux5~2_combout  & ((Mux38) # ((Mux381 & \Mux5~3_combout )))) # (!\Mux5~2_combout  & (((Mux381 & \Mux5~3_combout ))))

	.dataa(\Mux5~2_combout ),
	.datab(Mux38),
	.datac(Mux381),
	.datad(\Mux5~3_combout ),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hF888;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N6
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (Mux39 & \Mux5~3_combout )

	.dataa(gnd),
	.datab(Mux39),
	.datac(gnd),
	.datad(\Mux5~3_combout ),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hCC00;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N16
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// \Mux12~1_combout  = (\Mux5~1_combout ) # ((\Mux12~0_combout ) # ((\Mux5~2_combout  & Mux391)))

	.dataa(\Mux5~2_combout ),
	.datab(\Mux5~1_combout ),
	.datac(Mux391),
	.datad(\Mux12~0_combout ),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hFFEC;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N22
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// \Mux13~0_combout  = (\Mux5~3_combout  & ((Mux401) # ((Mux40 & \Mux5~2_combout )))) # (!\Mux5~3_combout  & (Mux40 & (\Mux5~2_combout )))

	.dataa(\Mux5~3_combout ),
	.datab(Mux40),
	.datac(\Mux5~2_combout ),
	.datad(Mux401),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hEAC0;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N16
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// \Mux14~0_combout  = (\Mux5~2_combout  & ((Mux41) # ((\Mux5~3_combout  & Mux411)))) # (!\Mux5~2_combout  & (\Mux5~3_combout  & (Mux411)))

	.dataa(\Mux5~2_combout ),
	.datab(\Mux5~3_combout ),
	.datac(Mux411),
	.datad(Mux41),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hEAC0;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N6
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// \Mux14~1_combout  = (\Mux5~1_combout ) # (\Mux14~0_combout )

	.dataa(\Mux5~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux14~0_combout ),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hFFAA;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N12
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// \Mux15~0_combout  = (\Mux5~3_combout  & ((Mux421) # ((\Mux5~2_combout  & Mux42)))) # (!\Mux5~3_combout  & (\Mux5~2_combout  & (Mux42)))

	.dataa(\Mux5~3_combout ),
	.datab(\Mux5~2_combout ),
	.datac(Mux42),
	.datad(Mux421),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hEAC0;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N14
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// \Mux15~1_combout  = (\Mux5~1_combout ) # (\Mux15~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Mux5~1_combout ),
	.datad(\Mux15~0_combout ),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'hFFF0;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N26
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// \Mux16~0_combout  = (\Mux5~2_combout  & ((Mux43) # ((Mux431 & \Mux5~3_combout )))) # (!\Mux5~2_combout  & (Mux431 & (\Mux5~3_combout )))

	.dataa(\Mux5~2_combout ),
	.datab(Mux431),
	.datac(\Mux5~3_combout ),
	.datad(Mux43),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'hEAC0;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N12
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// \Mux16~1_combout  = (\Mux16~0_combout ) # (\Mux5~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Mux16~0_combout ),
	.datad(\Mux5~1_combout ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hFFF0;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N14
cycloneive_lcell_comb \Mux36~0 (
// Equation(s):
// \Mux36~0_combout  = (!cuifregT_4 & (!cuifaluSrc_0 & !cuifaluSrc_1))

	.dataa(cuifregT_4),
	.datab(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.datac(gnd),
	.datad(\cu_dut|cuif.aluSrc[1]~1_combout ),
	.cin(gnd),
	.combout(\Mux36~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~0 .lut_mask = 16'h0011;
defparam \Mux36~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N10
cycloneive_lcell_comb \Mux31~0 (
// Equation(s):
// \Mux31~0_combout  = (cuifaluSrc_0 & ((dcifimemload_5) # ((\Mux36~0_combout  & Mux58)))) # (!cuifaluSrc_0 & (((\Mux36~0_combout  & Mux58))))

	.dataa(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.datab(dcifimemload_5),
	.datac(\Mux36~0_combout ),
	.datad(Mux58),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~0 .lut_mask = 16'hF888;
defparam \Mux31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N20
cycloneive_lcell_comb \Mux36~1 (
// Equation(s):
// \Mux36~1_combout  = (cuifregT_4 & (!cuifaluSrc_0 & !cuifaluSrc_1))

	.dataa(cuifregT_4),
	.datab(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.datac(gnd),
	.datad(\cu_dut|cuif.aluSrc[1]~1_combout ),
	.cin(gnd),
	.combout(\Mux36~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~1 .lut_mask = 16'h0022;
defparam \Mux36~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N12
cycloneive_lcell_comb \Mux31~1 (
// Equation(s):
// \Mux31~1_combout  = (\Mux31~0_combout ) # ((\Mux36~1_combout  & Mux581))

	.dataa(gnd),
	.datab(\Mux36~1_combout ),
	.datac(Mux581),
	.datad(\Mux31~0_combout ),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~1 .lut_mask = 16'hFFC0;
defparam \Mux31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N16
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// \Mux17~0_combout  = (\Mux5~2_combout  & ((Mux44) # ((\Mux5~3_combout  & Mux441)))) # (!\Mux5~2_combout  & (\Mux5~3_combout  & ((Mux441))))

	.dataa(\Mux5~2_combout ),
	.datab(\Mux5~3_combout ),
	.datac(Mux44),
	.datad(Mux441),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'hECA0;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N30
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// \Mux18~0_combout  = (\Mux5~2_combout  & ((Mux45) # ((\Mux5~3_combout  & Mux451)))) # (!\Mux5~2_combout  & (((\Mux5~3_combout  & Mux451))))

	.dataa(\Mux5~2_combout ),
	.datab(Mux45),
	.datac(\Mux5~3_combout ),
	.datad(Mux451),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'hF888;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N24
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (\Mux5~2_combout  & ((Mux46) # ((\Mux5~3_combout  & Mux461)))) # (!\Mux5~2_combout  & (\Mux5~3_combout  & (Mux461)))

	.dataa(\Mux5~2_combout ),
	.datab(\Mux5~3_combout ),
	.datac(Mux461),
	.datad(Mux46),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'hEAC0;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N12
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// \Mux20~0_combout  = (\Mux5~3_combout  & Mux47)

	.dataa(gnd),
	.datab(gnd),
	.datac(\Mux5~3_combout ),
	.datad(Mux47),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'hF000;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N20
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// \Mux20~1_combout  = (\Mux5~1_combout ) # ((\Mux20~0_combout ) # ((\Mux5~2_combout  & Mux471)))

	.dataa(\Mux5~2_combout ),
	.datab(Mux471),
	.datac(\Mux5~1_combout ),
	.datad(\Mux20~0_combout ),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'hFFF8;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N8
cycloneive_lcell_comb \Mux5~5 (
// Equation(s):
// \Mux5~5_combout  = (dcifimemload_15 & ((Equal2 & ((dcifimemload_29))) # (!Equal2 & (!cuifregT_0))))

	.dataa(\cu_dut|cuif.regT[0]~1_combout ),
	.datab(\cu_dut|Equal2~4_combout ),
	.datac(dcifimemload_15),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(\Mux5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~5 .lut_mask = 16'hD010;
defparam \Mux5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N22
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// \Mux21~0_combout  = (\Mux36~0_combout  & ((Mux48) # ((!cuifaluSrc_1 & \Mux5~5_combout )))) # (!\Mux36~0_combout  & (!cuifaluSrc_1 & (\Mux5~5_combout )))

	.dataa(\Mux36~0_combout ),
	.datab(\cu_dut|cuif.aluSrc[1]~1_combout ),
	.datac(\Mux5~5_combout ),
	.datad(Mux48),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hBA30;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N24
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// \Mux21~1_combout  = (\Mux21~0_combout ) # ((\Mux36~1_combout  & Mux481))

	.dataa(gnd),
	.datab(\Mux36~1_combout ),
	.datac(\Mux21~0_combout ),
	.datad(Mux481),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'hFCF0;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N0
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// \Mux22~0_combout  = (\Mux35~5_combout  & ((dcifimemload_14) # ((\Mux36~0_combout  & Mux49)))) # (!\Mux35~5_combout  & (((\Mux36~0_combout  & Mux49))))

	.dataa(\Mux35~5_combout ),
	.datab(dcifimemload_14),
	.datac(\Mux36~0_combout ),
	.datad(Mux49),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'hF888;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N24
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// \Mux22~1_combout  = (\Mux22~0_combout ) # ((\Mux36~1_combout  & Mux491))

	.dataa(gnd),
	.datab(\Mux36~1_combout ),
	.datac(Mux491),
	.datad(\Mux22~0_combout ),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'hFFC0;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N20
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// \Mux23~0_combout  = (\Mux36~0_combout  & ((Mux50) # ((dcifimemload_13 & \Mux35~5_combout )))) # (!\Mux36~0_combout  & (dcifimemload_13 & (\Mux35~5_combout )))

	.dataa(\Mux36~0_combout ),
	.datab(dcifimemload_13),
	.datac(\Mux35~5_combout ),
	.datad(Mux50),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hEAC0;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N22
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// \Mux23~1_combout  = (\Mux23~0_combout ) # ((Mux501 & \Mux36~1_combout ))

	.dataa(gnd),
	.datab(Mux501),
	.datac(\Mux36~1_combout ),
	.datad(\Mux23~0_combout ),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'hFFC0;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N12
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (dcifimemload_12 & ((\Mux35~5_combout ) # ((\Mux36~0_combout  & Mux51)))) # (!dcifimemload_12 & (((\Mux36~0_combout  & Mux51))))

	.dataa(dcifimemload_12),
	.datab(\Mux35~5_combout ),
	.datac(\Mux36~0_combout ),
	.datad(Mux51),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'hF888;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N10
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// \Mux24~1_combout  = (\Mux24~0_combout ) # ((\Mux36~1_combout  & Mux511))

	.dataa(\Mux36~1_combout ),
	.datab(gnd),
	.datac(Mux511),
	.datad(\Mux24~0_combout ),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'hFFA0;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N8
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (dcifimemload_11 & ((\Mux35~5_combout ) # ((Mux52 & \Mux36~0_combout )))) # (!dcifimemload_11 & (((Mux52 & \Mux36~0_combout ))))

	.dataa(dcifimemload_11),
	.datab(\Mux35~5_combout ),
	.datac(Mux52),
	.datad(\Mux36~0_combout ),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hF888;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N0
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// \Mux25~1_combout  = (\Mux25~0_combout ) # ((\Mux36~1_combout  & Mux521))

	.dataa(gnd),
	.datab(\Mux36~1_combout ),
	.datac(\Mux25~0_combout ),
	.datad(Mux521),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hFCF0;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N16
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (\Mux36~0_combout  & ((Mux53) # ((dcifimemload_10 & \Mux35~5_combout )))) # (!\Mux36~0_combout  & (dcifimemload_10 & (\Mux35~5_combout )))

	.dataa(\Mux36~0_combout ),
	.datab(dcifimemload_10),
	.datac(\Mux35~5_combout ),
	.datad(Mux53),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hEAC0;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N14
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// \Mux26~1_combout  = (\Mux26~0_combout ) # ((\Mux36~1_combout  & Mux531))

	.dataa(\Mux36~1_combout ),
	.datab(gnd),
	.datac(Mux531),
	.datad(\Mux26~0_combout ),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hFFA0;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N8
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (\Mux35~5_combout  & ((dcifimemload_9) # ((\Mux36~0_combout  & Mux54)))) # (!\Mux35~5_combout  & (\Mux36~0_combout  & ((Mux54))))

	.dataa(\Mux35~5_combout ),
	.datab(\Mux36~0_combout ),
	.datac(dcifimemload_9),
	.datad(Mux54),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'hECA0;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N18
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// \Mux27~1_combout  = (\Mux27~0_combout ) # ((Mux541 & \Mux36~1_combout ))

	.dataa(gnd),
	.datab(Mux541),
	.datac(\Mux27~0_combout ),
	.datad(\Mux36~1_combout ),
	.cin(gnd),
	.combout(\Mux27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hFCF0;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N16
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (\Mux35~5_combout  & ((dcifimemload_8) # ((\Mux36~0_combout  & Mux55)))) # (!\Mux35~5_combout  & (((\Mux36~0_combout  & Mux55))))

	.dataa(\Mux35~5_combout ),
	.datab(dcifimemload_8),
	.datac(\Mux36~0_combout ),
	.datad(Mux55),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'hF888;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N30
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// \Mux28~1_combout  = (\Mux28~0_combout ) # ((\Mux36~1_combout  & Mux551))

	.dataa(\Mux36~1_combout ),
	.datab(Mux551),
	.datac(gnd),
	.datad(\Mux28~0_combout ),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hFF88;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N2
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (\Mux35~5_combout  & ((dcifimemload_7) # ((\Mux36~0_combout  & Mux56)))) # (!\Mux35~5_combout  & (((\Mux36~0_combout  & Mux56))))

	.dataa(\Mux35~5_combout ),
	.datab(dcifimemload_7),
	.datac(\Mux36~0_combout ),
	.datad(Mux56),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'hF888;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N28
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// \Mux29~1_combout  = (\Mux29~0_combout ) # ((\Mux36~1_combout  & Mux561))

	.dataa(gnd),
	.datab(\Mux36~1_combout ),
	.datac(Mux561),
	.datad(\Mux29~0_combout ),
	.cin(gnd),
	.combout(\Mux29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'hFFC0;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N30
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// \Mux30~0_combout  = (\Mux36~0_combout  & ((Mux57) # ((dcifimemload_6 & \Mux35~5_combout )))) # (!\Mux36~0_combout  & (dcifimemload_6 & ((\Mux35~5_combout ))))

	.dataa(\Mux36~0_combout ),
	.datab(dcifimemload_6),
	.datac(Mux57),
	.datad(\Mux35~5_combout ),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'hECA0;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N20
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// \Mux30~1_combout  = (\Mux30~0_combout ) # ((\Mux36~1_combout  & Mux571))

	.dataa(gnd),
	.datab(\Mux36~1_combout ),
	.datac(\Mux30~0_combout ),
	.datad(Mux571),
	.cin(gnd),
	.combout(\Mux30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'hFCF0;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N30
cycloneive_lcell_comb \Mux36~2 (
// Equation(s):
// \Mux36~2_combout  = (!cuifaluSrc_1 & (!cuifaluSrc_0 & (cuifregT_4 & Mux63)))

	.dataa(\cu_dut|cuif.aluSrc[1]~1_combout ),
	.datab(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.datac(cuifregT_4),
	.datad(Mux63),
	.cin(gnd),
	.combout(\Mux36~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~2 .lut_mask = 16'h1000;
defparam \Mux36~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N10
cycloneive_lcell_comb \Mux32~2 (
// Equation(s):
// \Mux32~2_combout  = (!cuifaluSrc_0 & (!Equal0 & cuifaluSrc_1))

	.dataa(gnd),
	.datab(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.datac(\cu_dut|Equal0~0_combout ),
	.datad(\cu_dut|cuif.aluSrc[1]~1_combout ),
	.cin(gnd),
	.combout(\Mux32~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~2 .lut_mask = 16'h0300;
defparam \Mux32~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N4
cycloneive_lcell_comb \Mux36~3 (
// Equation(s):
// \Mux36~3_combout  = (\Mux32~2_combout  & ((dcifimemload_6) # ((dcifimemload_0 & cuifaluSrc_0)))) # (!\Mux32~2_combout  & (dcifimemload_0 & ((cuifaluSrc_0))))

	.dataa(\Mux32~2_combout ),
	.datab(dcifimemload_0),
	.datac(dcifimemload_6),
	.datad(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux36~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~3 .lut_mask = 16'hECA0;
defparam \Mux36~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N10
cycloneive_lcell_comb \Mux36~4 (
// Equation(s):
// \Mux36~4_combout  = (\Mux36~3_combout ) # ((\Mux36~2_combout ) # ((\Mux36~0_combout  & Mux631)))

	.dataa(\Mux36~3_combout ),
	.datab(\Mux36~0_combout ),
	.datac(\Mux36~2_combout ),
	.datad(Mux631),
	.cin(gnd),
	.combout(\Mux36~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~4 .lut_mask = 16'hFEFA;
defparam \Mux36~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N10
cycloneive_lcell_comb \Mux35~2 (
// Equation(s):
// \Mux35~2_combout  = (\Mux36~0_combout  & ((Mux62) # ((\Mux36~1_combout  & Mux621)))) # (!\Mux36~0_combout  & (\Mux36~1_combout  & (Mux621)))

	.dataa(\Mux36~0_combout ),
	.datab(\Mux36~1_combout ),
	.datac(Mux621),
	.datad(Mux62),
	.cin(gnd),
	.combout(\Mux35~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~2 .lut_mask = 16'hEAC0;
defparam \Mux35~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N16
cycloneive_lcell_comb \Mux35~3 (
// Equation(s):
// \Mux35~3_combout  = (dcifimemload_7 & ((\Mux32~2_combout ) # ((dcifimemload_1 & \Mux35~5_combout )))) # (!dcifimemload_7 & (dcifimemload_1 & (\Mux35~5_combout )))

	.dataa(dcifimemload_7),
	.datab(dcifimemload_1),
	.datac(\Mux35~5_combout ),
	.datad(\Mux32~2_combout ),
	.cin(gnd),
	.combout(\Mux35~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~3 .lut_mask = 16'hEAC0;
defparam \Mux35~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N20
cycloneive_lcell_comb \Mux35~4 (
// Equation(s):
// \Mux35~4_combout  = (\Mux35~3_combout ) # (\Mux35~2_combout )

	.dataa(gnd),
	.datab(\Mux35~3_combout ),
	.datac(gnd),
	.datad(\Mux35~2_combout ),
	.cin(gnd),
	.combout(\Mux35~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~4 .lut_mask = 16'hFFCC;
defparam \Mux35~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N8
cycloneive_lcell_comb \Mux34~2 (
// Equation(s):
// \Mux34~2_combout  = (dcifimemload_2 & ((cuifaluSrc_0) # ((dcifimemload_8 & \Mux32~2_combout )))) # (!dcifimemload_2 & (dcifimemload_8 & (\Mux32~2_combout )))

	.dataa(dcifimemload_2),
	.datab(dcifimemload_8),
	.datac(\Mux32~2_combout ),
	.datad(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux34~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~2 .lut_mask = 16'hEAC0;
defparam \Mux34~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N10
cycloneive_lcell_comb \Mux34~3 (
// Equation(s):
// \Mux34~3_combout  = (\Mux34~2_combout ) # ((\Mux34~4_combout ) # ((\Mux36~0_combout  & Mux611)))

	.dataa(\Mux36~0_combout ),
	.datab(\Mux34~2_combout ),
	.datac(\Mux34~4_combout ),
	.datad(Mux611),
	.cin(gnd),
	.combout(\Mux34~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~3 .lut_mask = 16'hFEFC;
defparam \Mux34~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N4
cycloneive_lcell_comb \Mux33~2 (
// Equation(s):
// \Mux33~2_combout  = (dcifimemload_3 & ((cuifaluSrc_0) # ((dcifimemload_9 & \Mux32~2_combout )))) # (!dcifimemload_3 & (((dcifimemload_9 & \Mux32~2_combout ))))

	.dataa(dcifimemload_3),
	.datab(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.datac(dcifimemload_9),
	.datad(\Mux32~2_combout ),
	.cin(gnd),
	.combout(\Mux33~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~2 .lut_mask = 16'hF888;
defparam \Mux33~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N20
cycloneive_lcell_comb \Mux33~3 (
// Equation(s):
// \Mux33~3_combout  = (\Mux33~2_combout ) # ((\Mux33~4_combout ) # ((\Mux36~0_combout  & Mux601)))

	.dataa(\Mux36~0_combout ),
	.datab(\Mux33~2_combout ),
	.datac(\Mux33~4_combout ),
	.datad(Mux601),
	.cin(gnd),
	.combout(\Mux33~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~3 .lut_mask = 16'hFEFC;
defparam \Mux33~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N28
cycloneive_lcell_comb \Mux32~3 (
// Equation(s):
// \Mux32~3_combout  = (cuifaluSrc_0 & ((dcifimemload_4) # ((\Mux32~2_combout  & dcifimemload_10)))) # (!cuifaluSrc_0 & (((\Mux32~2_combout  & dcifimemload_10))))

	.dataa(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.datab(dcifimemload_4),
	.datac(\Mux32~2_combout ),
	.datad(dcifimemload_10),
	.cin(gnd),
	.combout(\Mux32~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~3 .lut_mask = 16'hF888;
defparam \Mux32~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N6
cycloneive_lcell_comb \Mux32~4 (
// Equation(s):
// \Mux32~4_combout  = (\Mux32~3_combout ) # ((\Mux32~5_combout ) # ((\Mux36~0_combout  & Mux591)))

	.dataa(\Mux36~0_combout ),
	.datab(\Mux32~3_combout ),
	.datac(\Mux32~5_combout ),
	.datad(Mux591),
	.cin(gnd),
	.combout(\Mux32~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~4 .lut_mask = 16'hFEFC;
defparam \Mux32~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N8
cycloneive_lcell_comb \Mux5~6 (
// Equation(s):
// \Mux5~6_combout  = (\Mux5~1_combout ) # (\Mux5~4_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Mux5~1_combout ),
	.datad(\Mux5~4_combout ),
	.cin(gnd),
	.combout(\Mux5~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~6 .lut_mask = 16'hFFF0;
defparam \Mux5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N24
cycloneive_lcell_comb \Mux6~1 (
// Equation(s):
// \Mux6~1_combout  = (\Mux5~1_combout ) # (\Mux6~0_combout )

	.dataa(\Mux5~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux6~0_combout ),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~1 .lut_mask = 16'hFFAA;
defparam \Mux6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N2
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// \Mux8~1_combout  = (\Mux5~1_combout ) # (\Mux8~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Mux5~1_combout ),
	.datad(\Mux8~0_combout ),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'hFFF0;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N26
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// \Mux9~1_combout  = (\Mux5~1_combout ) # (\Mux9~0_combout )

	.dataa(\Mux5~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux9~0_combout ),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'hFFAA;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N12
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// \Mux10~1_combout  = (\Mux5~1_combout ) # (\Mux10~0_combout )

	.dataa(gnd),
	.datab(\Mux5~1_combout ),
	.datac(gnd),
	.datad(\Mux10~0_combout ),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'hFFCC;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N22
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// \Mux11~1_combout  = (\Mux5~1_combout ) # (\Mux11~0_combout )

	.dataa(gnd),
	.datab(\Mux5~1_combout ),
	.datac(gnd),
	.datad(\Mux11~0_combout ),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'hFFCC;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N24
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// \Mux13~1_combout  = (\Mux13~0_combout ) # (\Mux5~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Mux13~0_combout ),
	.datad(\Mux5~1_combout ),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'hFFF0;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N0
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// \Mux17~1_combout  = (\Mux17~0_combout ) # (\Mux5~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Mux17~0_combout ),
	.datad(\Mux5~1_combout ),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hFFF0;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N0
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// \Mux18~1_combout  = (\Mux5~1_combout ) # (\Mux18~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Mux5~1_combout ),
	.datad(\Mux18~0_combout ),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'hFFF0;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N6
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// \Mux19~1_combout  = (\Mux5~1_combout ) # (\Mux19~0_combout )

	.dataa(\Mux5~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Mux19~0_combout ),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'hFFAA;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N12
cycloneive_lcell_comb \Mux68~0 (
// Equation(s):
// \Mux68~0_combout  = (cuifMemtoReg_1 & (pcifimemaddr_0)) # (!cuifMemtoReg_1 & ((ramiframload_0)))

	.dataa(pcifimemaddr_0),
	.datab(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datac(gnd),
	.datad(ramiframload_0),
	.cin(gnd),
	.combout(\Mux68~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux68~0 .lut_mask = 16'hBB88;
defparam \Mux68~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N0
cycloneive_lcell_comb \Mux68~1 (
// Equation(s):
// \Mux68~1_combout  = (cuifMemtoReg_0 & (((\Mux68~0_combout )))) # (!cuifMemtoReg_0 & (!cuifMemtoReg_1 & ((Selector312))))

	.dataa(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datab(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datac(\Mux68~0_combout ),
	.datad(\alu_dut|Selector31~9_combout ),
	.cin(gnd),
	.combout(\Mux68~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux68~1 .lut_mask = 16'hB1A0;
defparam \Mux68~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N14
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// \Mux0~0_combout  = (!dcifimemload_27 & (!dcifimemload_28 & (!dcifimemload_26 & Equal22)))

	.dataa(dcifimemload_27),
	.datab(dcifimemload_28),
	.datac(dcifimemload_26),
	.datad(\cu_dut|Equal2~8_combout ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'h0100;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N8
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// \Mux4~0_combout  = (\Mux0~0_combout  & dcifimemload_11)

	.dataa(gnd),
	.datab(\Mux0~0_combout ),
	.datac(dcifimemload_11),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'hC0C0;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N14
cycloneive_lcell_comb \Mux4~1 (
// Equation(s):
// \Mux4~1_combout  = (\Mux4~0_combout ) # ((!cuifRegDst_0 & ((cuifregT_01) # (Equal23))))

	.dataa(\Mux4~0_combout ),
	.datab(\cu_dut|cuif.regT[0]~4_combout ),
	.datac(\cu_dut|Equal2~9_combout ),
	.datad(\cu_dut|cuif.RegDst[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~1 .lut_mask = 16'hAAFE;
defparam \Mux4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N6
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// \Mux2~0_combout  = (\Mux0~0_combout  & dcifimemload_13)

	.dataa(gnd),
	.datab(\Mux0~0_combout ),
	.datac(gnd),
	.datad(dcifimemload_13),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'hCC00;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N24
cycloneive_lcell_comb \Mux2~1 (
// Equation(s):
// \Mux2~1_combout  = (\Mux2~0_combout ) # ((!cuifRegDst_0 & ((Equal23) # (cuifregT_2))))

	.dataa(\Mux2~0_combout ),
	.datab(\cu_dut|Equal2~9_combout ),
	.datac(\cu_dut|cuif.regT[2]~3_combout ),
	.datad(\cu_dut|cuif.RegDst[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~1 .lut_mask = 16'hAAFE;
defparam \Mux2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N18
cycloneive_lcell_comb \Mux0~1 (
// Equation(s):
// \Mux0~1_combout  = (\Mux0~0_combout  & dcifimemload_15)

	.dataa(gnd),
	.datab(gnd),
	.datac(\Mux0~0_combout ),
	.datad(dcifimemload_15),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~1 .lut_mask = 16'hF000;
defparam \Mux0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N0
cycloneive_lcell_comb \Mux0~2 (
// Equation(s):
// \Mux0~2_combout  = (\Mux0~1_combout ) # ((!cuifRegDst_0 & ((cuifregT_4) # (Equal23))))

	.dataa(cuifregT_4),
	.datab(\cu_dut|cuif.RegDst[0]~0_combout ),
	.datac(\cu_dut|Equal2~9_combout ),
	.datad(\Mux0~1_combout ),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~2 .lut_mask = 16'hFF32;
defparam \Mux0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N10
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// \Mux1~0_combout  = (dcifimemload_14 & (!Equal0 & ((!Equal22) # (!Equal21))))

	.dataa(dcifimemload_14),
	.datab(\cu_dut|Equal0~0_combout ),
	.datac(\cu_dut|Equal2~7_combout ),
	.datad(\cu_dut|Equal2~8_combout ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'h0222;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N22
cycloneive_lcell_comb \Mux1~1 (
// Equation(s):
// \Mux1~1_combout  = (\Mux1~0_combout ) # ((!cuifRegDst_0 & ((cuifregT_3) # (Equal23))))

	.dataa(\Mux1~0_combout ),
	.datab(\cu_dut|cuif.regT[3]~2_combout ),
	.datac(\cu_dut|Equal2~9_combout ),
	.datad(\cu_dut|cuif.RegDst[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~1 .lut_mask = 16'hAAFE;
defparam \Mux1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N22
cycloneive_lcell_comb \WEN~2 (
// Equation(s):
// \WEN~2_combout  = (dcifimemload_5 & (((!dcifimemload_2 & dcifimemload_1)) # (!dcifimemload_3)))

	.dataa(dcifimemload_5),
	.datab(dcifimemload_3),
	.datac(dcifimemload_2),
	.datad(dcifimemload_1),
	.cin(gnd),
	.combout(\WEN~2_combout ),
	.cout());
// synopsys translate_off
defparam \WEN~2 .lut_mask = 16'h2A22;
defparam \WEN~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N8
cycloneive_lcell_comb \WEN~3 (
// Equation(s):
// \WEN~3_combout  = (dcifimemload_29) # ((cuifaluOp_3 & ((WideOr4) # (\WEN~2_combout ))))

	.dataa(\cu_dut|WideOr4~2_combout ),
	.datab(\cu_dut|cuif.aluOp[3]~1_combout ),
	.datac(dcifimemload_29),
	.datad(\WEN~2_combout ),
	.cin(gnd),
	.combout(\WEN~3_combout ),
	.cout());
// synopsys translate_off
defparam \WEN~3 .lut_mask = 16'hFCF8;
defparam \WEN~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N10
cycloneive_lcell_comb \WEN~4 (
// Equation(s):
// \WEN~4_combout  = (dcifimemload_31 & (Equal21 & ((\WEN~6_combout )))) # (!dcifimemload_31 & ((Equal21) # ((\WEN~3_combout ))))

	.dataa(dcifimemload_31),
	.datab(\cu_dut|Equal2~7_combout ),
	.datac(\WEN~3_combout ),
	.datad(\WEN~6_combout ),
	.cin(gnd),
	.combout(\WEN~4_combout ),
	.cout());
// synopsys translate_off
defparam \WEN~4 .lut_mask = 16'hDC54;
defparam \WEN~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N12
cycloneive_lcell_comb \WEN~5 (
// Equation(s):
// \WEN~5_combout  = (dcifimemload_30 & (dcifimemload_31 & (Equal12))) # (!dcifimemload_30 & (((\WEN~4_combout ))))

	.dataa(dcifimemload_30),
	.datab(dcifimemload_31),
	.datac(\cu_dut|Equal12~2_combout ),
	.datad(\WEN~4_combout ),
	.cin(gnd),
	.combout(\WEN~5_combout ),
	.cout());
// synopsys translate_off
defparam \WEN~5 .lut_mask = 16'hD580;
defparam \WEN~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N28
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (\Mux0~0_combout  & dcifimemload_12)

	.dataa(gnd),
	.datab(gnd),
	.datac(\Mux0~0_combout ),
	.datad(dcifimemload_12),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hF000;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N30
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// \Mux3~1_combout  = (\Mux3~0_combout ) # ((!cuifRegDst_0 & ((cuifregT_1) # (Equal23))))

	.dataa(\Mux3~0_combout ),
	.datab(\cu_dut|cuif.regT[1]~5_combout ),
	.datac(\cu_dut|Equal2~9_combout ),
	.datad(\cu_dut|cuif.RegDst[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'hAAFE;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N28
cycloneive_lcell_comb \Mux37~0 (
// Equation(s):
// \Mux37~0_combout  = (cuifMemtoReg_0 & (((cuifMemtoReg_1)))) # (!cuifMemtoReg_0 & ((cuifMemtoReg_1 & (dcifimemload_15)) # (!cuifMemtoReg_1 & ((Selector0)))))

	.dataa(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datab(dcifimemload_15),
	.datac(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datad(Selector0),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~0 .lut_mask = 16'hE5E0;
defparam \Mux37~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N26
cycloneive_lcell_comb \Mux37~1 (
// Equation(s):
// \Mux37~1_combout  = (cuifMemtoReg_0 & ((\Mux37~0_combout  & (\Add0~58_combout )) # (!\Mux37~0_combout  & ((ramiframload_311))))) # (!cuifMemtoReg_0 & (((\Mux37~0_combout ))))

	.dataa(\Add0~58_combout ),
	.datab(ramiframload_311),
	.datac(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\Mux37~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~1 .lut_mask = 16'hAFC0;
defparam \Mux37~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N18
cycloneive_lcell_comb \Mux38~0 (
// Equation(s):
// \Mux38~0_combout  = (cuifMemtoReg_0 & ((ramiframload_301) # ((cuifMemtoReg_1)))) # (!cuifMemtoReg_0 & (((!cuifMemtoReg_1 & Selector1))))

	.dataa(ramiframload_301),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datad(Selector1),
	.cin(gnd),
	.combout(\Mux38~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~0 .lut_mask = 16'hCBC8;
defparam \Mux38~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N24
cycloneive_lcell_comb \Mux38~1 (
// Equation(s):
// \Mux38~1_combout  = (\Mux38~0_combout  & ((\Add0~56_combout ) # ((!cuifMemtoReg_1)))) # (!\Mux38~0_combout  & (((dcifimemload_14 & cuifMemtoReg_1))))

	.dataa(\Add0~56_combout ),
	.datab(\Mux38~0_combout ),
	.datac(dcifimemload_14),
	.datad(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.cin(gnd),
	.combout(\Mux38~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~1 .lut_mask = 16'hB8CC;
defparam \Mux38~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N30
cycloneive_lcell_comb \Mux39~0 (
// Equation(s):
// \Mux39~0_combout  = (cuifMemtoReg_1 & ((dcifimemload_13) # ((cuifMemtoReg_0)))) # (!cuifMemtoReg_1 & (((!cuifMemtoReg_0 & Selector2))))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(dcifimemload_13),
	.datac(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datad(Selector2),
	.cin(gnd),
	.combout(\Mux39~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~0 .lut_mask = 16'hADA8;
defparam \Mux39~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N2
cycloneive_lcell_comb \Mux39~1 (
// Equation(s):
// \Mux39~1_combout  = (cuifMemtoReg_0 & ((\Mux39~0_combout  & ((\Add0~54_combout ))) # (!\Mux39~0_combout  & (ramiframload_291)))) # (!cuifMemtoReg_0 & (((\Mux39~0_combout ))))

	.dataa(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datab(ramiframload_291),
	.datac(\Mux39~0_combout ),
	.datad(\Add0~54_combout ),
	.cin(gnd),
	.combout(\Mux39~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~1 .lut_mask = 16'hF858;
defparam \Mux39~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N14
cycloneive_lcell_comb \Mux40~0 (
// Equation(s):
// \Mux40~0_combout  = (cuifMemtoReg_0 & ((ramiframload_281) # ((cuifMemtoReg_1)))) # (!cuifMemtoReg_0 & (((!cuifMemtoReg_1 & Selector3))))

	.dataa(ramiframload_281),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datad(Selector3),
	.cin(gnd),
	.combout(\Mux40~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~0 .lut_mask = 16'hCBC8;
defparam \Mux40~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N12
cycloneive_lcell_comb \Mux40~1 (
// Equation(s):
// \Mux40~1_combout  = (cuifMemtoReg_1 & ((\Mux40~0_combout  & (\Add0~52_combout )) # (!\Mux40~0_combout  & ((dcifimemload_12))))) # (!cuifMemtoReg_1 & (((\Mux40~0_combout ))))

	.dataa(\Add0~52_combout ),
	.datab(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datac(dcifimemload_12),
	.datad(\Mux40~0_combout ),
	.cin(gnd),
	.combout(\Mux40~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~1 .lut_mask = 16'hBBC0;
defparam \Mux40~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N14
cycloneive_lcell_comb \Mux41~0 (
// Equation(s):
// \Mux41~0_combout  = (cuifMemtoReg_1 & ((dcifimemload_11) # ((cuifMemtoReg_0)))) # (!cuifMemtoReg_1 & (((Selector41 & !cuifMemtoReg_0))))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(dcifimemload_11),
	.datac(Selector41),
	.datad(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.cin(gnd),
	.combout(\Mux41~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~0 .lut_mask = 16'hAAD8;
defparam \Mux41~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N18
cycloneive_lcell_comb \Mux41~1 (
// Equation(s):
// \Mux41~1_combout  = (cuifMemtoReg_0 & ((\Mux41~0_combout  & ((\Add0~50_combout ))) # (!\Mux41~0_combout  & (ramiframload_271)))) # (!cuifMemtoReg_0 & (((\Mux41~0_combout ))))

	.dataa(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datab(ramiframload_271),
	.datac(\Add0~50_combout ),
	.datad(\Mux41~0_combout ),
	.cin(gnd),
	.combout(\Mux41~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~1 .lut_mask = 16'hF588;
defparam \Mux41~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N16
cycloneive_lcell_comb \Mux42~0 (
// Equation(s):
// \Mux42~0_combout  = (cuifMemtoReg_1 & (((cuifMemtoReg_0)))) # (!cuifMemtoReg_1 & ((cuifMemtoReg_0 & (ramiframload_261)) # (!cuifMemtoReg_0 & ((Selector5)))))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(ramiframload_261),
	.datac(Selector5),
	.datad(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.cin(gnd),
	.combout(\Mux42~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~0 .lut_mask = 16'hEE50;
defparam \Mux42~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N2
cycloneive_lcell_comb \Mux42~1 (
// Equation(s):
// \Mux42~1_combout  = (cuifMemtoReg_1 & ((\Mux42~0_combout  & (\Add0~48_combout )) # (!\Mux42~0_combout  & ((dcifimemload_10))))) # (!cuifMemtoReg_1 & (((\Mux42~0_combout ))))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(\Add0~48_combout ),
	.datac(dcifimemload_10),
	.datad(\Mux42~0_combout ),
	.cin(gnd),
	.combout(\Mux42~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~1 .lut_mask = 16'hDDA0;
defparam \Mux42~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N30
cycloneive_lcell_comb \Mux43~0 (
// Equation(s):
// \Mux43~0_combout  = (cuifMemtoReg_1 & ((cuifMemtoReg_0) # ((dcifimemload_9)))) # (!cuifMemtoReg_1 & (!cuifMemtoReg_0 & ((Selector6))))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(dcifimemload_9),
	.datad(Selector6),
	.cin(gnd),
	.combout(\Mux43~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~0 .lut_mask = 16'hB9A8;
defparam \Mux43~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N24
cycloneive_lcell_comb \Mux43~1 (
// Equation(s):
// \Mux43~1_combout  = (\Mux43~0_combout  & ((\Add0~46_combout ) # ((!cuifMemtoReg_0)))) # (!\Mux43~0_combout  & (((ramiframload_25 & cuifMemtoReg_0))))

	.dataa(\Add0~46_combout ),
	.datab(ramiframload_25),
	.datac(\Mux43~0_combout ),
	.datad(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.cin(gnd),
	.combout(\Mux43~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~1 .lut_mask = 16'hACF0;
defparam \Mux43~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N4
cycloneive_lcell_comb \Mux44~0 (
// Equation(s):
// \Mux44~0_combout  = (cuifMemtoReg_1 & (cuifMemtoReg_0)) # (!cuifMemtoReg_1 & ((cuifMemtoReg_0 & (ramiframload_24)) # (!cuifMemtoReg_0 & ((Selector71)))))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(ramiframload_24),
	.datad(\alu_dut|Selector7~8_combout ),
	.cin(gnd),
	.combout(\Mux44~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~0 .lut_mask = 16'hD9C8;
defparam \Mux44~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N30
cycloneive_lcell_comb \Mux44~1 (
// Equation(s):
// \Mux44~1_combout  = (\Mux44~0_combout  & (((\Add0~44_combout ) # (!cuifMemtoReg_1)))) # (!\Mux44~0_combout  & (dcifimemload_8 & ((cuifMemtoReg_1))))

	.dataa(dcifimemload_8),
	.datab(\Add0~44_combout ),
	.datac(\Mux44~0_combout ),
	.datad(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.cin(gnd),
	.combout(\Mux44~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~1 .lut_mask = 16'hCAF0;
defparam \Mux44~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N26
cycloneive_lcell_comb \Mux45~0 (
// Equation(s):
// \Mux45~0_combout  = (cuifMemtoReg_1 & ((dcifimemload_7) # ((cuifMemtoReg_0)))) # (!cuifMemtoReg_1 & (((!cuifMemtoReg_0 & Selector83))))

	.dataa(dcifimemload_7),
	.datab(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datac(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datad(\alu_dut|Selector8~11_combout ),
	.cin(gnd),
	.combout(\Mux45~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~0 .lut_mask = 16'hCBC8;
defparam \Mux45~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N8
cycloneive_lcell_comb \Mux45~1 (
// Equation(s):
// \Mux45~1_combout  = (cuifMemtoReg_0 & ((\Mux45~0_combout  & (\Add0~42_combout )) # (!\Mux45~0_combout  & ((ramiframload_23))))) # (!cuifMemtoReg_0 & (((\Mux45~0_combout ))))

	.dataa(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datab(\Add0~42_combout ),
	.datac(\Mux45~0_combout ),
	.datad(ramiframload_23),
	.cin(gnd),
	.combout(\Mux45~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~1 .lut_mask = 16'hDAD0;
defparam \Mux45~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N22
cycloneive_lcell_comb \Mux46~0 (
// Equation(s):
// \Mux46~0_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1) # ((ramiframload_22)))) # (!cuifMemtoReg_0 & (!cuifMemtoReg_1 & ((Selector9))))

	.dataa(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datab(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datac(ramiframload_22),
	.datad(Selector9),
	.cin(gnd),
	.combout(\Mux46~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~0 .lut_mask = 16'hB9A8;
defparam \Mux46~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N20
cycloneive_lcell_comb \Mux46~1 (
// Equation(s):
// \Mux46~1_combout  = (\Mux46~0_combout  & (((\Add0~40_combout ) # (!cuifMemtoReg_1)))) # (!\Mux46~0_combout  & (dcifimemload_6 & ((cuifMemtoReg_1))))

	.dataa(dcifimemload_6),
	.datab(\Add0~40_combout ),
	.datac(\Mux46~0_combout ),
	.datad(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.cin(gnd),
	.combout(\Mux46~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~1 .lut_mask = 16'hCAF0;
defparam \Mux46~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N8
cycloneive_lcell_comb \Mux47~0 (
// Equation(s):
// \Mux47~0_combout  = (cuifMemtoReg_0 & (((cuifMemtoReg_1)))) # (!cuifMemtoReg_0 & ((cuifMemtoReg_1 & (dcifimemload_5)) # (!cuifMemtoReg_1 & ((Selector10)))))

	.dataa(dcifimemload_5),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(Selector10),
	.datad(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.cin(gnd),
	.combout(\Mux47~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~0 .lut_mask = 16'hEE30;
defparam \Mux47~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N6
cycloneive_lcell_comb \Mux47~1 (
// Equation(s):
// \Mux47~1_combout  = (cuifMemtoReg_0 & ((\Mux47~0_combout  & (\Add0~38_combout )) # (!\Mux47~0_combout  & ((ramiframload_21))))) # (!cuifMemtoReg_0 & (((\Mux47~0_combout ))))

	.dataa(\Add0~38_combout ),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(\Mux47~0_combout ),
	.datad(ramiframload_21),
	.cin(gnd),
	.combout(\Mux47~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~1 .lut_mask = 16'hBCB0;
defparam \Mux47~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N20
cycloneive_lcell_comb \Mux48~0 (
// Equation(s):
// \Mux48~0_combout  = (cuifMemtoReg_0 & ((ramiframload_20) # ((cuifMemtoReg_1)))) # (!cuifMemtoReg_0 & (((!cuifMemtoReg_1 & Selector11))))

	.dataa(ramiframload_20),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datad(Selector11),
	.cin(gnd),
	.combout(\Mux48~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~0 .lut_mask = 16'hCBC8;
defparam \Mux48~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N30
cycloneive_lcell_comb \Mux48~1 (
// Equation(s):
// \Mux48~1_combout  = (cuifMemtoReg_1 & ((\Mux48~0_combout  & ((\Add0~36_combout ))) # (!\Mux48~0_combout  & (dcifimemload_4)))) # (!cuifMemtoReg_1 & (((\Mux48~0_combout ))))

	.dataa(dcifimemload_4),
	.datab(\Add0~36_combout ),
	.datac(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datad(\Mux48~0_combout ),
	.cin(gnd),
	.combout(\Mux48~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~1 .lut_mask = 16'hCFA0;
defparam \Mux48~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N22
cycloneive_lcell_comb \Mux63~0 (
// Equation(s):
// \Mux63~0_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & (\Add0~6_combout )) # (!cuifMemtoReg_1 & ((ramiframload_5)))))

	.dataa(\Add0~6_combout ),
	.datab(ramiframload_5),
	.datac(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datad(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.cin(gnd),
	.combout(\Mux63~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~0 .lut_mask = 16'hAC00;
defparam \Mux63~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N8
cycloneive_lcell_comb \Mux63~1 (
// Equation(s):
// \Mux63~1_combout  = (\Mux63~0_combout ) # ((Selector261 & (!cuifMemtoReg_1 & !cuifMemtoReg_0)))

	.dataa(\alu_dut|Selector26~7_combout ),
	.datab(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datac(\Mux63~0_combout ),
	.datad(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.cin(gnd),
	.combout(\Mux63~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~1 .lut_mask = 16'hF0F2;
defparam \Mux63~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N22
cycloneive_lcell_comb \Mux49~0 (
// Equation(s):
// \Mux49~0_combout  = (cuifMemtoReg_1 & ((cuifMemtoReg_0) # ((dcifimemload_3)))) # (!cuifMemtoReg_1 & (!cuifMemtoReg_0 & ((Selector12))))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(dcifimemload_3),
	.datad(Selector12),
	.cin(gnd),
	.combout(\Mux49~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~0 .lut_mask = 16'hB9A8;
defparam \Mux49~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N24
cycloneive_lcell_comb \Mux49~1 (
// Equation(s):
// \Mux49~1_combout  = (\Mux49~0_combout  & (((\Add0~34_combout ) # (!cuifMemtoReg_0)))) # (!\Mux49~0_combout  & (ramiframload_19 & ((cuifMemtoReg_0))))

	.dataa(ramiframload_19),
	.datab(\Add0~34_combout ),
	.datac(\Mux49~0_combout ),
	.datad(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.cin(gnd),
	.combout(\Mux49~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~1 .lut_mask = 16'hCAF0;
defparam \Mux49~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N18
cycloneive_lcell_comb \Mux50~0 (
// Equation(s):
// \Mux50~0_combout  = (cuifMemtoReg_0 & ((ramiframload_18) # ((cuifMemtoReg_1)))) # (!cuifMemtoReg_0 & (((Selector13 & !cuifMemtoReg_1))))

	.dataa(ramiframload_18),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(Selector13),
	.datad(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.cin(gnd),
	.combout(\Mux50~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~0 .lut_mask = 16'hCCB8;
defparam \Mux50~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N4
cycloneive_lcell_comb \Mux50~1 (
// Equation(s):
// \Mux50~1_combout  = (cuifMemtoReg_1 & ((\Mux50~0_combout  & ((\Add0~32_combout ))) # (!\Mux50~0_combout  & (dcifimemload_2)))) # (!cuifMemtoReg_1 & (((\Mux50~0_combout ))))

	.dataa(dcifimemload_2),
	.datab(\Add0~32_combout ),
	.datac(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datad(\Mux50~0_combout ),
	.cin(gnd),
	.combout(\Mux50~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~1 .lut_mask = 16'hCFA0;
defparam \Mux50~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N8
cycloneive_lcell_comb \Mux51~0 (
// Equation(s):
// \Mux51~0_combout  = (cuifMemtoReg_1 & ((dcifimemload_1) # ((cuifMemtoReg_0)))) # (!cuifMemtoReg_1 & (((Selector14 & !cuifMemtoReg_0))))

	.dataa(dcifimemload_1),
	.datab(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datac(Selector14),
	.datad(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.cin(gnd),
	.combout(\Mux51~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~0 .lut_mask = 16'hCCB8;
defparam \Mux51~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N30
cycloneive_lcell_comb \Mux51~1 (
// Equation(s):
// \Mux51~1_combout  = (\Mux51~0_combout  & ((\Add0~30_combout ) # ((!cuifMemtoReg_0)))) # (!\Mux51~0_combout  & (((ramiframload_17 & cuifMemtoReg_0))))

	.dataa(\Add0~30_combout ),
	.datab(ramiframload_17),
	.datac(\Mux51~0_combout ),
	.datad(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.cin(gnd),
	.combout(\Mux51~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~1 .lut_mask = 16'hACF0;
defparam \Mux51~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N14
cycloneive_lcell_comb \Mux52~0 (
// Equation(s):
// \Mux52~0_combout  = (cuifMemtoReg_0 & ((ramiframload_16) # ((cuifMemtoReg_1)))) # (!cuifMemtoReg_0 & (((!cuifMemtoReg_1 & Selector15))))

	.dataa(ramiframload_16),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datad(Selector15),
	.cin(gnd),
	.combout(\Mux52~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~0 .lut_mask = 16'hCBC8;
defparam \Mux52~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N14
cycloneive_lcell_comb \Mux52~1 (
// Equation(s):
// \Mux52~1_combout  = (cuifMemtoReg_1 & ((\Mux52~0_combout  & ((\Add0~28_combout ))) # (!\Mux52~0_combout  & (dcifimemload_0)))) # (!cuifMemtoReg_1 & (((\Mux52~0_combout ))))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(dcifimemload_0),
	.datac(\Mux52~0_combout ),
	.datad(\Add0~28_combout ),
	.cin(gnd),
	.combout(\Mux52~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~1 .lut_mask = 16'hF858;
defparam \Mux52~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N24
cycloneive_lcell_comb \Mux53~0 (
// Equation(s):
// \Mux53~0_combout  = (cuifMemtoReg_1 & ((\Add0~26_combout ))) # (!cuifMemtoReg_1 & (ramiframload_15))

	.dataa(gnd),
	.datab(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datac(ramiframload_15),
	.datad(\Add0~26_combout ),
	.cin(gnd),
	.combout(\Mux53~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~0 .lut_mask = 16'hFC30;
defparam \Mux53~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N10
cycloneive_lcell_comb \Mux53~1 (
// Equation(s):
// \Mux53~1_combout  = (cuifMemtoReg_0 & (\Mux53~0_combout )) # (!cuifMemtoReg_0 & (((Selector16 & !cuifMemtoReg_1))))

	.dataa(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datab(\Mux53~0_combout ),
	.datac(Selector16),
	.datad(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.cin(gnd),
	.combout(\Mux53~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~1 .lut_mask = 16'h88D8;
defparam \Mux53~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N4
cycloneive_lcell_comb \Mux54~0 (
// Equation(s):
// \Mux54~0_combout  = (cuifMemtoReg_1 & (\Add0~24_combout )) # (!cuifMemtoReg_1 & ((ramiframload_14)))

	.dataa(\Add0~24_combout ),
	.datab(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datac(gnd),
	.datad(ramiframload_14),
	.cin(gnd),
	.combout(\Mux54~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~0 .lut_mask = 16'hBB88;
defparam \Mux54~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N6
cycloneive_lcell_comb \Mux54~1 (
// Equation(s):
// \Mux54~1_combout  = (cuifMemtoReg_0 & (((\Mux54~0_combout )))) # (!cuifMemtoReg_0 & (Selector17 & (!cuifMemtoReg_1)))

	.dataa(Selector17),
	.datab(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datac(\Mux54~0_combout ),
	.datad(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.cin(gnd),
	.combout(\Mux54~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~1 .lut_mask = 16'hF022;
defparam \Mux54~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N20
cycloneive_lcell_comb \Mux55~0 (
// Equation(s):
// \Mux55~0_combout  = (cuifMemtoReg_1 & (\Add0~22_combout )) # (!cuifMemtoReg_1 & ((ramiframload_13)))

	.dataa(\Add0~22_combout ),
	.datab(ramiframload_13),
	.datac(gnd),
	.datad(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.cin(gnd),
	.combout(\Mux55~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~0 .lut_mask = 16'hAACC;
defparam \Mux55~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N24
cycloneive_lcell_comb \Mux55~1 (
// Equation(s):
// \Mux55~1_combout  = (cuifMemtoReg_0 & (((\Mux55~0_combout )))) # (!cuifMemtoReg_0 & (Selector18 & (!cuifMemtoReg_1)))

	.dataa(Selector18),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datad(\Mux55~0_combout ),
	.cin(gnd),
	.combout(\Mux55~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~1 .lut_mask = 16'hCE02;
defparam \Mux55~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N14
cycloneive_lcell_comb \Mux56~0 (
// Equation(s):
// \Mux56~0_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & ((\Add0~20_combout ))) # (!cuifMemtoReg_1 & (ramiframload_12))))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(ramiframload_12),
	.datac(\Add0~20_combout ),
	.datad(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.cin(gnd),
	.combout(\Mux56~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~0 .lut_mask = 16'hE400;
defparam \Mux56~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N24
cycloneive_lcell_comb \Mux56~1 (
// Equation(s):
// \Mux56~1_combout  = (\Mux56~0_combout ) # ((!cuifMemtoReg_1 & (!cuifMemtoReg_0 & Selector19)))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(\Mux56~0_combout ),
	.datad(Selector19),
	.cin(gnd),
	.combout(\Mux56~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~1 .lut_mask = 16'hF1F0;
defparam \Mux56~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y35_N14
cycloneive_lcell_comb \Mux57~0 (
// Equation(s):
// \Mux57~0_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & ((\Add0~18_combout ))) # (!cuifMemtoReg_1 & (ramiframload_11))))

	.dataa(ramiframload_11),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datad(\Add0~18_combout ),
	.cin(gnd),
	.combout(\Mux57~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~0 .lut_mask = 16'hC808;
defparam \Mux57~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N30
cycloneive_lcell_comb \Mux57~1 (
// Equation(s):
// \Mux57~1_combout  = (\Mux57~0_combout ) # ((!cuifMemtoReg_1 & (!cuifMemtoReg_0 & Selector20)))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(\Mux57~0_combout ),
	.datad(Selector20),
	.cin(gnd),
	.combout(\Mux57~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~1 .lut_mask = 16'hF1F0;
defparam \Mux57~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y34_N0
cycloneive_lcell_comb \Mux58~0 (
// Equation(s):
// \Mux58~0_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & ((\Add0~16_combout ))) # (!cuifMemtoReg_1 & (ramiframload_10))))

	.dataa(ramiframload_10),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datad(\Add0~16_combout ),
	.cin(gnd),
	.combout(\Mux58~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~0 .lut_mask = 16'hC808;
defparam \Mux58~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N16
cycloneive_lcell_comb \Mux58~1 (
// Equation(s):
// \Mux58~1_combout  = (\Mux58~0_combout ) # ((!cuifMemtoReg_1 & (!cuifMemtoReg_0 & Selector21)))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(\Mux58~0_combout ),
	.datad(Selector21),
	.cin(gnd),
	.combout(\Mux58~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~1 .lut_mask = 16'hF1F0;
defparam \Mux58~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N10
cycloneive_lcell_comb \Mux59~0 (
// Equation(s):
// \Mux59~0_combout  = (cuifMemtoReg_1 & (\Add0~14_combout )) # (!cuifMemtoReg_1 & ((ramiframload_9)))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(\Add0~14_combout ),
	.datac(gnd),
	.datad(ramiframload_9),
	.cin(gnd),
	.combout(\Mux59~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~0 .lut_mask = 16'hDD88;
defparam \Mux59~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N20
cycloneive_lcell_comb \Mux59~1 (
// Equation(s):
// \Mux59~1_combout  = (cuifMemtoReg_0 & (((\Mux59~0_combout )))) # (!cuifMemtoReg_0 & (!cuifMemtoReg_1 & ((Selector22))))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(\Mux59~0_combout ),
	.datac(Selector22),
	.datad(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.cin(gnd),
	.combout(\Mux59~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~1 .lut_mask = 16'hCC50;
defparam \Mux59~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N4
cycloneive_lcell_comb \Mux60~0 (
// Equation(s):
// \Mux60~0_combout  = (cuifMemtoReg_1 & ((\Add0~12_combout ))) # (!cuifMemtoReg_1 & (ramiframload_8))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(ramiframload_8),
	.datac(gnd),
	.datad(\Add0~12_combout ),
	.cin(gnd),
	.combout(\Mux60~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~0 .lut_mask = 16'hEE44;
defparam \Mux60~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N24
cycloneive_lcell_comb \Mux60~1 (
// Equation(s):
// \Mux60~1_combout  = (cuifMemtoReg_0 & (((\Mux60~0_combout )))) # (!cuifMemtoReg_0 & (!cuifMemtoReg_1 & (Selector23)))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(Selector23),
	.datac(\Mux60~0_combout ),
	.datad(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.cin(gnd),
	.combout(\Mux60~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~1 .lut_mask = 16'hF044;
defparam \Mux60~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N18
cycloneive_lcell_comb \Mux61~0 (
// Equation(s):
// \Mux61~0_combout  = (cuifMemtoReg_1 & ((\Add0~10_combout ))) # (!cuifMemtoReg_1 & (ramiframload_7))

	.dataa(ramiframload_7),
	.datab(\Add0~10_combout ),
	.datac(gnd),
	.datad(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.cin(gnd),
	.combout(\Mux61~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~0 .lut_mask = 16'hCCAA;
defparam \Mux61~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N20
cycloneive_lcell_comb \Mux61~1 (
// Equation(s):
// \Mux61~1_combout  = (cuifMemtoReg_0 & (\Mux61~0_combout )) # (!cuifMemtoReg_0 & (((!cuifMemtoReg_1 & Selector242))))

	.dataa(\Mux61~0_combout ),
	.datab(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datac(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datad(\alu_dut|Selector24~9_combout ),
	.cin(gnd),
	.combout(\Mux61~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~1 .lut_mask = 16'hA3A0;
defparam \Mux61~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N4
cycloneive_lcell_comb \Mux62~0 (
// Equation(s):
// \Mux62~0_combout  = (cuifMemtoReg_1 & (\Add0~8_combout )) # (!cuifMemtoReg_1 & ((ramiframload_6)))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(\Add0~8_combout ),
	.datac(gnd),
	.datad(ramiframload_6),
	.cin(gnd),
	.combout(\Mux62~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~0 .lut_mask = 16'hDD88;
defparam \Mux62~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N14
cycloneive_lcell_comb \Mux62~1 (
// Equation(s):
// \Mux62~1_combout  = (cuifMemtoReg_0 & (((\Mux62~0_combout )))) # (!cuifMemtoReg_0 & (!cuifMemtoReg_1 & ((Selector251))))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(\Mux62~0_combout ),
	.datad(\alu_dut|Selector25~7_combout ),
	.cin(gnd),
	.combout(\Mux62~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~1 .lut_mask = 16'hD1C0;
defparam \Mux62~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N10
cycloneive_lcell_comb \Mux66~0 (
// Equation(s):
// \Mux66~0_combout  = (cuifMemtoReg_1 & (\Add0~0_combout )) # (!cuifMemtoReg_1 & ((ramiframload_2)))

	.dataa(\Add0~0_combout ),
	.datab(ramiframload_2),
	.datac(gnd),
	.datad(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.cin(gnd),
	.combout(\Mux66~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux66~0 .lut_mask = 16'hAACC;
defparam \Mux66~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N2
cycloneive_lcell_comb \Mux66~1 (
// Equation(s):
// \Mux66~1_combout  = (cuifMemtoReg_0 & (((\Mux66~0_combout )))) # (!cuifMemtoReg_0 & (!cuifMemtoReg_1 & ((Selector29))))

	.dataa(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datab(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datac(\Mux66~0_combout ),
	.datad(Selector29),
	.cin(gnd),
	.combout(\Mux66~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux66~1 .lut_mask = 16'hB1A0;
defparam \Mux66~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N10
cycloneive_lcell_comb \Mux67~0 (
// Equation(s):
// \Mux67~0_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & (pcifimemaddr_1)) # (!cuifMemtoReg_1 & ((ramiframload_1)))))

	.dataa(pcifimemaddr_1),
	.datab(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datac(ramiframload_1),
	.datad(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.cin(gnd),
	.combout(\Mux67~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux67~0 .lut_mask = 16'hB800;
defparam \Mux67~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N16
cycloneive_lcell_comb \Mux67~1 (
// Equation(s):
// \Mux67~1_combout  = (\Mux67~0_combout ) # ((!cuifMemtoReg_1 & (Selector30 & !cuifMemtoReg_0)))

	.dataa(\Mux67~0_combout ),
	.datab(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datac(Selector30),
	.datad(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.cin(gnd),
	.combout(\Mux67~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux67~1 .lut_mask = 16'hAABA;
defparam \Mux67~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N2
cycloneive_lcell_comb \Mux64~0 (
// Equation(s):
// \Mux64~0_combout  = (cuifMemtoReg_0 & ((cuifMemtoReg_1 & ((\Add0~4_combout ))) # (!cuifMemtoReg_1 & (ramiframload_4))))

	.dataa(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datab(ramiframload_4),
	.datac(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datad(\Add0~4_combout ),
	.cin(gnd),
	.combout(\Mux64~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux64~0 .lut_mask = 16'hA808;
defparam \Mux64~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N16
cycloneive_lcell_comb \Mux64~1 (
// Equation(s):
// \Mux64~1_combout  = (\Mux64~0_combout ) # ((!cuifMemtoReg_0 & (!cuifMemtoReg_1 & Selector271)))

	.dataa(\Mux64~0_combout ),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datad(\alu_dut|Selector27~8_combout ),
	.cin(gnd),
	.combout(\Mux64~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux64~1 .lut_mask = 16'hABAA;
defparam \Mux64~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y33_N14
cycloneive_lcell_comb \Mux65~0 (
// Equation(s):
// \Mux65~0_combout  = (cuifMemtoReg_1 & ((\Add0~2_combout ))) # (!cuifMemtoReg_1 & (ramiframload_3))

	.dataa(gnd),
	.datab(ramiframload_3),
	.datac(\Add0~2_combout ),
	.datad(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.cin(gnd),
	.combout(\Mux65~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux65~0 .lut_mask = 16'hF0CC;
defparam \Mux65~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N20
cycloneive_lcell_comb \Mux65~1 (
// Equation(s):
// \Mux65~1_combout  = (cuifMemtoReg_0 & (((\Mux65~0_combout )))) # (!cuifMemtoReg_0 & (!cuifMemtoReg_1 & (Selector28)))

	.dataa(\cu_dut|cuif.MemtoReg[1]~2_combout ),
	.datab(\cu_dut|cuif.MemtoReg[0]~4_combout ),
	.datac(Selector28),
	.datad(\Mux65~0_combout ),
	.cin(gnd),
	.combout(\Mux65~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux65~1 .lut_mask = 16'hDC10;
defparam \Mux65~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N8
cycloneive_lcell_comb \Mux35~5 (
// Equation(s):
// \Mux35~5_combout  = (!cuifaluSrc_1 & ((Equal2 & (dcifimemload_29)) # (!Equal2 & ((!cuifregT_0)))))

	.dataa(dcifimemload_29),
	.datab(\cu_dut|cuif.regT[0]~1_combout ),
	.datac(\cu_dut|Equal2~4_combout ),
	.datad(\cu_dut|cuif.aluSrc[1]~1_combout ),
	.cin(gnd),
	.combout(\Mux35~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~5 .lut_mask = 16'h00A3;
defparam \Mux35~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N22
cycloneive_lcell_comb \Mux34~4 (
// Equation(s):
// \Mux34~4_combout  = (cuifregT_4 & (!cuifaluSrc_1 & (Mux61 & !cuifaluSrc_0)))

	.dataa(cuifregT_4),
	.datab(\cu_dut|cuif.aluSrc[1]~1_combout ),
	.datac(Mux61),
	.datad(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.cin(gnd),
	.combout(\Mux34~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~4 .lut_mask = 16'h0020;
defparam \Mux34~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N26
cycloneive_lcell_comb \Mux33~4 (
// Equation(s):
// \Mux33~4_combout  = (!cuifaluSrc_0 & (cuifregT_4 & (!cuifaluSrc_1 & Mux60)))

	.dataa(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.datab(cuifregT_4),
	.datac(\cu_dut|cuif.aluSrc[1]~1_combout ),
	.datad(Mux60),
	.cin(gnd),
	.combout(\Mux33~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~4 .lut_mask = 16'h0400;
defparam \Mux33~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N22
cycloneive_lcell_comb \Mux32~5 (
// Equation(s):
// \Mux32~5_combout  = (!cuifaluSrc_0 & (!cuifaluSrc_1 & (cuifregT_4 & Mux59)))

	.dataa(\cu_dut|cuif.aluSrc[0]~0_combout ),
	.datab(\cu_dut|cuif.aluSrc[1]~1_combout ),
	.datac(cuifregT_4),
	.datad(Mux59),
	.cin(gnd),
	.combout(\Mux32~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~5 .lut_mask = 16'h1000;
defparam \Mux32~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N30
cycloneive_lcell_comb \WEN~6 (
// Equation(s):
// \WEN~6_combout  = (always1 & (!instr_29 & ((ruifdmemWEN) # (ruifdmemREN))))

	.dataa(always1),
	.datab(instr_29),
	.datac(ruifdmemWEN),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(\WEN~6_combout ),
	.cout());
// synopsys translate_off
defparam \WEN~6 .lut_mask = 16'h2220;
defparam \WEN~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: DDIOOUTCELL_X0_Y32_N18
dffeas \dpif.halt (
	.clk(CLK),
	.d(\dpif.halt~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dpifhalt),
	.prn(vcc));
// synopsys translate_off
defparam \dpif.halt .is_wysiwyg = "true";
defparam \dpif.halt .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N6
cycloneive_lcell_comb \dpif.halt~_Duplicate_1feeder (
// Equation(s):
// \dpif.halt~_Duplicate_1feeder_combout  = \dpif.halt~0_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\dpif.halt~0_combout ),
	.cin(gnd),
	.combout(\dpif.halt~_Duplicate_1feeder_combout ),
	.cout());
// synopsys translate_off
defparam \dpif.halt~_Duplicate_1feeder .lut_mask = 16'hFF00;
defparam \dpif.halt~_Duplicate_1feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y32_N7
dffeas \dpif.halt~_Duplicate_1 (
	.clk(CLK),
	.d(\dpif.halt~_Duplicate_1feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\dpif.halt~_Duplicate_1_q ),
	.prn(vcc));
// synopsys translate_off
defparam \dpif.halt~_Duplicate_1 .is_wysiwyg = "true";
defparam \dpif.halt~_Duplicate_1 .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N2
cycloneive_lcell_comb \dpif.halt~0 (
// Equation(s):
// \dpif.halt~0_combout  = (\dpif.halt~_Duplicate_1_q ) # ((dcifimemload_30 & (dcifimemload_31 & Equal12)))

	.dataa(dcifimemload_30),
	.datab(dcifimemload_31),
	.datac(\cu_dut|Equal12~2_combout ),
	.datad(\dpif.halt~_Duplicate_1_q ),
	.cin(gnd),
	.combout(\dpif.halt~0_combout ),
	.cout());
// synopsys translate_off
defparam \dpif.halt~0 .lut_mask = 16'hFF80;
defparam \dpif.halt~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module alu (
	cuifaluOp_3,
	cuifaluOp_2,
	cuifaluOp_1,
	cuifaluOp_0,
	Mux5,
	Mux51,
	Mux6,
	Mux7,
	Mux8,
	Mux9,
	Mux10,
	Mux11,
	Mux12,
	Mux13,
	Mux14,
	Mux15,
	Mux151,
	Mux16,
	Mux31,
	Mux17,
	Mux18,
	Mux19,
	Mux20,
	Mux21,
	Mux22,
	Mux23,
	Mux24,
	Mux25,
	Mux26,
	Mux27,
	Mux28,
	Mux29,
	Mux30,
	Mux291,
	Mux301,
	Mux36,
	Mux35,
	Mux351,
	Mux352,
	Mux271,
	Mux281,
	Mux34,
	Mux231,
	Mux241,
	Mux251,
	Mux261,
	Mux33,
	Mux152,
	Mux161,
	Mux171,
	Mux181,
	Mux191,
	Mux201,
	Mux211,
	Mux221,
	Mux32,
	Mux0,
	Mux2,
	Mux1,
	Mux3,
	Mux4,
	Mux52,
	Mux61,
	Mux71,
	Mux81,
	Mux91,
	Mux101,
	Mux111,
	Mux121,
	Mux131,
	Mux141,
	Mux311,
	Selector30,
	ShiftRight0,
	Mux53,
	Mux62,
	Mux82,
	Mux92,
	Mux102,
	Mux112,
	Mux132,
	Mux172,
	Mux182,
	Mux192,
	Selector31,
	Selector311,
	Selector28,
	ShiftLeft0,
	Selector0,
	ShiftLeft01,
	Selector2,
	Selector29,
	Selector4,
	Selector5,
	ShiftLeft02,
	Selector3,
	ShiftLeft03,
	Selector1,
	Selector41,
	Selector10,
	Selector6,
	Selector7,
	Selector71,
	Selector11,
	Selector24,
	Selector241,
	Selector242,
	Selector25,
	Selector251,
	Selector13,
	Selector12,
	Selector26,
	Selector261,
	Selector27,
	Selector271,
	Equal10,
	Selector14,
	Selector15,
	Selector16,
	Selector17,
	Equal101,
	Selector20,
	Selector21,
	Selector18,
	Selector19,
	Selector8,
	Selector81,
	Selector82,
	Selector9,
	Selector312,
	Selector22,
	Selector23,
	Equal102,
	Selector83,
	devpor,
	devclrn,
	devoe);
input 	cuifaluOp_3;
input 	cuifaluOp_2;
input 	cuifaluOp_1;
input 	cuifaluOp_0;
input 	Mux5;
input 	Mux51;
input 	Mux6;
input 	Mux7;
input 	Mux8;
input 	Mux9;
input 	Mux10;
input 	Mux11;
input 	Mux12;
input 	Mux13;
input 	Mux14;
input 	Mux15;
input 	Mux151;
input 	Mux16;
input 	Mux31;
input 	Mux17;
input 	Mux18;
input 	Mux19;
input 	Mux20;
input 	Mux21;
input 	Mux22;
input 	Mux23;
input 	Mux24;
input 	Mux25;
input 	Mux26;
input 	Mux27;
input 	Mux28;
input 	Mux29;
input 	Mux30;
input 	Mux291;
input 	Mux301;
input 	Mux36;
input 	Mux35;
input 	Mux351;
input 	Mux352;
input 	Mux271;
input 	Mux281;
input 	Mux34;
input 	Mux231;
input 	Mux241;
input 	Mux251;
input 	Mux261;
input 	Mux33;
input 	Mux152;
input 	Mux161;
input 	Mux171;
input 	Mux181;
input 	Mux191;
input 	Mux201;
input 	Mux211;
input 	Mux221;
input 	Mux32;
input 	Mux0;
input 	Mux2;
input 	Mux1;
input 	Mux3;
input 	Mux4;
input 	Mux52;
input 	Mux61;
input 	Mux71;
input 	Mux81;
input 	Mux91;
input 	Mux101;
input 	Mux111;
input 	Mux121;
input 	Mux131;
input 	Mux141;
input 	Mux311;
output 	Selector30;
output 	ShiftRight0;
input 	Mux53;
input 	Mux62;
input 	Mux82;
input 	Mux92;
input 	Mux102;
input 	Mux112;
input 	Mux132;
input 	Mux172;
input 	Mux182;
input 	Mux192;
output 	Selector31;
output 	Selector311;
output 	Selector28;
output 	ShiftLeft0;
output 	Selector0;
output 	ShiftLeft01;
output 	Selector2;
output 	Selector29;
output 	Selector4;
output 	Selector5;
output 	ShiftLeft02;
output 	Selector3;
output 	ShiftLeft03;
output 	Selector1;
output 	Selector41;
output 	Selector10;
output 	Selector6;
output 	Selector7;
output 	Selector71;
output 	Selector11;
output 	Selector24;
output 	Selector241;
output 	Selector242;
output 	Selector25;
output 	Selector251;
output 	Selector13;
output 	Selector12;
output 	Selector26;
output 	Selector261;
output 	Selector27;
output 	Selector271;
output 	Equal10;
output 	Selector14;
output 	Selector15;
output 	Selector16;
output 	Selector17;
output 	Equal101;
output 	Selector20;
output 	Selector21;
output 	Selector18;
output 	Selector19;
output 	Selector8;
output 	Selector81;
output 	Selector82;
output 	Selector9;
output 	Selector312;
output 	Selector22;
output 	Selector23;
output 	Equal102;
output 	Selector83;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add0~10_combout ;
wire \Add0~14_combout ;
wire \Add0~18_combout ;
wire \Add0~24_combout ;
wire \Add0~32_combout ;
wire \Add0~44_combout ;
wire \Add1~10_combout ;
wire \Add1~20_combout ;
wire \Add1~34_combout ;
wire \Add1~36_combout ;
wire \ShiftRight0~52_combout ;
wire \ShiftRight0~63_combout ;
wire \ShiftRight0~103_combout ;
wire \Selector31~2_combout ;
wire \Selector0~31_combout ;
wire \Selector2~6_combout ;
wire \ShiftLeft0~72_combout ;
wire \Selector29~2_combout ;
wire \Selector1~1_combout ;
wire \Selector4~1_combout ;
wire \Selector11~5_combout ;
wire \Selector11~6_combout ;
wire \Selector13~4_combout ;
wire \Selector12~3_combout ;
wire \Selector26~1_combout ;
wire \Selector14~3_combout ;
wire \Selector15~3_combout ;
wire \Selector20~3_combout ;
wire \Selector21~2_combout ;
wire \Selector18~1_combout ;
wire \Selector8~7_combout ;
wire \Selector9~5_combout ;
wire \Selector9~6_combout ;
wire \Selector23~2_combout ;
wire \Selector0~9_combout ;
wire \Selector30~3_combout ;
wire \Selector0~10_combout ;
wire \Selector30~4_combout ;
wire \Selector0~8_combout ;
wire \Selector0~12_combout ;
wire \Add1~1 ;
wire \Add1~2_combout ;
wire \Add0~1 ;
wire \Add0~2_combout ;
wire \Selector30~6_combout ;
wire \Selector0~11_combout ;
wire \Selector30~5_combout ;
wire \Selector30~7_combout ;
wire \ShiftRight0~71_combout ;
wire \ShiftRight0~70_combout ;
wire \ShiftRight0~130_combout ;
wire \ShiftRight0~68_combout ;
wire \ShiftRight0~69_combout ;
wire \ShiftRight0~129_combout ;
wire \ShiftRight0~72_combout ;
wire \ShiftRight0~62_combout ;
wire \ShiftRight0~64_combout ;
wire \ShiftRight0~66_combout ;
wire \ShiftRight0~65_combout ;
wire \ShiftRight0~128_combout ;
wire \ShiftRight0~67_combout ;
wire \ShiftRight0~73_combout ;
wire \ShiftRight0~77_combout ;
wire \ShiftRight0~76_combout ;
wire \ShiftRight0~131_combout ;
wire \ShiftRight0~74_combout ;
wire \ShiftRight0~75_combout ;
wire \ShiftRight0~78_combout ;
wire \ShiftRight0~79_combout ;
wire \ShiftRight0~80_combout ;
wire \ShiftRight0~132_combout ;
wire \ShiftRight0~82_combout ;
wire \ShiftRight0~133_combout ;
wire \Selector22~0_combout ;
wire \ShiftRight0~83_combout ;
wire \Selector0~6_combout ;
wire \Selector24~0_combout ;
wire \Selector30~0_combout ;
wire \ShiftLeft0~52_combout ;
wire \Selector30~1_combout ;
wire \Selector0~7_combout ;
wire \ShiftRight0~53_combout ;
wire \ShiftRight0~54_combout ;
wire \ShiftRight0~55_combout ;
wire \ShiftRight0~56_combout ;
wire \ShiftRight0~57_combout ;
wire \ShiftRight0~59_combout ;
wire \ShiftRight0~58_combout ;
wire \ShiftRight0~60_combout ;
wire \ShiftRight0~61_combout ;
wire \Selector30~2_combout ;
wire \ShiftRight0~96_combout ;
wire \ShiftRight0~97_combout ;
wire \ShiftRight0~137_combout ;
wire \ShiftRight0~98_combout ;
wire \ShiftRight0~99_combout ;
wire \ShiftRight0~138_combout ;
wire \ShiftRight0~90_combout ;
wire \ShiftRight0~91_combout ;
wire \ShiftRight0~135_combout ;
wire \ShiftRight0~93_combout ;
wire \ShiftRight0~92_combout ;
wire \ShiftRight0~136_combout ;
wire \ShiftRight0~94_combout ;
wire \ShiftRight0~88_combout ;
wire \ShiftRight0~87_combout ;
wire \ShiftRight0~134_combout ;
wire \ShiftRight0~85_combout ;
wire \ShiftRight0~84_combout ;
wire \ShiftRight0~86_combout ;
wire \ShiftRight0~89_combout ;
wire \ShiftRight0~95_combout ;
wire \ShiftRight0~102_combout ;
wire \ShiftRight0~101_combout ;
wire \ShiftRight0~139_combout ;
wire \ShiftRight0~104_combout ;
wire \ShiftRight0~140_combout ;
wire \Selector23~0_combout ;
wire \ShiftRight0~105_combout ;
wire \Selector31~0_combout ;
wire \Selector0~13_combout ;
wire \Add0~0_combout ;
wire \Selector31~1_combout ;
wire \Add1~0_combout ;
wire \LessThan1~1_cout ;
wire \LessThan1~3_cout ;
wire \LessThan1~5_cout ;
wire \LessThan1~7_cout ;
wire \LessThan1~9_cout ;
wire \LessThan1~11_cout ;
wire \LessThan1~13_cout ;
wire \LessThan1~15_cout ;
wire \LessThan1~17_cout ;
wire \LessThan1~19_cout ;
wire \LessThan1~21_cout ;
wire \LessThan1~23_cout ;
wire \LessThan1~25_cout ;
wire \LessThan1~27_cout ;
wire \LessThan1~29_cout ;
wire \LessThan1~31_cout ;
wire \LessThan1~33_cout ;
wire \LessThan1~35_cout ;
wire \LessThan1~37_cout ;
wire \LessThan1~39_cout ;
wire \LessThan1~41_cout ;
wire \LessThan1~43_cout ;
wire \LessThan1~45_cout ;
wire \LessThan1~47_cout ;
wire \LessThan1~49_cout ;
wire \LessThan1~51_cout ;
wire \LessThan1~53_cout ;
wire \LessThan1~55_cout ;
wire \LessThan1~57_cout ;
wire \LessThan1~59_cout ;
wire \LessThan1~61_cout ;
wire \LessThan1~62_combout ;
wire \LessThan0~1_cout ;
wire \LessThan0~3_cout ;
wire \LessThan0~5_cout ;
wire \LessThan0~7_cout ;
wire \LessThan0~9_cout ;
wire \LessThan0~11_cout ;
wire \LessThan0~13_cout ;
wire \LessThan0~15_cout ;
wire \LessThan0~17_cout ;
wire \LessThan0~19_cout ;
wire \LessThan0~21_cout ;
wire \LessThan0~23_cout ;
wire \LessThan0~25_cout ;
wire \LessThan0~27_cout ;
wire \LessThan0~29_cout ;
wire \LessThan0~31_cout ;
wire \LessThan0~33_cout ;
wire \LessThan0~35_cout ;
wire \LessThan0~37_cout ;
wire \LessThan0~39_cout ;
wire \LessThan0~41_cout ;
wire \LessThan0~43_cout ;
wire \LessThan0~45_cout ;
wire \LessThan0~47_cout ;
wire \LessThan0~49_cout ;
wire \LessThan0~51_cout ;
wire \LessThan0~53_cout ;
wire \LessThan0~55_cout ;
wire \LessThan0~57_cout ;
wire \LessThan0~59_cout ;
wire \LessThan0~61_cout ;
wire \LessThan0~62_combout ;
wire \Selector31~3_combout ;
wire \Selector31~4_combout ;
wire \Selector31~5_combout ;
wire \ShiftRight0~106_combout ;
wire \Selector31~7_combout ;
wire \ShiftRight0~109_combout ;
wire \ShiftRight0~145_combout ;
wire \ShiftRight0~144_combout ;
wire \ShiftRight0~110_combout ;
wire \ShiftRight0~146_combout ;
wire \ShiftRight0~81_combout ;
wire \ShiftRight0~147_combout ;
wire \Selector20~1_combout ;
wire \ShiftRight0~111_combout ;
wire \ShiftLeft0~53_combout ;
wire \ShiftLeft0~106_combout ;
wire \Selector0~14_combout ;
wire \Selector16~0_combout ;
wire \Selector28~12_combout ;
wire \Selector0~21_combout ;
wire \Selector20~0_combout ;
wire \Selector2~2_combout ;
wire \Selector28~7_combout ;
wire \Selector0~17_combout ;
wire \Selector0~15_combout ;
wire \Selector28~2_combout ;
wire \Selector28~3_combout ;
wire \ShiftRight0~107_combout ;
wire \Selector2~14_combout ;
wire \ShiftRight0~141_combout ;
wire \Selector28~8_combout ;
wire \ShiftRight0~142_combout ;
wire \ShiftRight0~143_combout ;
wire \ShiftRight0~108_combout ;
wire \Selector28~9_combout ;
wire \Selector0~18_combout ;
wire \Selector28~4_combout ;
wire \Selector0~20_combout ;
wire \Add0~3 ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \Add1~3 ;
wire \Add1~5 ;
wire \Add1~6_combout ;
wire \Selector28~5_combout ;
wire \Selector28~6_combout ;
wire \Selector28~10_combout ;
wire \ShiftLeft0~58_combout ;
wire \ShiftLeft0~59_combout ;
wire \ShiftLeft0~109_combout ;
wire \Selector0~23_combout ;
wire \Selector0~16_combout ;
wire \Selector0~24_combout ;
wire \Selector0~25_combout ;
wire \Selector8~0_combout ;
wire \Selector0~26_combout ;
wire \Selector0~22_combout ;
wire \ShiftLeft0~57_combout ;
wire \ShiftLeft0~56_combout ;
wire \ShiftLeft0~108_combout ;
wire \ShiftLeft0~55_combout ;
wire \ShiftLeft0~54_combout ;
wire \ShiftLeft0~107_combout ;
wire \Selector0~28_combout ;
wire \ShiftLeft0~68_combout ;
wire \ShiftLeft0~67_combout ;
wire \ShiftLeft0~112_combout ;
wire \Selector0~41_combout ;
wire \Selector0~32_combout ;
wire \Selector0~33_combout ;
wire \Selector16~1_combout ;
wire \Selector0~34_combout ;
wire \ShiftLeft0~64_combout ;
wire \ShiftLeft0~63_combout ;
wire \ShiftLeft0~111_combout ;
wire \Selector8~1_combout ;
wire \ShiftLeft0~65_combout ;
wire \Selector0~40_combout ;
wire \Selector0~35_combout ;
wire \Selector0~36_combout ;
wire \Selector0~19_combout ;
wire \Add1~7 ;
wire \Add1~9 ;
wire \Add1~11 ;
wire \Add1~13 ;
wire \Add1~15 ;
wire \Add1~17 ;
wire \Add1~19 ;
wire \Add1~21 ;
wire \Add1~23 ;
wire \Add1~25 ;
wire \Add1~27 ;
wire \Add1~29 ;
wire \Add1~31 ;
wire \Add1~33 ;
wire \Add1~35 ;
wire \Add1~37 ;
wire \Add1~39 ;
wire \Add1~41 ;
wire \Add1~43 ;
wire \Add1~45 ;
wire \Add1~47 ;
wire \Add1~49 ;
wire \Add1~51 ;
wire \Add1~53 ;
wire \Add1~55 ;
wire \Add1~57 ;
wire \Add1~59 ;
wire \Add1~61 ;
wire \Add1~62_combout ;
wire \Selector0~37_combout ;
wire \Add0~7 ;
wire \Add0~9 ;
wire \Add0~11 ;
wire \Add0~13 ;
wire \Add0~15 ;
wire \Add0~17 ;
wire \Add0~19 ;
wire \Add0~21 ;
wire \Add0~23 ;
wire \Add0~25 ;
wire \Add0~27 ;
wire \Add0~29 ;
wire \Add0~31 ;
wire \Add0~33 ;
wire \Add0~35 ;
wire \Add0~37 ;
wire \Add0~39 ;
wire \Add0~41 ;
wire \Add0~43 ;
wire \Add0~45 ;
wire \Add0~47 ;
wire \Add0~49 ;
wire \Add0~51 ;
wire \Add0~53 ;
wire \Add0~55 ;
wire \Add0~57 ;
wire \Add0~59 ;
wire \Add0~61 ;
wire \Add0~62_combout ;
wire \ShiftLeft0~113_combout ;
wire \Selector2~12_combout ;
wire \Selector2~3_combout ;
wire \ShiftLeft0~70_combout ;
wire \Selector0~29_combout ;
wire \Selector2~4_combout ;
wire \Selector2~5_combout ;
wire \Selector2~7_combout ;
wire \Add0~58_combout ;
wire \Add1~58_combout ;
wire \Selector2~8_combout ;
wire \Selector2~9_combout ;
wire \ShiftLeft0~118_combout ;
wire \ShiftLeft0~117_combout ;
wire \ShiftLeft0~71_combout ;
wire \ShiftLeft0~116_combout ;
wire \ShiftLeft0~66_combout ;
wire \Selector2~10_combout ;
wire \Selector2~11_combout ;
wire \ShiftLeft0~73_combout ;
wire \Selector29~11_combout ;
wire \ShiftRight0~152_combout ;
wire \ShiftRight0~153_combout ;
wire \Selector21~0_combout ;
wire \ShiftRight0~151_combout ;
wire \ShiftRight0~113_combout ;
wire \ShiftRight0~114_combout ;
wire \Selector29~3_combout ;
wire \ShiftRight0~150_combout ;
wire \ShiftRight0~149_combout ;
wire \ShiftRight0~112_combout ;
wire \ShiftRight0~148_combout ;
wire \Selector29~7_combout ;
wire \Selector29~8_combout ;
wire \Selector29~4_combout ;
wire \Add1~4_combout ;
wire \Add0~4_combout ;
wire \Selector29~5_combout ;
wire \Selector29~6_combout ;
wire \Selector29~9_combout ;
wire \Selector5~6_combout ;
wire \Selector5~7_combout ;
wire \Selector5~8_combout ;
wire \Add0~52_combout ;
wire \Add1~52_combout ;
wire \Selector5~5_combout ;
wire \Selector5~9_combout ;
wire \Selector5~0_combout ;
wire \Selector5~1_combout ;
wire \ShiftLeft0~76_combout ;
wire \ShiftLeft0~77_combout ;
wire \ShiftLeft0~120_combout ;
wire \ShiftLeft0~78_combout ;
wire \ShiftLeft0~79_combout ;
wire \ShiftLeft0~121_combout ;
wire \ShiftLeft0~80_combout ;
wire \Selector5~2_combout ;
wire \ShiftLeft0~84_combout ;
wire \ShiftLeft0~123_combout ;
wire \ShiftLeft0~87_combout ;
wire \ShiftLeft0~88_combout ;
wire \Selector5~3_combout ;
wire \Selector5~4_combout ;
wire \ShiftLeft0~125_combout ;
wire \ShiftLeft0~89_combout ;
wire \ShiftLeft0~83_combout ;
wire \ShiftLeft0~126_combout ;
wire \ShiftLeft0~82_combout ;
wire \ShiftLeft0~81_combout ;
wire \ShiftLeft0~75_combout ;
wire \ShiftLeft0~129_combout ;
wire \ShiftLeft0~92_combout ;
wire \Selector3~6_combout ;
wire \ShiftLeft0~130_combout ;
wire \ShiftLeft0~74_combout ;
wire \ShiftLeft0~131_combout ;
wire \ShiftLeft0~93_combout ;
wire \Selector3~7_combout ;
wire \ShiftLeft0~86_combout ;
wire \ShiftLeft0~128_combout ;
wire \ShiftLeft0~85_combout ;
wire \ShiftLeft0~127_combout ;
wire \Selector11~0_combout ;
wire \ShiftLeft0~91_combout ;
wire \Selector3~0_combout ;
wire \Selector3~4_combout ;
wire \Selector3~2_combout ;
wire \Selector3~3_combout ;
wire \Add1~56_combout ;
wire \Add0~56_combout ;
wire \Selector3~1_combout ;
wire \Selector3~5_combout ;
wire \Selector0~30_combout ;
wire \Selector1~0_combout ;
wire \Add0~60_combout ;
wire \Selector1~9_combout ;
wire \Add1~60_combout ;
wire \Selector1~2_combout ;
wire \ShiftLeft0~122_combout ;
wire \Selector1~3_combout ;
wire \Selector1~4_combout ;
wire \Selector1~5_combout ;
wire \ShiftLeft0~119_combout ;
wire \Selector1~6_combout ;
wire \Selector0~27_combout ;
wire \Selector1~7_combout ;
wire \Selector1~8_combout ;
wire \Selector1~10_combout ;
wire \ShiftLeft0~96_combout ;
wire \ShiftLeft0~61_combout ;
wire \ShiftLeft0~62_combout ;
wire \ShiftLeft0~110_combout ;
wire \ShiftLeft0~97_combout ;
wire \ShiftLeft0~98_combout ;
wire \Selector4~2_combout ;
wire \Selector4~3_combout ;
wire \Selector4~7_combout ;
wire \Selector4~6_combout ;
wire \Selector4~5_combout ;
wire \Add1~54_combout ;
wire \Add0~54_combout ;
wire \Selector4~4_combout ;
wire \Selector4~8_combout ;
wire \ShiftLeft0~115_combout ;
wire \ShiftLeft0~114_combout ;
wire \Selector10~0_combout ;
wire \Selector10~1_combout ;
wire \Selector10~5_combout ;
wire \Selector10~3_combout ;
wire \Selector10~4_combout ;
wire \Selector10~6_combout ;
wire \Add0~42_combout ;
wire \Add1~42_combout ;
wire \Selector10~2_combout ;
wire \Selector10~7_combout ;
wire \Selector10~8_combout ;
wire \ShiftLeft0~100_combout ;
wire \ShiftLeft0~101_combout ;
wire \ShiftLeft0~102_combout ;
wire \Selector6~0_combout ;
wire \ShiftLeft0~99_combout ;
wire \Selector6~1_combout ;
wire \Selector6~2_combout ;
wire \Selector6~6_combout ;
wire \Selector6~4_combout ;
wire \Selector6~5_combout ;
wire \Add1~50_combout ;
wire \Add0~50_combout ;
wire \Selector6~3_combout ;
wire \Selector6~7_combout ;
wire \Selector7~5_combout ;
wire \Selector7~6_combout ;
wire \Selector7~4_combout ;
wire \Add1~48_combout ;
wire \Add0~48_combout ;
wire \Selector7~3_combout ;
wire \ShiftLeft0~104_combout ;
wire \ShiftLeft0~105_combout ;
wire \ShiftLeft0~103_combout ;
wire \Selector7~0_combout ;
wire \Selector7~1_combout ;
wire \Selector7~2_combout ;
wire \Selector11~1_combout ;
wire \Selector11~4_combout ;
wire \ShiftRight0~117_combout ;
wire \ShiftRight0~118_combout ;
wire \Selector11~2_combout ;
wire \Add1~40_combout ;
wire \Add0~40_combout ;
wire \Selector11~3_combout ;
wire \Selector11~7_combout ;
wire \Selector11~8_combout ;
wire \Add1~14_combout ;
wire \Selector24~2_combout ;
wire \Selector24~3_combout ;
wire \Selector24~4_combout ;
wire \Selector24~1_combout ;
wire \ShiftRight0~119_combout ;
wire \Selector24~5_combout ;
wire \ShiftRight0~120_combout ;
wire \ShiftRight0~121_combout ;
wire \Selector24~6_combout ;
wire \ShiftRight0~124_combout ;
wire \ShiftRight0~125_combout ;
wire \ShiftRight0~122_combout ;
wire \Selector25~4_combout ;
wire \Selector25~5_combout ;
wire \Selector25~0_combout ;
wire \Add0~12_combout ;
wire \Add1~12_combout ;
wire \Selector25~1_combout ;
wire \Selector25~2_combout ;
wire \Selector25~3_combout ;
wire \Selector13~3_combout ;
wire \Selector13~2_combout ;
wire \Add0~36_combout ;
wire \Selector13~1_combout ;
wire \Selector13~5_combout ;
wire \ShiftLeft0~124_combout ;
wire \Selector13~0_combout ;
wire \Selector13~6_combout ;
wire \Selector13~7_combout ;
wire \Selector12~2_combout ;
wire \Selector12~4_combout ;
wire \Add0~38_combout ;
wire \Add1~38_combout ;
wire \Selector12~1_combout ;
wire \Selector12~5_combout ;
wire \Selector12~0_combout ;
wire \Selector12~6_combout ;
wire \Selector12~7_combout ;
wire \Selector26~0_combout ;
wire \Selector26~2_combout ;
wire \Selector26~3_combout ;
wire \Selector26~4_combout ;
wire \ShiftRight0~126_combout ;
wire \ShiftRight0~115_combout ;
wire \ShiftRight0~116_combout ;
wire \Selector26~5_combout ;
wire \Selector27~0_combout ;
wire \Selector27~1_combout ;
wire \Selector27~2_combout ;
wire \Add0~8_combout ;
wire \Add1~8_combout ;
wire \Selector27~3_combout ;
wire \Selector27~4_combout ;
wire \ShiftRight0~127_combout ;
wire \Selector27~5_combout ;
wire \Selector27~6_combout ;
wire \Equal10~5_combout ;
wire \Equal10~3_combout ;
wire \Equal10~4_combout ;
wire \Equal10~0_combout ;
wire \Equal10~1_combout ;
wire \Equal10~2_combout ;
wire \Selector14~4_combout ;
wire \Selector14~5_combout ;
wire \Selector14~1_combout ;
wire \Add0~34_combout ;
wire \Selector14~2_combout ;
wire \Selector14~6_combout ;
wire \Selector14~0_combout ;
wire \Selector14~7_combout ;
wire \Selector15~0_combout ;
wire \Selector15~4_combout ;
wire \Selector15~2_combout ;
wire \Add1~32_combout ;
wire \Selector15~1_combout ;
wire \Selector15~5_combout ;
wire \Selector15~6_combout ;
wire \Selector15~7_combout ;
wire \Selector16~10_combout ;
wire \Selector0~39_combout ;
wire \Selector16~2_combout ;
wire \Selector16~3_combout ;
wire \Selector16~4_combout ;
wire \Add1~30_combout ;
wire \Add0~30_combout ;
wire \Selector16~5_combout ;
wire \Selector16~6_combout ;
wire \Selector16~7_combout ;
wire \Selector16~8_combout ;
wire \Selector16~9_combout ;
wire \ShiftRight0~123_combout ;
wire \Selector9~0_combout ;
wire \ShiftLeft0~95_combout ;
wire \Selector17~0_combout ;
wire \Selector17~1_combout ;
wire \Add0~28_combout ;
wire \Add1~28_combout ;
wire \Selector17~2_combout ;
wire \Selector17~3_combout ;
wire \Selector17~4_combout ;
wire \Selector17~5_combout ;
wire \Selector17~6_combout ;
wire \Selector20~2_combout ;
wire \Add1~22_combout ;
wire \Add0~22_combout ;
wire \Selector20~4_combout ;
wire \Selector20~5_combout ;
wire \Selector20~6_combout ;
wire \Selector20~7_combout ;
wire \Selector20~8_combout ;
wire \Add0~20_combout ;
wire \Selector21~3_combout ;
wire \Selector21~4_combout ;
wire \Selector21~5_combout ;
wire \Selector21~6_combout ;
wire \Selector21~7_combout ;
wire \Selector21~1_combout ;
wire \Selector18~0_combout ;
wire \Add0~26_combout ;
wire \Add1~26_combout ;
wire \Selector18~2_combout ;
wire \Selector18~3_combout ;
wire \Selector18~4_combout ;
wire \Selector18~5_combout ;
wire \Selector18~6_combout ;
wire \Selector19~1_combout ;
wire \Add1~24_combout ;
wire \Selector19~2_combout ;
wire \Selector19~3_combout ;
wire \Selector19~4_combout ;
wire \Selector19~5_combout ;
wire \Selector19~0_combout ;
wire \Selector19~6_combout ;
wire \Selector8~5_combout ;
wire \Selector8~6_combout ;
wire \Selector8~8_combout ;
wire \Add0~46_combout ;
wire \Add1~46_combout ;
wire \Selector8~4_combout ;
wire \Selector8~9_combout ;
wire \Selector9~1_combout ;
wire \Selector9~4_combout ;
wire \Add1~44_combout ;
wire \Selector9~3_combout ;
wire \Selector9~2_combout ;
wire \Selector9~7_combout ;
wire \Selector9~8_combout ;
wire \Selector22~2_combout ;
wire \Add1~18_combout ;
wire \Selector22~3_combout ;
wire \Selector22~4_combout ;
wire \Selector22~5_combout ;
wire \Selector22~6_combout ;
wire \Selector22~7_combout ;
wire \Selector22~1_combout ;
wire \Selector23~1_combout ;
wire \Add1~16_combout ;
wire \Add0~16_combout ;
wire \Selector23~3_combout ;
wire \Selector23~4_combout ;
wire \Selector23~5_combout ;
wire \Selector23~6_combout ;
wire \Selector23~7_combout ;
wire \Equal10~8_combout ;


// Location: LCCOMB_X53_Y41_N10
cycloneive_lcell_comb \Add0~10 (
// Equation(s):
// \Add0~10_combout  = (\Mux31~1_combout  & ((Mux26 & (\Add0~9  & VCC)) # (!Mux26 & (!\Add0~9 )))) # (!\Mux31~1_combout  & ((Mux26 & (!\Add0~9 )) # (!Mux26 & ((\Add0~9 ) # (GND)))))
// \Add0~11  = CARRY((\Mux31~1_combout  & (!Mux26 & !\Add0~9 )) # (!\Mux31~1_combout  & ((!\Add0~9 ) # (!Mux26))))

	.dataa(Mux31),
	.datab(Mux261),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
// synopsys translate_off
defparam \Add0~10 .lut_mask = 16'h9617;
defparam \Add0~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N14
cycloneive_lcell_comb \Add0~14 (
// Equation(s):
// \Add0~14_combout  = (\Mux29~1_combout  & ((Mux24 & (\Add0~13  & VCC)) # (!Mux24 & (!\Add0~13 )))) # (!\Mux29~1_combout  & ((Mux24 & (!\Add0~13 )) # (!Mux24 & ((\Add0~13 ) # (GND)))))
// \Add0~15  = CARRY((\Mux29~1_combout  & (!Mux24 & !\Add0~13 )) # (!\Mux29~1_combout  & ((!\Add0~13 ) # (!Mux24))))

	.dataa(Mux29),
	.datab(Mux241),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
// synopsys translate_off
defparam \Add0~14 .lut_mask = 16'h9617;
defparam \Add0~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N18
cycloneive_lcell_comb \Add0~18 (
// Equation(s):
// \Add0~18_combout  = (Mux22 & ((\Mux27~1_combout  & (\Add0~17  & VCC)) # (!\Mux27~1_combout  & (!\Add0~17 )))) # (!Mux22 & ((\Mux27~1_combout  & (!\Add0~17 )) # (!\Mux27~1_combout  & ((\Add0~17 ) # (GND)))))
// \Add0~19  = CARRY((Mux22 & (!\Mux27~1_combout  & !\Add0~17 )) # (!Mux22 & ((!\Add0~17 ) # (!\Mux27~1_combout ))))

	.dataa(Mux221),
	.datab(Mux27),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
// synopsys translate_off
defparam \Add0~18 .lut_mask = 16'h9617;
defparam \Add0~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N24
cycloneive_lcell_comb \Add0~24 (
// Equation(s):
// \Add0~24_combout  = ((\Mux24~1_combout  $ (Mux19 $ (!\Add0~23 )))) # (GND)
// \Add0~25  = CARRY((\Mux24~1_combout  & ((Mux19) # (!\Add0~23 ))) # (!\Mux24~1_combout  & (Mux19 & !\Add0~23 )))

	.dataa(Mux24),
	.datab(Mux191),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
// synopsys translate_off
defparam \Add0~24 .lut_mask = 16'h698E;
defparam \Add0~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N0
cycloneive_lcell_comb \Add0~32 (
// Equation(s):
// \Add0~32_combout  = ((\Mux20~1_combout  $ (Mux15 $ (!\Add0~31 )))) # (GND)
// \Add0~33  = CARRY((\Mux20~1_combout  & ((Mux15) # (!\Add0~31 ))) # (!\Mux20~1_combout  & (Mux15 & !\Add0~31 )))

	.dataa(Mux20),
	.datab(Mux152),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~31 ),
	.combout(\Add0~32_combout ),
	.cout(\Add0~33 ));
// synopsys translate_off
defparam \Add0~32 .lut_mask = 16'h698E;
defparam \Add0~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N12
cycloneive_lcell_comb \Add0~44 (
// Equation(s):
// \Add0~44_combout  = ((Mux9 $ (\Mux14~1_combout  $ (!\Add0~43 )))) # (GND)
// \Add0~45  = CARRY((Mux9 & ((\Mux14~1_combout ) # (!\Add0~43 ))) # (!Mux9 & (\Mux14~1_combout  & !\Add0~43 )))

	.dataa(Mux91),
	.datab(Mux14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~43 ),
	.combout(\Add0~44_combout ),
	.cout(\Add0~45 ));
// synopsys translate_off
defparam \Add0~44 .lut_mask = 16'h698E;
defparam \Add0~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N10
cycloneive_lcell_comb \Add1~10 (
// Equation(s):
// \Add1~10_combout  = (\Mux31~1_combout  & ((Mux26 & (!\Add1~9 )) # (!Mux26 & ((\Add1~9 ) # (GND))))) # (!\Mux31~1_combout  & ((Mux26 & (\Add1~9  & VCC)) # (!Mux26 & (!\Add1~9 ))))
// \Add1~11  = CARRY((\Mux31~1_combout  & ((!\Add1~9 ) # (!Mux26))) # (!\Mux31~1_combout  & (!Mux26 & !\Add1~9 )))

	.dataa(Mux31),
	.datab(Mux261),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h692B;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N20
cycloneive_lcell_comb \Add1~20 (
// Equation(s):
// \Add1~20_combout  = ((Mux21 $ (\Mux26~1_combout  $ (\Add1~19 )))) # (GND)
// \Add1~21  = CARRY((Mux21 & ((!\Add1~19 ) # (!\Mux26~1_combout ))) # (!Mux21 & (!\Mux26~1_combout  & !\Add1~19 )))

	.dataa(Mux211),
	.datab(Mux26),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~19 ),
	.combout(\Add1~20_combout ),
	.cout(\Add1~21 ));
// synopsys translate_off
defparam \Add1~20 .lut_mask = 16'h962B;
defparam \Add1~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N2
cycloneive_lcell_comb \Add1~34 (
// Equation(s):
// \Add1~34_combout  = (Mux14 & ((\Mux19~1_combout  & (!\Add1~33 )) # (!\Mux19~1_combout  & (\Add1~33  & VCC)))) # (!Mux14 & ((\Mux19~1_combout  & ((\Add1~33 ) # (GND))) # (!\Mux19~1_combout  & (!\Add1~33 ))))
// \Add1~35  = CARRY((Mux14 & (\Mux19~1_combout  & !\Add1~33 )) # (!Mux14 & ((\Mux19~1_combout ) # (!\Add1~33 ))))

	.dataa(Mux141),
	.datab(Mux192),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~33 ),
	.combout(\Add1~34_combout ),
	.cout(\Add1~35 ));
// synopsys translate_off
defparam \Add1~34 .lut_mask = 16'h694D;
defparam \Add1~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N4
cycloneive_lcell_comb \Add1~36 (
// Equation(s):
// \Add1~36_combout  = ((\Mux18~1_combout  $ (Mux13 $ (\Add1~35 )))) # (GND)
// \Add1~37  = CARRY((\Mux18~1_combout  & (Mux13 & !\Add1~35 )) # (!\Mux18~1_combout  & ((Mux13) # (!\Add1~35 ))))

	.dataa(Mux182),
	.datab(Mux131),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~35 ),
	.combout(\Add1~36_combout ),
	.cout(\Add1~37 ));
// synopsys translate_off
defparam \Add1~36 .lut_mask = 16'h964D;
defparam \Add1~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N22
cycloneive_lcell_comb \ShiftRight0~52 (
// Equation(s):
// \ShiftRight0~52_combout  = (\Mux5~4_combout ) # ((\Mux5~1_combout ) # ((\Mux7~1_combout ) # (\Mux6~0_combout )))

	.dataa(Mux51),
	.datab(Mux5),
	.datac(Mux7),
	.datad(Mux6),
	.cin(gnd),
	.combout(\ShiftRight0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~52 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N6
cycloneive_lcell_comb \ShiftRight0~63 (
// Equation(s):
// \ShiftRight0~63_combout  = (\Mux36~4_combout  & (Mux27)) # (!\Mux36~4_combout  & ((Mux28)))

	.dataa(Mux36),
	.datab(gnd),
	.datac(Mux271),
	.datad(Mux281),
	.cin(gnd),
	.combout(\ShiftRight0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~63 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N6
cycloneive_lcell_comb \ShiftRight0~103 (
// Equation(s):
// \ShiftRight0~103_combout  = (\Mux36~4_combout  & (Mux12)) # (!\Mux36~4_combout  & ((Mux13)))

	.dataa(Mux36),
	.datab(gnd),
	.datac(Mux121),
	.datad(Mux131),
	.cin(gnd),
	.combout(\ShiftRight0~103_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~103 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N26
cycloneive_lcell_comb \Selector31~2 (
// Equation(s):
// \Selector31~2_combout  = (!Mux31 & (\Selector0~11_combout  & !\Mux36~4_combout ))

	.dataa(Mux311),
	.datab(gnd),
	.datac(\Selector0~11_combout ),
	.datad(Mux36),
	.cin(gnd),
	.combout(\Selector31~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~2 .lut_mask = 16'h0050;
defparam \Selector31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N6
cycloneive_lcell_comb \Selector0~31 (
// Equation(s):
// \Selector0~31_combout  = (\Selector0~30_combout  & ((\ShiftLeft0~66_combout ) # ((\Selector0~41_combout )))) # (!\Selector0~30_combout  & (((Mux0 & !\Selector0~41_combout ))))

	.dataa(\Selector0~30_combout ),
	.datab(\ShiftLeft0~66_combout ),
	.datac(Mux0),
	.datad(\Selector0~41_combout ),
	.cin(gnd),
	.combout(\Selector0~31_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~31 .lut_mask = 16'hAAD8;
defparam \Selector0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N10
cycloneive_lcell_comb \Selector2~6 (
// Equation(s):
// \Selector2~6_combout  = (Mux2) # ((\Selector0~18_combout ) # (\Mux7~1_combout ))

	.dataa(Mux2),
	.datab(gnd),
	.datac(\Selector0~18_combout ),
	.datad(Mux7),
	.cin(gnd),
	.combout(\Selector2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~6 .lut_mask = 16'hFFFA;
defparam \Selector2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N22
cycloneive_lcell_comb \ShiftLeft0~72 (
// Equation(s):
// \ShiftLeft0~72_combout  = (!\Mux36~4_combout  & ((\Mux35~4_combout  & (Mux31)) # (!\Mux35~4_combout  & ((Mux29)))))

	.dataa(Mux311),
	.datab(Mux352),
	.datac(Mux36),
	.datad(Mux291),
	.cin(gnd),
	.combout(\ShiftLeft0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~72 .lut_mask = 16'h0B08;
defparam \ShiftLeft0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N30
cycloneive_lcell_comb \Selector29~2 (
// Equation(s):
// \Selector29~2_combout  = (\Selector0~15_combout ) # ((Mux29 & \Selector0~16_combout ))

	.dataa(Mux291),
	.datab(gnd),
	.datac(\Selector0~15_combout ),
	.datad(\Selector0~16_combout ),
	.cin(gnd),
	.combout(\Selector29~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~2 .lut_mask = 16'hFAF0;
defparam \Selector29~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N30
cycloneive_lcell_comb \Selector1~1 (
// Equation(s):
// \Selector1~1_combout  = (\Selector0~17_combout  & (Mux1 $ (((\Mux5~1_combout ) # (\Mux6~0_combout )))))

	.dataa(Mux5),
	.datab(Mux6),
	.datac(Mux1),
	.datad(\Selector0~17_combout ),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~1 .lut_mask = 16'h1E00;
defparam \Selector1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N12
cycloneive_lcell_comb \Selector4~1 (
// Equation(s):
// \Selector4~1_combout  = (\Selector5~0_combout  & (((\Selector5~1_combout ) # (\ShiftLeft0~108_combout )))) # (!\Selector5~0_combout  & (\ShiftLeft0~112_combout  & (!\Selector5~1_combout )))

	.dataa(\Selector5~0_combout ),
	.datab(\ShiftLeft0~112_combout ),
	.datac(\Selector5~1_combout ),
	.datad(\ShiftLeft0~108_combout ),
	.cin(gnd),
	.combout(\Selector4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~1 .lut_mask = 16'hAEA4;
defparam \Selector4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N28
cycloneive_lcell_comb \Selector11~5 (
// Equation(s):
// \Selector11~5_combout  = (\Mux16~1_combout  & (\Selector0~15_combout )) # (!\Mux16~1_combout  & (((\Selector0~18_combout  & !Mux11))))

	.dataa(\Selector0~15_combout ),
	.datab(\Selector0~18_combout ),
	.datac(Mux16),
	.datad(Mux111),
	.cin(gnd),
	.combout(\Selector11~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~5 .lut_mask = 16'hA0AC;
defparam \Selector11~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N10
cycloneive_lcell_comb \Selector11~6 (
// Equation(s):
// \Selector11~6_combout  = (\Selector11~5_combout ) # ((\Selector0~17_combout  & (\Mux16~1_combout  $ (Mux11))))

	.dataa(Mux16),
	.datab(\Selector11~5_combout ),
	.datac(\Selector0~17_combout ),
	.datad(Mux111),
	.cin(gnd),
	.combout(\Selector11~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~6 .lut_mask = 16'hDCEC;
defparam \Selector11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N26
cycloneive_lcell_comb \Selector13~4 (
// Equation(s):
// \Selector13~4_combout  = (\Mux18~1_combout  & (((\Selector0~15_combout )))) # (!\Mux18~1_combout  & (\Selector0~18_combout  & ((!Mux13))))

	.dataa(\Selector0~18_combout ),
	.datab(\Selector0~15_combout ),
	.datac(Mux131),
	.datad(Mux182),
	.cin(gnd),
	.combout(\Selector13~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~4 .lut_mask = 16'hCC0A;
defparam \Selector13~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N10
cycloneive_lcell_comb \Selector12~3 (
// Equation(s):
// \Selector12~3_combout  = (\Selector0~17_combout  & (Mux12 $ (((\Mux5~1_combout ) # (\Mux17~0_combout )))))

	.dataa(Mux121),
	.datab(Mux5),
	.datac(Mux17),
	.datad(\Selector0~17_combout ),
	.cin(gnd),
	.combout(\Selector12~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~3 .lut_mask = 16'h5600;
defparam \Selector12~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N10
cycloneive_lcell_comb \Selector26~1 (
// Equation(s):
// \Selector26~1_combout  = (\Selector0~13_combout  & ((\Add0~10_combout ) # ((\Selector0~12_combout  & \Add1~10_combout )))) # (!\Selector0~13_combout  & (\Selector0~12_combout  & (\Add1~10_combout )))

	.dataa(\Selector0~13_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Add1~10_combout ),
	.datad(\Add0~10_combout ),
	.cin(gnd),
	.combout(\Selector26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~1 .lut_mask = 16'hEAC0;
defparam \Selector26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N14
cycloneive_lcell_comb \Selector14~3 (
// Equation(s):
// \Selector14~3_combout  = (Mux14 & ((\Selector0~15_combout ) # ((\Selector0~16_combout  & \Mux19~1_combout ))))

	.dataa(\Selector0~15_combout ),
	.datab(\Selector0~16_combout ),
	.datac(Mux141),
	.datad(Mux192),
	.cin(gnd),
	.combout(\Selector14~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~3 .lut_mask = 16'hE0A0;
defparam \Selector14~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N30
cycloneive_lcell_comb \Selector15~3 (
// Equation(s):
// \Selector15~3_combout  = (\Selector0~17_combout  & (\Mux20~1_combout  $ (Mux15)))

	.dataa(\Selector0~17_combout ),
	.datab(Mux20),
	.datac(Mux152),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector15~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~3 .lut_mask = 16'h2828;
defparam \Selector15~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N10
cycloneive_lcell_comb \Selector20~3 (
// Equation(s):
// \Selector20~3_combout  = (\Selector0~15_combout  & (((Mux20) # (\Mux25~1_combout )))) # (!\Selector0~15_combout  & (\Selector0~16_combout  & (Mux20 & \Mux25~1_combout )))

	.dataa(\Selector0~15_combout ),
	.datab(\Selector0~16_combout ),
	.datac(Mux201),
	.datad(Mux25),
	.cin(gnd),
	.combout(\Selector20~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~3 .lut_mask = 16'hEAA0;
defparam \Selector20~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N14
cycloneive_lcell_comb \Selector21~2 (
// Equation(s):
// \Selector21~2_combout  = (\Selector0~15_combout  & (((\Mux26~1_combout ) # (Mux21)))) # (!\Selector0~15_combout  & (\Selector0~16_combout  & (\Mux26~1_combout  & Mux21)))

	.dataa(\Selector0~15_combout ),
	.datab(\Selector0~16_combout ),
	.datac(Mux26),
	.datad(Mux211),
	.cin(gnd),
	.combout(\Selector21~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~2 .lut_mask = 16'hEAA0;
defparam \Selector21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N2
cycloneive_lcell_comb \Selector18~1 (
// Equation(s):
// \Selector18~1_combout  = (\Selector0~15_combout  & (((\Mux23~1_combout ) # (Mux18)))) # (!\Selector0~15_combout  & (\Selector0~16_combout  & (\Mux23~1_combout  & Mux18)))

	.dataa(\Selector0~16_combout ),
	.datab(\Selector0~15_combout ),
	.datac(Mux23),
	.datad(Mux181),
	.cin(gnd),
	.combout(\Selector18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~1 .lut_mask = 16'hECC0;
defparam \Selector18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N26
cycloneive_lcell_comb \Selector8~7 (
// Equation(s):
// \Selector8~7_combout  = (\Mux13~1_combout  & (((\Selector0~15_combout )))) # (!\Mux13~1_combout  & (!Mux8 & ((\Selector0~18_combout ))))

	.dataa(Mux81),
	.datab(\Selector0~15_combout ),
	.datac(\Selector0~18_combout ),
	.datad(Mux132),
	.cin(gnd),
	.combout(\Selector8~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~7 .lut_mask = 16'hCC50;
defparam \Selector8~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N0
cycloneive_lcell_comb \Selector9~5 (
// Equation(s):
// \Selector9~5_combout  = (\Mux14~1_combout  & (\Selector0~15_combout )) # (!\Mux14~1_combout  & (((!Mux9 & \Selector0~18_combout ))))

	.dataa(Mux14),
	.datab(\Selector0~15_combout ),
	.datac(Mux91),
	.datad(\Selector0~18_combout ),
	.cin(gnd),
	.combout(\Selector9~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~5 .lut_mask = 16'h8D88;
defparam \Selector9~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N30
cycloneive_lcell_comb \Selector9~6 (
// Equation(s):
// \Selector9~6_combout  = (\Selector9~5_combout ) # ((\Selector0~17_combout  & (Mux9 $ (\Mux14~1_combout ))))

	.dataa(\Selector0~17_combout ),
	.datab(\Selector9~5_combout ),
	.datac(Mux91),
	.datad(Mux14),
	.cin(gnd),
	.combout(\Selector9~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~6 .lut_mask = 16'hCEEC;
defparam \Selector9~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N6
cycloneive_lcell_comb \Selector23~2 (
// Equation(s):
// \Selector23~2_combout  = (\Mux28~1_combout  & ((\Selector0~15_combout ) # ((\Selector0~16_combout  & Mux23)))) # (!\Mux28~1_combout  & (((\Selector0~15_combout  & Mux23))))

	.dataa(Mux28),
	.datab(\Selector0~16_combout ),
	.datac(\Selector0~15_combout ),
	.datad(Mux231),
	.cin(gnd),
	.combout(\Selector23~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~2 .lut_mask = 16'hF8A0;
defparam \Selector23~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N14
cycloneive_lcell_comb \Selector30~8 (
// Equation(s):
// Selector30 = (\Selector30~4_combout ) # ((\Selector30~7_combout ) # ((\Selector30~0_combout ) # (\Selector30~2_combout )))

	.dataa(\Selector30~4_combout ),
	.datab(\Selector30~7_combout ),
	.datac(\Selector30~0_combout ),
	.datad(\Selector30~2_combout ),
	.cin(gnd),
	.combout(Selector30),
	.cout());
// synopsys translate_off
defparam \Selector30~8 .lut_mask = 16'hFFFE;
defparam \Selector30~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N6
cycloneive_lcell_comb \ShiftRight0~100 (
// Equation(s):
// ShiftRight0 = (\Mux34~3_combout  & (\ShiftRight0~137_combout )) # (!\Mux34~3_combout  & ((\ShiftRight0~138_combout )))

	.dataa(Mux34),
	.datab(gnd),
	.datac(\ShiftRight0~137_combout ),
	.datad(\ShiftRight0~138_combout ),
	.cin(gnd),
	.combout(ShiftRight0),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~100 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N6
cycloneive_lcell_comb \Selector31~6 (
// Equation(s):
// Selector31 = (\Selector31~0_combout ) # ((\Selector31~5_combout ) # ((\Mux36~4_combout  & \Selector0~8_combout )))

	.dataa(Mux36),
	.datab(\Selector0~8_combout ),
	.datac(\Selector31~0_combout ),
	.datad(\Selector31~5_combout ),
	.cin(gnd),
	.combout(Selector31),
	.cout());
// synopsys translate_off
defparam \Selector31~6 .lut_mask = 16'hFFF8;
defparam \Selector31~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N8
cycloneive_lcell_comb \Selector31~8 (
// Equation(s):
// Selector311 = (\Selector0~8_combout ) # ((\Selector31~7_combout ) # ((\Mux36~4_combout  & \Selector0~9_combout )))

	.dataa(Mux36),
	.datab(\Selector0~8_combout ),
	.datac(\Selector31~7_combout ),
	.datad(\Selector0~9_combout ),
	.cin(gnd),
	.combout(Selector311),
	.cout());
// synopsys translate_off
defparam \Selector31~8 .lut_mask = 16'hFEFC;
defparam \Selector31~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N2
cycloneive_lcell_comb \Selector28~11 (
// Equation(s):
// Selector28 = (\Selector28~12_combout ) # ((\Selector28~10_combout ) # ((\ShiftRight0~111_combout  & \Selector20~0_combout )))

	.dataa(\ShiftRight0~111_combout ),
	.datab(\Selector28~12_combout ),
	.datac(\Selector20~0_combout ),
	.datad(\Selector28~10_combout ),
	.cin(gnd),
	.combout(Selector28),
	.cout());
// synopsys translate_off
defparam \Selector28~11 .lut_mask = 16'hFFEC;
defparam \Selector28~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N0
cycloneive_lcell_comb \ShiftLeft0~60 (
// Equation(s):
// ShiftLeft0 = (\Mux34~3_combout  & (\ShiftLeft0~106_combout )) # (!\Mux34~3_combout  & ((\ShiftLeft0~109_combout )))

	.dataa(Mux34),
	.datab(\ShiftLeft0~106_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~109_combout ),
	.cin(gnd),
	.combout(ShiftLeft0),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~60 .lut_mask = 16'hDD88;
defparam \ShiftLeft0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N20
cycloneive_lcell_comb \Selector0~38 (
// Equation(s):
// Selector0 = (\Selector0~36_combout ) # ((\Selector0~37_combout ) # ((\Selector0~20_combout  & \Add0~62_combout )))

	.dataa(\Selector0~36_combout ),
	.datab(\Selector0~20_combout ),
	.datac(\Selector0~37_combout ),
	.datad(\Add0~62_combout ),
	.cin(gnd),
	.combout(Selector0),
	.cout());
// synopsys translate_off
defparam \Selector0~38 .lut_mask = 16'hFEFA;
defparam \Selector0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N6
cycloneive_lcell_comb \ShiftLeft0~69 (
// Equation(s):
// ShiftLeft01 = (\Mux34~3_combout  & (((\ShiftLeft0~52_combout  & !\Mux35~4_combout )))) # (!\Mux34~3_combout  & (\ShiftLeft0~113_combout ))

	.dataa(Mux34),
	.datab(\ShiftLeft0~113_combout ),
	.datac(\ShiftLeft0~52_combout ),
	.datad(Mux352),
	.cin(gnd),
	.combout(ShiftLeft01),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~69 .lut_mask = 16'h44E4;
defparam \ShiftLeft0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N26
cycloneive_lcell_comb \Selector2~13 (
// Equation(s):
// Selector2 = (\Selector2~4_combout ) # ((\Selector2~9_combout ) # ((\Selector2~12_combout  & \Selector2~11_combout )))

	.dataa(\Selector2~12_combout ),
	.datab(\Selector2~4_combout ),
	.datac(\Selector2~9_combout ),
	.datad(\Selector2~11_combout ),
	.cin(gnd),
	.combout(Selector2),
	.cout());
// synopsys translate_off
defparam \Selector2~13 .lut_mask = 16'hFEFC;
defparam \Selector2~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N10
cycloneive_lcell_comb \Selector29~10 (
// Equation(s):
// Selector29 = (\Selector29~11_combout ) # ((\Selector29~9_combout ) # ((\Selector20~0_combout  & \ShiftRight0~114_combout )))

	.dataa(\Selector29~11_combout ),
	.datab(\Selector20~0_combout ),
	.datac(\ShiftRight0~114_combout ),
	.datad(\Selector29~9_combout ),
	.cin(gnd),
	.combout(Selector29),
	.cout());
// synopsys translate_off
defparam \Selector29~10 .lut_mask = 16'hFFEA;
defparam \Selector29~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N6
cycloneive_lcell_comb \Selector4~0 (
// Equation(s):
// Selector4 = (\Selector0~6_combout  & (!\Mux32~4_combout  & (!\ShiftRight0~61_combout  & !\Mux33~3_combout )))

	.dataa(\Selector0~6_combout ),
	.datab(Mux32),
	.datac(\ShiftRight0~61_combout ),
	.datad(Mux33),
	.cin(gnd),
	.combout(Selector4),
	.cout());
// synopsys translate_off
defparam \Selector4~0 .lut_mask = 16'h0002;
defparam \Selector4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N30
cycloneive_lcell_comb \Selector5~10 (
// Equation(s):
// Selector5 = (\Selector5~9_combout ) # ((\Selector5~4_combout ) # ((\ShiftRight0~113_combout  & Selector4)))

	.dataa(\ShiftRight0~113_combout ),
	.datab(Selector4),
	.datac(\Selector5~9_combout ),
	.datad(\Selector5~4_combout ),
	.cin(gnd),
	.combout(Selector5),
	.cout());
// synopsys translate_off
defparam \Selector5~10 .lut_mask = 16'hFFF8;
defparam \Selector5~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N4
cycloneive_lcell_comb \ShiftLeft0~90 (
// Equation(s):
// ShiftLeft02 = (\Mux34~3_combout  & (\ShiftLeft0~125_combout )) # (!\Mux34~3_combout  & ((\ShiftLeft0~126_combout )))

	.dataa(gnd),
	.datab(Mux34),
	.datac(\ShiftLeft0~125_combout ),
	.datad(\ShiftLeft0~126_combout ),
	.cin(gnd),
	.combout(ShiftLeft02),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~90 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N2
cycloneive_lcell_comb \Selector3~8 (
// Equation(s):
// Selector3 = (\Selector3~0_combout ) # ((\Selector3~5_combout ) # ((\Selector2~12_combout  & \Selector3~7_combout )))

	.dataa(\Selector2~12_combout ),
	.datab(\Selector3~7_combout ),
	.datac(\Selector3~0_combout ),
	.datad(\Selector3~5_combout ),
	.cin(gnd),
	.combout(Selector3),
	.cout());
// synopsys translate_off
defparam \Selector3~8 .lut_mask = 16'hFFF8;
defparam \Selector3~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N26
cycloneive_lcell_comb \ShiftLeft0~94 (
// Equation(s):
// ShiftLeft03 = (\Mux34~3_combout  & (\ShiftLeft0~73_combout )) # (!\Mux34~3_combout  & ((\ShiftLeft0~123_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~73_combout ),
	.datac(Mux34),
	.datad(\ShiftLeft0~123_combout ),
	.cin(gnd),
	.combout(ShiftLeft03),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~94 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N20
cycloneive_lcell_comb \Selector1~11 (
// Equation(s):
// Selector1 = (\Selector1~0_combout ) # ((\Selector1~10_combout ) # ((\Selector0~20_combout  & \Add0~60_combout )))

	.dataa(\Selector1~0_combout ),
	.datab(\Selector0~20_combout ),
	.datac(\Add0~60_combout ),
	.datad(\Selector1~10_combout ),
	.cin(gnd),
	.combout(Selector1),
	.cout());
// synopsys translate_off
defparam \Selector1~11 .lut_mask = 16'hFFEA;
defparam \Selector1~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N26
cycloneive_lcell_comb \Selector4~9 (
// Equation(s):
// Selector41 = (\Selector4~3_combout ) # ((\Selector4~8_combout ) # ((\ShiftRight0~110_combout  & Selector4)))

	.dataa(\Selector4~3_combout ),
	.datab(\ShiftRight0~110_combout ),
	.datac(Selector4),
	.datad(\Selector4~8_combout ),
	.cin(gnd),
	.combout(Selector41),
	.cout());
// synopsys translate_off
defparam \Selector4~9 .lut_mask = 16'hFFEA;
defparam \Selector4~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N12
cycloneive_lcell_comb \Selector10~9 (
// Equation(s):
// Selector10 = (\Selector10~8_combout ) # ((ShiftLeft01 & (!\Mux33~3_combout  & \Selector0~29_combout )))

	.dataa(ShiftLeft01),
	.datab(Mux33),
	.datac(\Selector0~29_combout ),
	.datad(\Selector10~8_combout ),
	.cin(gnd),
	.combout(Selector10),
	.cout());
// synopsys translate_off
defparam \Selector10~9 .lut_mask = 16'hFF20;
defparam \Selector10~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N28
cycloneive_lcell_comb \Selector6~8 (
// Equation(s):
// Selector6 = (\Selector6~2_combout ) # ((\Selector6~7_combout ) # ((Selector4 & \ShiftRight0~78_combout )))

	.dataa(Selector4),
	.datab(\Selector6~2_combout ),
	.datac(\Selector6~7_combout ),
	.datad(\ShiftRight0~78_combout ),
	.cin(gnd),
	.combout(Selector6),
	.cout());
// synopsys translate_off
defparam \Selector6~8 .lut_mask = 16'hFEFC;
defparam \Selector6~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N24
cycloneive_lcell_comb \Selector7~7 (
// Equation(s):
// Selector7 = (\Selector7~6_combout ) # ((\Selector7~4_combout ) # ((\Selector7~3_combout ) # (\Selector7~2_combout )))

	.dataa(\Selector7~6_combout ),
	.datab(\Selector7~4_combout ),
	.datac(\Selector7~3_combout ),
	.datad(\Selector7~2_combout ),
	.cin(gnd),
	.combout(Selector7),
	.cout());
// synopsys translate_off
defparam \Selector7~7 .lut_mask = 16'hFFFE;
defparam \Selector7~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N26
cycloneive_lcell_comb \Selector7~8 (
// Equation(s):
// Selector71 = (Selector7) # ((Selector4 & ShiftRight0))

	.dataa(Selector4),
	.datab(gnd),
	.datac(ShiftRight0),
	.datad(Selector7),
	.cin(gnd),
	.combout(Selector71),
	.cout());
// synopsys translate_off
defparam \Selector7~8 .lut_mask = 16'hFFA0;
defparam \Selector7~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N14
cycloneive_lcell_comb \Selector11~9 (
// Equation(s):
// Selector11 = (\Selector11~8_combout ) # ((\Selector0~29_combout  & (!\Mux33~3_combout  & ShiftLeft02)))

	.dataa(\Selector0~29_combout ),
	.datab(Mux33),
	.datac(ShiftLeft02),
	.datad(\Selector11~8_combout ),
	.cin(gnd),
	.combout(Selector11),
	.cout());
// synopsys translate_off
defparam \Selector11~9 .lut_mask = 16'hFF20;
defparam \Selector11~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N14
cycloneive_lcell_comb \Selector24~7 (
// Equation(s):
// Selector24 = (\Selector24~4_combout ) # ((\Selector24~1_combout ) # ((\Selector24~6_combout  & \Selector24~0_combout )))

	.dataa(\Selector24~4_combout ),
	.datab(\Selector24~1_combout ),
	.datac(\Selector24~6_combout ),
	.datad(\Selector24~0_combout ),
	.cin(gnd),
	.combout(Selector24),
	.cout());
// synopsys translate_off
defparam \Selector24~7 .lut_mask = 16'hFEEE;
defparam \Selector24~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N26
cycloneive_lcell_comb \Selector24~8 (
// Equation(s):
// Selector241 = (!\ShiftRight0~61_combout  & (\Selector0~7_combout  & (!\Mux32~4_combout  & !\Mux33~3_combout )))

	.dataa(\ShiftRight0~61_combout ),
	.datab(\Selector0~7_combout ),
	.datac(Mux32),
	.datad(Mux33),
	.cin(gnd),
	.combout(Selector241),
	.cout());
// synopsys translate_off
defparam \Selector24~8 .lut_mask = 16'h0004;
defparam \Selector24~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N8
cycloneive_lcell_comb \Selector24~9 (
// Equation(s):
// Selector242 = (Selector24) # ((Selector241 & ShiftLeft0))

	.dataa(Selector241),
	.datab(ShiftLeft0),
	.datac(gnd),
	.datad(Selector24),
	.cin(gnd),
	.combout(Selector242),
	.cout());
// synopsys translate_off
defparam \Selector24~9 .lut_mask = 16'hFF88;
defparam \Selector24~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N18
cycloneive_lcell_comb \Selector25~6 (
// Equation(s):
// Selector25 = (\Selector25~0_combout ) # ((\Selector25~3_combout ) # ((\Selector25~5_combout  & \Selector24~0_combout )))

	.dataa(\Selector25~5_combout ),
	.datab(\Selector25~0_combout ),
	.datac(\Selector25~3_combout ),
	.datad(\Selector24~0_combout ),
	.cin(gnd),
	.combout(Selector25),
	.cout());
// synopsys translate_off
defparam \Selector25~6 .lut_mask = 16'hFEFC;
defparam \Selector25~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N18
cycloneive_lcell_comb \Selector25~7 (
// Equation(s):
// Selector251 = (Selector25) # ((ShiftLeft03 & Selector241))

	.dataa(gnd),
	.datab(ShiftLeft03),
	.datac(Selector25),
	.datad(Selector241),
	.cin(gnd),
	.combout(Selector251),
	.cout());
// synopsys translate_off
defparam \Selector25~7 .lut_mask = 16'hFCF0;
defparam \Selector25~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N8
cycloneive_lcell_comb \Selector13~8 (
// Equation(s):
// Selector13 = (\Selector13~7_combout ) # ((\Selector0~29_combout  & (\ShiftRight0~107_combout  & \ShiftLeft0~73_combout )))

	.dataa(\Selector0~29_combout ),
	.datab(\ShiftRight0~107_combout ),
	.datac(\Selector13~7_combout ),
	.datad(\ShiftLeft0~73_combout ),
	.cin(gnd),
	.combout(Selector13),
	.cout());
// synopsys translate_off
defparam \Selector13~8 .lut_mask = 16'hF8F0;
defparam \Selector13~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N12
cycloneive_lcell_comb \Selector12~8 (
// Equation(s):
// Selector12 = (\Selector12~7_combout ) # ((\ShiftLeft0~106_combout  & (\ShiftRight0~107_combout  & \Selector0~29_combout )))

	.dataa(\ShiftLeft0~106_combout ),
	.datab(\ShiftRight0~107_combout ),
	.datac(\Selector12~7_combout ),
	.datad(\Selector0~29_combout ),
	.cin(gnd),
	.combout(Selector12),
	.cout());
// synopsys translate_off
defparam \Selector12~8 .lut_mask = 16'hF8F0;
defparam \Selector12~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N24
cycloneive_lcell_comb \Selector26~6 (
// Equation(s):
// Selector26 = (\Selector26~0_combout ) # ((\Selector26~3_combout ) # ((\Selector24~0_combout  & \Selector26~5_combout )))

	.dataa(\Selector24~0_combout ),
	.datab(\Selector26~0_combout ),
	.datac(\Selector26~3_combout ),
	.datad(\Selector26~5_combout ),
	.cin(gnd),
	.combout(Selector26),
	.cout());
// synopsys translate_off
defparam \Selector26~6 .lut_mask = 16'hFEFC;
defparam \Selector26~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N30
cycloneive_lcell_comb \Selector26~7 (
// Equation(s):
// Selector261 = (Selector26) # ((ShiftLeft01 & Selector241))

	.dataa(gnd),
	.datab(ShiftLeft01),
	.datac(Selector241),
	.datad(Selector26),
	.cin(gnd),
	.combout(Selector261),
	.cout());
// synopsys translate_off
defparam \Selector26~7 .lut_mask = 16'hFFC0;
defparam \Selector26~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N20
cycloneive_lcell_comb \Selector27~7 (
// Equation(s):
// Selector27 = (\Selector27~1_combout ) # ((\Selector27~4_combout ) # ((\Selector27~6_combout  & \Selector24~0_combout )))

	.dataa(\Selector27~1_combout ),
	.datab(\Selector27~4_combout ),
	.datac(\Selector27~6_combout ),
	.datad(\Selector24~0_combout ),
	.cin(gnd),
	.combout(Selector27),
	.cout());
// synopsys translate_off
defparam \Selector27~7 .lut_mask = 16'hFEEE;
defparam \Selector27~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N30
cycloneive_lcell_comb \Selector27~8 (
// Equation(s):
// Selector271 = (Selector27) # ((ShiftLeft02 & Selector241))

	.dataa(Selector27),
	.datab(ShiftLeft02),
	.datac(Selector241),
	.datad(gnd),
	.cin(gnd),
	.combout(Selector271),
	.cout());
// synopsys translate_off
defparam \Selector27~8 .lut_mask = 16'hEAEA;
defparam \Selector27~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N20
cycloneive_lcell_comb \Equal10~6 (
// Equation(s):
// Equal10 = (\Equal10~5_combout  & (\Equal10~4_combout  & \Equal10~2_combout ))

	.dataa(\Equal10~5_combout ),
	.datab(gnd),
	.datac(\Equal10~4_combout ),
	.datad(\Equal10~2_combout ),
	.cin(gnd),
	.combout(Equal10),
	.cout());
// synopsys translate_off
defparam \Equal10~6 .lut_mask = 16'hA000;
defparam \Equal10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N22
cycloneive_lcell_comb \Selector14~8 (
// Equation(s):
// Selector14 = (\Selector14~7_combout ) # ((\ShiftLeft0~100_combout  & (!\Mux33~3_combout  & \Selector0~29_combout )))

	.dataa(\ShiftLeft0~100_combout ),
	.datab(Mux33),
	.datac(\Selector0~29_combout ),
	.datad(\Selector14~7_combout ),
	.cin(gnd),
	.combout(Selector14),
	.cout());
// synopsys translate_off
defparam \Selector14~8 .lut_mask = 16'hFF20;
defparam \Selector14~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N28
cycloneive_lcell_comb \Selector15~8 (
// Equation(s):
// Selector15 = (\Selector15~0_combout ) # ((\Selector15~7_combout ) # ((\ShiftRight0~105_combout  & \Selector8~0_combout )))

	.dataa(\ShiftRight0~105_combout ),
	.datab(\Selector8~0_combout ),
	.datac(\Selector15~0_combout ),
	.datad(\Selector15~7_combout ),
	.cin(gnd),
	.combout(Selector15),
	.cout());
// synopsys translate_off
defparam \Selector15~8 .lut_mask = 16'hFFF8;
defparam \Selector15~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N26
cycloneive_lcell_comb \Selector16~11 (
// Equation(s):
// Selector16 = (\Selector16~3_combout ) # ((\Selector16~9_combout ) # ((\Selector16~10_combout  & \ShiftRight0~119_combout )))

	.dataa(\Selector16~10_combout ),
	.datab(\ShiftRight0~119_combout ),
	.datac(\Selector16~3_combout ),
	.datad(\Selector16~9_combout ),
	.cin(gnd),
	.combout(Selector16),
	.cout());
// synopsys translate_off
defparam \Selector16~11 .lut_mask = 16'hFFF8;
defparam \Selector16~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N0
cycloneive_lcell_comb \Selector17~7 (
// Equation(s):
// Selector17 = (\Selector17~6_combout ) # ((\ShiftRight0~123_combout  & (\Selector20~0_combout  & !\Mux33~3_combout )))

	.dataa(\ShiftRight0~123_combout ),
	.datab(\Selector20~0_combout ),
	.datac(Mux33),
	.datad(\Selector17~6_combout ),
	.cin(gnd),
	.combout(Selector17),
	.cout());
// synopsys translate_off
defparam \Selector17~7 .lut_mask = 16'hFF08;
defparam \Selector17~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N2
cycloneive_lcell_comb \Equal10~7 (
// Equation(s):
// Equal101 = (!Selector16 & (!Selector15 & (!Selector14 & !Selector17)))

	.dataa(Selector16),
	.datab(Selector15),
	.datac(Selector14),
	.datad(Selector17),
	.cin(gnd),
	.combout(Equal101),
	.cout());
// synopsys translate_off
defparam \Equal10~7 .lut_mask = 16'h0001;
defparam \Equal10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N22
cycloneive_lcell_comb \Selector20~9 (
// Equation(s):
// Selector20 = (\Selector20~2_combout ) # ((\Selector20~8_combout ) # ((\ShiftRight0~108_combout  & \Selector16~10_combout )))

	.dataa(\ShiftRight0~108_combout ),
	.datab(\Selector16~10_combout ),
	.datac(\Selector20~2_combout ),
	.datad(\Selector20~8_combout ),
	.cin(gnd),
	.combout(Selector20),
	.cout());
// synopsys translate_off
defparam \Selector20~9 .lut_mask = 16'hFFF8;
defparam \Selector20~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N28
cycloneive_lcell_comb \Selector21~8 (
// Equation(s):
// Selector21 = (\Selector21~7_combout ) # ((\Selector21~1_combout ) # ((\ShiftRight0~112_combout  & \Selector16~10_combout )))

	.dataa(\Selector21~7_combout ),
	.datab(\ShiftRight0~112_combout ),
	.datac(\Selector21~1_combout ),
	.datad(\Selector16~10_combout ),
	.cin(gnd),
	.combout(Selector21),
	.cout());
// synopsys translate_off
defparam \Selector21~8 .lut_mask = 16'hFEFA;
defparam \Selector21~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N22
cycloneive_lcell_comb \Selector18~7 (
// Equation(s):
// Selector18 = (\Selector18~6_combout ) # ((\ShiftRight0~107_combout  & (\ShiftRight0~75_combout  & \Selector20~0_combout )))

	.dataa(\ShiftRight0~107_combout ),
	.datab(\ShiftRight0~75_combout ),
	.datac(\Selector20~0_combout ),
	.datad(\Selector18~6_combout ),
	.cin(gnd),
	.combout(Selector18),
	.cout());
// synopsys translate_off
defparam \Selector18~7 .lut_mask = 16'hFF80;
defparam \Selector18~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N28
cycloneive_lcell_comb \Selector19~7 (
// Equation(s):
// Selector19 = (\Selector19~6_combout ) # ((\Selector20~0_combout  & (\ShiftRight0~107_combout  & \ShiftRight0~137_combout )))

	.dataa(\Selector20~0_combout ),
	.datab(\ShiftRight0~107_combout ),
	.datac(\ShiftRight0~137_combout ),
	.datad(\Selector19~6_combout ),
	.cin(gnd),
	.combout(Selector19),
	.cout());
// synopsys translate_off
defparam \Selector19~7 .lut_mask = 16'hFF80;
defparam \Selector19~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N8
cycloneive_lcell_comb \Selector8~2 (
// Equation(s):
// Selector8 = (!\Mux33~3_combout  & (ShiftLeft0 & \Selector0~29_combout ))

	.dataa(gnd),
	.datab(Mux33),
	.datac(ShiftLeft0),
	.datad(\Selector0~29_combout ),
	.cin(gnd),
	.combout(Selector8),
	.cout());
// synopsys translate_off
defparam \Selector8~2 .lut_mask = 16'h3000;
defparam \Selector8~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N8
cycloneive_lcell_comb \Selector8~3 (
// Equation(s):
// Selector81 = (\Selector16~1_combout  & (!cuifaluOp_0 & \Selector0~28_combout ))

	.dataa(\Selector16~1_combout ),
	.datab(cuifaluOp_0),
	.datac(gnd),
	.datad(\Selector0~28_combout ),
	.cin(gnd),
	.combout(Selector81),
	.cout());
// synopsys translate_off
defparam \Selector8~3 .lut_mask = 16'h2200;
defparam \Selector8~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N26
cycloneive_lcell_comb \Selector8~10 (
// Equation(s):
// Selector82 = (\Selector8~9_combout ) # ((\Selector0~27_combout  & \Selector8~1_combout ))

	.dataa(\Selector0~27_combout ),
	.datab(gnd),
	.datac(\Selector8~1_combout ),
	.datad(\Selector8~9_combout ),
	.cin(gnd),
	.combout(Selector82),
	.cout());
// synopsys translate_off
defparam \Selector8~10 .lut_mask = 16'hFFA0;
defparam \Selector8~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N28
cycloneive_lcell_comb \Selector9~9 (
// Equation(s):
// Selector9 = (\Selector9~8_combout ) # ((!\Mux33~3_combout  & (ShiftLeft03 & \Selector0~29_combout )))

	.dataa(Mux33),
	.datab(ShiftLeft03),
	.datac(\Selector0~29_combout ),
	.datad(\Selector9~8_combout ),
	.cin(gnd),
	.combout(Selector9),
	.cout());
// synopsys translate_off
defparam \Selector9~9 .lut_mask = 16'hFF40;
defparam \Selector9~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N14
cycloneive_lcell_comb \Selector31~9 (
// Equation(s):
// Selector312 = (Selector31) # ((Mux31 & Selector311))

	.dataa(gnd),
	.datab(Mux311),
	.datac(Selector311),
	.datad(Selector31),
	.cin(gnd),
	.combout(Selector312),
	.cout());
// synopsys translate_off
defparam \Selector31~9 .lut_mask = 16'hFFC0;
defparam \Selector31~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N4
cycloneive_lcell_comb \Selector22~8 (
// Equation(s):
// Selector22 = (\Selector22~7_combout ) # ((\Selector22~1_combout ) # ((\ShiftRight0~72_combout  & \Selector16~10_combout )))

	.dataa(\ShiftRight0~72_combout ),
	.datab(\Selector16~10_combout ),
	.datac(\Selector22~7_combout ),
	.datad(\Selector22~1_combout ),
	.cin(gnd),
	.combout(Selector22),
	.cout());
// synopsys translate_off
defparam \Selector22~8 .lut_mask = 16'hFFF8;
defparam \Selector22~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N16
cycloneive_lcell_comb \Selector23~8 (
// Equation(s):
// Selector23 = (\Selector23~1_combout ) # ((\Selector23~7_combout ) # ((\ShiftRight0~94_combout  & \Selector16~10_combout )))

	.dataa(\ShiftRight0~94_combout ),
	.datab(\Selector23~1_combout ),
	.datac(\Selector16~10_combout ),
	.datad(\Selector23~7_combout ),
	.cin(gnd),
	.combout(Selector23),
	.cout());
// synopsys translate_off
defparam \Selector23~8 .lut_mask = 16'hFFEC;
defparam \Selector23~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N4
cycloneive_lcell_comb \Equal10~9 (
// Equation(s):
// Equal102 = (!Selector22 & (!Selector312 & (\Equal10~8_combout  & !Selector23)))

	.dataa(Selector22),
	.datab(Selector312),
	.datac(\Equal10~8_combout ),
	.datad(Selector23),
	.cin(gnd),
	.combout(Equal102),
	.cout());
// synopsys translate_off
defparam \Equal10~9 .lut_mask = 16'h0010;
defparam \Equal10~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N16
cycloneive_lcell_comb \Selector8~11 (
// Equation(s):
// Selector83 = (Selector8) # ((Selector82) # (Selector81))

	.dataa(Selector8),
	.datab(gnd),
	.datac(Selector82),
	.datad(Selector81),
	.cin(gnd),
	.combout(Selector83),
	.cout());
// synopsys translate_off
defparam \Selector8~11 .lut_mask = 16'hFFFA;
defparam \Selector8~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N2
cycloneive_lcell_comb \Selector0~9 (
// Equation(s):
// \Selector0~9_combout  = (!cuifaluOp_0 & (!cuifaluOp_31 & (!cuifaluOp_1 & !cuifaluOp_2)))

	.dataa(cuifaluOp_0),
	.datab(cuifaluOp_3),
	.datac(cuifaluOp_1),
	.datad(cuifaluOp_2),
	.cin(gnd),
	.combout(\Selector0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~9 .lut_mask = 16'h0001;
defparam \Selector0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N12
cycloneive_lcell_comb \Selector30~3 (
// Equation(s):
// \Selector30~3_combout  = (\Mux35~4_combout  & ((\Selector0~8_combout ) # ((\Selector0~9_combout  & Mux30))))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~9_combout ),
	.datac(Mux301),
	.datad(Mux352),
	.cin(gnd),
	.combout(\Selector30~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~3 .lut_mask = 16'hEA00;
defparam \Selector30~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N28
cycloneive_lcell_comb \Selector0~10 (
// Equation(s):
// \Selector0~10_combout  = (cuifaluOp_1 & (!cuifaluOp_31 & (!cuifaluOp_0 & !cuifaluOp_2)))

	.dataa(cuifaluOp_1),
	.datab(cuifaluOp_3),
	.datac(cuifaluOp_0),
	.datad(cuifaluOp_2),
	.cin(gnd),
	.combout(\Selector0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~10 .lut_mask = 16'h0002;
defparam \Selector0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N22
cycloneive_lcell_comb \Selector30~4 (
// Equation(s):
// \Selector30~4_combout  = (\Selector30~3_combout ) # ((\Selector0~10_combout  & (Mux30 $ (\Mux35~4_combout ))))

	.dataa(\Selector30~3_combout ),
	.datab(\Selector0~10_combout ),
	.datac(Mux301),
	.datad(Mux352),
	.cin(gnd),
	.combout(\Selector30~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~4 .lut_mask = 16'hAEEA;
defparam \Selector30~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N8
cycloneive_lcell_comb \Selector0~8 (
// Equation(s):
// \Selector0~8_combout  = (cuifaluOp_0 & (!cuifaluOp_31 & (!cuifaluOp_1 & !cuifaluOp_2)))

	.dataa(cuifaluOp_0),
	.datab(cuifaluOp_3),
	.datac(cuifaluOp_1),
	.datad(cuifaluOp_2),
	.cin(gnd),
	.combout(\Selector0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~8 .lut_mask = 16'h0002;
defparam \Selector0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N16
cycloneive_lcell_comb \Selector0~12 (
// Equation(s):
// \Selector0~12_combout  = (cuifaluOp_0 & (!cuifaluOp_31 & (cuifaluOp_1 & cuifaluOp_2)))

	.dataa(cuifaluOp_0),
	.datab(cuifaluOp_3),
	.datac(cuifaluOp_1),
	.datad(cuifaluOp_2),
	.cin(gnd),
	.combout(\Selector0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~12 .lut_mask = 16'h2000;
defparam \Selector0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N0
cycloneive_lcell_comb \Add1~0 (
// Equation(s):
// \Add1~0_combout  = (Mux31 & ((GND) # (!\Mux36~4_combout ))) # (!Mux31 & (\Mux36~4_combout  $ (GND)))
// \Add1~1  = CARRY((Mux31) # (!\Mux36~4_combout ))

	.dataa(Mux311),
	.datab(Mux36),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h66BB;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N2
cycloneive_lcell_comb \Add1~2 (
// Equation(s):
// \Add1~2_combout  = (\Mux35~4_combout  & ((Mux30 & (!\Add1~1 )) # (!Mux30 & ((\Add1~1 ) # (GND))))) # (!\Mux35~4_combout  & ((Mux30 & (\Add1~1  & VCC)) # (!Mux30 & (!\Add1~1 ))))
// \Add1~3  = CARRY((\Mux35~4_combout  & ((!\Add1~1 ) # (!Mux30))) # (!\Mux35~4_combout  & (!Mux30 & !\Add1~1 )))

	.dataa(Mux352),
	.datab(Mux301),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h692B;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N0
cycloneive_lcell_comb \Add0~0 (
// Equation(s):
// \Add0~0_combout  = (\Mux36~4_combout  & (Mux31 $ (VCC))) # (!\Mux36~4_combout  & (Mux31 & VCC))
// \Add0~1  = CARRY((\Mux36~4_combout  & Mux31))

	.dataa(Mux36),
	.datab(Mux311),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
// synopsys translate_off
defparam \Add0~0 .lut_mask = 16'h6688;
defparam \Add0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N2
cycloneive_lcell_comb \Add0~2 (
// Equation(s):
// \Add0~2_combout  = (Mux30 & ((\Mux35~4_combout  & (\Add0~1  & VCC)) # (!\Mux35~4_combout  & (!\Add0~1 )))) # (!Mux30 & ((\Mux35~4_combout  & (!\Add0~1 )) # (!\Mux35~4_combout  & ((\Add0~1 ) # (GND)))))
// \Add0~3  = CARRY((Mux30 & (!\Mux35~4_combout  & !\Add0~1 )) # (!Mux30 & ((!\Add0~1 ) # (!\Mux35~4_combout ))))

	.dataa(Mux301),
	.datab(Mux352),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
// synopsys translate_off
defparam \Add0~2 .lut_mask = 16'h9617;
defparam \Add0~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N14
cycloneive_lcell_comb \Selector30~6 (
// Equation(s):
// \Selector30~6_combout  = (\Selector0~13_combout  & ((\Add0~2_combout ) # ((\Selector0~12_combout  & \Add1~2_combout )))) # (!\Selector0~13_combout  & (\Selector0~12_combout  & (\Add1~2_combout )))

	.dataa(\Selector0~13_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Add1~2_combout ),
	.datad(\Add0~2_combout ),
	.cin(gnd),
	.combout(\Selector30~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~6 .lut_mask = 16'hEAC0;
defparam \Selector30~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N30
cycloneive_lcell_comb \Selector0~11 (
// Equation(s):
// \Selector0~11_combout  = (cuifaluOp_0 & (!cuifaluOp_31 & (cuifaluOp_1 & !cuifaluOp_2)))

	.dataa(cuifaluOp_0),
	.datab(cuifaluOp_3),
	.datac(cuifaluOp_1),
	.datad(cuifaluOp_2),
	.cin(gnd),
	.combout(\Selector0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~11 .lut_mask = 16'h0020;
defparam \Selector0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N0
cycloneive_lcell_comb \Selector30~5 (
// Equation(s):
// \Selector30~5_combout  = (!\Mux35~2_combout  & (!Mux30 & (\Selector0~11_combout  & !\Mux35~3_combout )))

	.dataa(Mux35),
	.datab(Mux301),
	.datac(\Selector0~11_combout ),
	.datad(Mux351),
	.cin(gnd),
	.combout(\Selector30~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~5 .lut_mask = 16'h0010;
defparam \Selector30~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N4
cycloneive_lcell_comb \Selector30~7 (
// Equation(s):
// \Selector30~7_combout  = (\Selector30~6_combout ) # ((\Selector30~5_combout ) # ((\Selector0~8_combout  & Mux30)))

	.dataa(\Selector0~8_combout ),
	.datab(Mux301),
	.datac(\Selector30~6_combout ),
	.datad(\Selector30~5_combout ),
	.cin(gnd),
	.combout(\Selector30~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~7 .lut_mask = 16'hFFF8;
defparam \Selector30~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N2
cycloneive_lcell_comb \ShiftRight0~71 (
// Equation(s):
// \ShiftRight0~71_combout  = (\Mux36~4_combout  & (Mux21)) # (!\Mux36~4_combout  & ((Mux22)))

	.dataa(gnd),
	.datab(Mux36),
	.datac(Mux211),
	.datad(Mux221),
	.cin(gnd),
	.combout(\ShiftRight0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~71 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N12
cycloneive_lcell_comb \ShiftRight0~70 (
// Equation(s):
// \ShiftRight0~70_combout  = (\Mux36~4_combout  & (Mux19)) # (!\Mux36~4_combout  & ((Mux20)))

	.dataa(Mux191),
	.datab(gnd),
	.datac(Mux201),
	.datad(Mux36),
	.cin(gnd),
	.combout(\ShiftRight0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~70 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N30
cycloneive_lcell_comb \ShiftRight0~130 (
// Equation(s):
// \ShiftRight0~130_combout  = (\Mux35~3_combout  & (((\ShiftRight0~70_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftRight0~70_combout ))) # (!\Mux35~2_combout  & (\ShiftRight0~71_combout ))))

	.dataa(Mux351),
	.datab(\ShiftRight0~71_combout ),
	.datac(Mux35),
	.datad(\ShiftRight0~70_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~130_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~130 .lut_mask = 16'hFE04;
defparam \ShiftRight0~130 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N6
cycloneive_lcell_comb \ShiftRight0~68 (
// Equation(s):
// \ShiftRight0~68_combout  = (\Mux36~4_combout  & ((Mux15))) # (!\Mux36~4_combout  & (Mux16))

	.dataa(Mux161),
	.datab(Mux152),
	.datac(gnd),
	.datad(Mux36),
	.cin(gnd),
	.combout(\ShiftRight0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~68 .lut_mask = 16'hCCAA;
defparam \ShiftRight0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N16
cycloneive_lcell_comb \ShiftRight0~69 (
// Equation(s):
// \ShiftRight0~69_combout  = (\Mux36~4_combout  & (Mux17)) # (!\Mux36~4_combout  & ((Mux18)))

	.dataa(Mux171),
	.datab(gnd),
	.datac(Mux181),
	.datad(Mux36),
	.cin(gnd),
	.combout(\ShiftRight0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~69 .lut_mask = 16'hAAF0;
defparam \ShiftRight0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N22
cycloneive_lcell_comb \ShiftRight0~129 (
// Equation(s):
// \ShiftRight0~129_combout  = (\Mux35~3_combout  & (((\ShiftRight0~68_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & (\ShiftRight0~68_combout )) # (!\Mux35~2_combout  & ((\ShiftRight0~69_combout )))))

	.dataa(Mux351),
	.datab(Mux35),
	.datac(\ShiftRight0~68_combout ),
	.datad(\ShiftRight0~69_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~129_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~129 .lut_mask = 16'hF1E0;
defparam \ShiftRight0~129 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N12
cycloneive_lcell_comb \ShiftRight0~72 (
// Equation(s):
// \ShiftRight0~72_combout  = (\Mux34~3_combout  & ((\ShiftRight0~129_combout ))) # (!\Mux34~3_combout  & (\ShiftRight0~130_combout ))

	.dataa(gnd),
	.datab(Mux34),
	.datac(\ShiftRight0~130_combout ),
	.datad(\ShiftRight0~129_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~72 .lut_mask = 16'hFC30;
defparam \ShiftRight0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N4
cycloneive_lcell_comb \ShiftRight0~62 (
// Equation(s):
// \ShiftRight0~62_combout  = (!\Mux35~4_combout  & ((\Mux36~4_combout  & ((Mux29))) # (!\Mux36~4_combout  & (Mux30))))

	.dataa(Mux36),
	.datab(Mux352),
	.datac(Mux301),
	.datad(Mux291),
	.cin(gnd),
	.combout(\ShiftRight0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~62 .lut_mask = 16'h3210;
defparam \ShiftRight0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N30
cycloneive_lcell_comb \ShiftRight0~64 (
// Equation(s):
// \ShiftRight0~64_combout  = (!\Mux34~3_combout  & ((\ShiftRight0~62_combout ) # ((\ShiftRight0~63_combout  & \Mux35~4_combout ))))

	.dataa(\ShiftRight0~63_combout ),
	.datab(Mux34),
	.datac(\ShiftRight0~62_combout ),
	.datad(Mux352),
	.cin(gnd),
	.combout(\ShiftRight0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~64 .lut_mask = 16'h3230;
defparam \ShiftRight0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N22
cycloneive_lcell_comb \ShiftRight0~66 (
// Equation(s):
// \ShiftRight0~66_combout  = (\Mux36~4_combout  & ((Mux25))) # (!\Mux36~4_combout  & (Mux26))

	.dataa(gnd),
	.datab(Mux261),
	.datac(Mux36),
	.datad(Mux251),
	.cin(gnd),
	.combout(\ShiftRight0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~66 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N0
cycloneive_lcell_comb \ShiftRight0~65 (
// Equation(s):
// \ShiftRight0~65_combout  = (\Mux36~4_combout  & ((Mux23))) # (!\Mux36~4_combout  & (Mux24))

	.dataa(gnd),
	.datab(Mux36),
	.datac(Mux241),
	.datad(Mux231),
	.cin(gnd),
	.combout(\ShiftRight0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~65 .lut_mask = 16'hFC30;
defparam \ShiftRight0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N4
cycloneive_lcell_comb \ShiftRight0~128 (
// Equation(s):
// \ShiftRight0~128_combout  = (\Mux35~2_combout  & (((\ShiftRight0~65_combout )))) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & ((\ShiftRight0~65_combout ))) # (!\Mux35~3_combout  & (\ShiftRight0~66_combout ))))

	.dataa(Mux35),
	.datab(Mux351),
	.datac(\ShiftRight0~66_combout ),
	.datad(\ShiftRight0~65_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~128_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~128 .lut_mask = 16'hFE10;
defparam \ShiftRight0~128 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N24
cycloneive_lcell_comb \ShiftRight0~67 (
// Equation(s):
// \ShiftRight0~67_combout  = (!\Mux33~3_combout  & ((\ShiftRight0~64_combout ) # ((\Mux34~3_combout  & \ShiftRight0~128_combout ))))

	.dataa(Mux33),
	.datab(Mux34),
	.datac(\ShiftRight0~64_combout ),
	.datad(\ShiftRight0~128_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~67 .lut_mask = 16'h5450;
defparam \ShiftRight0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N10
cycloneive_lcell_comb \ShiftRight0~73 (
// Equation(s):
// \ShiftRight0~73_combout  = (!\Mux32~4_combout  & ((\ShiftRight0~67_combout ) # ((\Mux33~3_combout  & \ShiftRight0~72_combout ))))

	.dataa(Mux33),
	.datab(Mux32),
	.datac(\ShiftRight0~72_combout ),
	.datad(\ShiftRight0~67_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~73 .lut_mask = 16'h3320;
defparam \ShiftRight0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N6
cycloneive_lcell_comb \ShiftRight0~77 (
// Equation(s):
// \ShiftRight0~77_combout  = (\Mux36~4_combout  & ((Mux5))) # (!\Mux36~4_combout  & (Mux6))

	.dataa(gnd),
	.datab(Mux61),
	.datac(Mux36),
	.datad(Mux52),
	.cin(gnd),
	.combout(\ShiftRight0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~77 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N28
cycloneive_lcell_comb \ShiftRight0~76 (
// Equation(s):
// \ShiftRight0~76_combout  = (\Mux36~4_combout  & (Mux3)) # (!\Mux36~4_combout  & ((Mux4)))

	.dataa(Mux36),
	.datab(gnd),
	.datac(Mux3),
	.datad(Mux4),
	.cin(gnd),
	.combout(\ShiftRight0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~76 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N16
cycloneive_lcell_comb \ShiftRight0~131 (
// Equation(s):
// \ShiftRight0~131_combout  = (\Mux35~3_combout  & (((\ShiftRight0~76_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftRight0~76_combout ))) # (!\Mux35~2_combout  & (\ShiftRight0~77_combout ))))

	.dataa(Mux351),
	.datab(Mux35),
	.datac(\ShiftRight0~77_combout ),
	.datad(\ShiftRight0~76_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~131_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~131 .lut_mask = 16'hFE10;
defparam \ShiftRight0~131 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N20
cycloneive_lcell_comb \ShiftRight0~74 (
// Equation(s):
// \ShiftRight0~74_combout  = (!\Mux36~4_combout  & ((\Mux35~4_combout  & ((Mux0))) # (!\Mux35~4_combout  & (Mux2))))

	.dataa(Mux2),
	.datab(Mux36),
	.datac(Mux0),
	.datad(Mux352),
	.cin(gnd),
	.combout(\ShiftRight0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~74 .lut_mask = 16'h3022;
defparam \ShiftRight0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N18
cycloneive_lcell_comb \ShiftRight0~75 (
// Equation(s):
// \ShiftRight0~75_combout  = (\ShiftRight0~74_combout ) # ((\Mux36~4_combout  & (!\Mux35~4_combout  & Mux1)))

	.dataa(Mux36),
	.datab(Mux352),
	.datac(Mux1),
	.datad(\ShiftRight0~74_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~75 .lut_mask = 16'hFF20;
defparam \ShiftRight0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N30
cycloneive_lcell_comb \ShiftRight0~78 (
// Equation(s):
// \ShiftRight0~78_combout  = (\Mux34~3_combout  & ((\ShiftRight0~75_combout ))) # (!\Mux34~3_combout  & (\ShiftRight0~131_combout ))

	.dataa(Mux34),
	.datab(gnd),
	.datac(\ShiftRight0~131_combout ),
	.datad(\ShiftRight0~75_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~78 .lut_mask = 16'hFA50;
defparam \ShiftRight0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N30
cycloneive_lcell_comb \ShiftRight0~79 (
// Equation(s):
// \ShiftRight0~79_combout  = (\Mux36~4_combout  & ((Mux7))) # (!\Mux36~4_combout  & (Mux8))

	.dataa(Mux36),
	.datab(gnd),
	.datac(Mux81),
	.datad(Mux71),
	.cin(gnd),
	.combout(\ShiftRight0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~79 .lut_mask = 16'hFA50;
defparam \ShiftRight0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N20
cycloneive_lcell_comb \ShiftRight0~80 (
// Equation(s):
// \ShiftRight0~80_combout  = (\Mux36~4_combout  & (Mux9)) # (!\Mux36~4_combout  & ((Mux10)))

	.dataa(Mux36),
	.datab(gnd),
	.datac(Mux91),
	.datad(Mux101),
	.cin(gnd),
	.combout(\ShiftRight0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~80 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N26
cycloneive_lcell_comb \ShiftRight0~132 (
// Equation(s):
// \ShiftRight0~132_combout  = (\Mux35~3_combout  & (((\ShiftRight0~79_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & (\ShiftRight0~79_combout )) # (!\Mux35~2_combout  & ((\ShiftRight0~80_combout )))))

	.dataa(Mux351),
	.datab(Mux35),
	.datac(\ShiftRight0~79_combout ),
	.datad(\ShiftRight0~80_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~132_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~132 .lut_mask = 16'hF1E0;
defparam \ShiftRight0~132 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N12
cycloneive_lcell_comb \ShiftRight0~82 (
// Equation(s):
// \ShiftRight0~82_combout  = (\Mux36~4_combout  & (Mux13)) # (!\Mux36~4_combout  & ((Mux14)))

	.dataa(gnd),
	.datab(Mux131),
	.datac(Mux36),
	.datad(Mux141),
	.cin(gnd),
	.combout(\ShiftRight0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~82 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N16
cycloneive_lcell_comb \ShiftRight0~133 (
// Equation(s):
// \ShiftRight0~133_combout  = (\Mux35~3_combout  & (\ShiftRight0~81_combout )) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & (\ShiftRight0~81_combout )) # (!\Mux35~2_combout  & ((\ShiftRight0~82_combout )))))

	.dataa(\ShiftRight0~81_combout ),
	.datab(Mux351),
	.datac(\ShiftRight0~82_combout ),
	.datad(Mux35),
	.cin(gnd),
	.combout(\ShiftRight0~133_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~133 .lut_mask = 16'hAAB8;
defparam \ShiftRight0~133 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N12
cycloneive_lcell_comb \Selector22~0 (
// Equation(s):
// \Selector22~0_combout  = (\Mux34~3_combout  & (\ShiftRight0~132_combout )) # (!\Mux34~3_combout  & ((\ShiftRight0~133_combout )))

	.dataa(gnd),
	.datab(Mux34),
	.datac(\ShiftRight0~132_combout ),
	.datad(\ShiftRight0~133_combout ),
	.cin(gnd),
	.combout(\Selector22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~0 .lut_mask = 16'hF3C0;
defparam \Selector22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N8
cycloneive_lcell_comb \ShiftRight0~83 (
// Equation(s):
// \ShiftRight0~83_combout  = (\Mux33~3_combout  & (\ShiftRight0~78_combout )) # (!\Mux33~3_combout  & ((\Selector22~0_combout )))

	.dataa(Mux33),
	.datab(gnd),
	.datac(\ShiftRight0~78_combout ),
	.datad(\Selector22~0_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~83 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N28
cycloneive_lcell_comb \Selector0~6 (
// Equation(s):
// \Selector0~6_combout  = (cuifaluOp_2 & (cuifaluOp_0 & (!cuifaluOp_31 & !cuifaluOp_1)))

	.dataa(cuifaluOp_2),
	.datab(cuifaluOp_0),
	.datac(cuifaluOp_3),
	.datad(cuifaluOp_1),
	.cin(gnd),
	.combout(\Selector0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~6 .lut_mask = 16'h0008;
defparam \Selector0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N18
cycloneive_lcell_comb \Selector24~0 (
// Equation(s):
// \Selector24~0_combout  = (!\ShiftRight0~61_combout  & \Selector0~6_combout )

	.dataa(\ShiftRight0~61_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\Selector0~6_combout ),
	.cin(gnd),
	.combout(\Selector24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~0 .lut_mask = 16'h5500;
defparam \Selector24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N22
cycloneive_lcell_comb \Selector30~0 (
// Equation(s):
// \Selector30~0_combout  = (\Selector24~0_combout  & ((\ShiftRight0~73_combout ) # ((\Mux32~4_combout  & \ShiftRight0~83_combout ))))

	.dataa(\ShiftRight0~73_combout ),
	.datab(Mux32),
	.datac(\ShiftRight0~83_combout ),
	.datad(\Selector24~0_combout ),
	.cin(gnd),
	.combout(\Selector30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~0 .lut_mask = 16'hEA00;
defparam \Selector30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N30
cycloneive_lcell_comb \ShiftLeft0~52 (
// Equation(s):
// \ShiftLeft0~52_combout  = (\Mux36~4_combout  & ((Mux31))) # (!\Mux36~4_combout  & (Mux30))

	.dataa(gnd),
	.datab(Mux301),
	.datac(Mux36),
	.datad(Mux311),
	.cin(gnd),
	.combout(\ShiftLeft0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~52 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N16
cycloneive_lcell_comb \Selector30~1 (
// Equation(s):
// \Selector30~1_combout  = (!\Mux33~3_combout  & (!\Mux35~4_combout  & (\ShiftLeft0~52_combout  & !\Mux34~3_combout )))

	.dataa(Mux33),
	.datab(Mux352),
	.datac(\ShiftLeft0~52_combout ),
	.datad(Mux34),
	.cin(gnd),
	.combout(\Selector30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~1 .lut_mask = 16'h0010;
defparam \Selector30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N28
cycloneive_lcell_comb \Selector0~7 (
// Equation(s):
// \Selector0~7_combout  = (!cuifaluOp_0 & (!cuifaluOp_1 & (!cuifaluOp_31 & cuifaluOp_2)))

	.dataa(cuifaluOp_0),
	.datab(cuifaluOp_1),
	.datac(cuifaluOp_3),
	.datad(cuifaluOp_2),
	.cin(gnd),
	.combout(\Selector0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~7 .lut_mask = 16'h0100;
defparam \Selector0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N20
cycloneive_lcell_comb \ShiftRight0~53 (
// Equation(s):
// \ShiftRight0~53_combout  = (\Mux9~0_combout ) # ((\Mux5~1_combout ) # ((\Mux8~0_combout ) # (\Mux10~0_combout )))

	.dataa(Mux9),
	.datab(Mux5),
	.datac(Mux8),
	.datad(Mux10),
	.cin(gnd),
	.combout(\ShiftRight0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~53 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N8
cycloneive_lcell_comb \ShiftRight0~54 (
// Equation(s):
// \ShiftRight0~54_combout  = (\Mux13~0_combout ) # ((\Mux11~0_combout ) # ((\Mux5~1_combout ) # (\Mux12~1_combout )))

	.dataa(Mux13),
	.datab(Mux11),
	.datac(Mux5),
	.datad(Mux12),
	.cin(gnd),
	.combout(\ShiftRight0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~54 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N14
cycloneive_lcell_comb \ShiftRight0~55 (
// Equation(s):
// \ShiftRight0~55_combout  = (\Mux16~1_combout ) # ((\ShiftRight0~54_combout ) # ((\Mux14~1_combout ) # (\Mux15~1_combout )))

	.dataa(Mux16),
	.datab(\ShiftRight0~54_combout ),
	.datac(Mux14),
	.datad(Mux151),
	.cin(gnd),
	.combout(\ShiftRight0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~55 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N18
cycloneive_lcell_comb \ShiftRight0~56 (
// Equation(s):
// \ShiftRight0~56_combout  = (\Mux5~1_combout ) # ((\Mux19~0_combout ) # ((\Mux18~0_combout ) # (\Mux17~0_combout )))

	.dataa(Mux5),
	.datab(Mux19),
	.datac(Mux18),
	.datad(Mux17),
	.cin(gnd),
	.combout(\ShiftRight0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~56 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N4
cycloneive_lcell_comb \ShiftRight0~57 (
// Equation(s):
// \ShiftRight0~57_combout  = (\Mux21~1_combout ) # ((\ShiftRight0~56_combout ) # ((\Mux22~1_combout ) # (\Mux20~1_combout )))

	.dataa(Mux21),
	.datab(\ShiftRight0~56_combout ),
	.datac(Mux22),
	.datad(Mux20),
	.cin(gnd),
	.combout(\ShiftRight0~57_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~57 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N4
cycloneive_lcell_comb \ShiftRight0~59 (
// Equation(s):
// \ShiftRight0~59_combout  = (\Mux30~1_combout ) # ((\Mux27~1_combout ) # ((\Mux28~1_combout ) # (\Mux29~1_combout )))

	.dataa(Mux30),
	.datab(Mux27),
	.datac(Mux28),
	.datad(Mux29),
	.cin(gnd),
	.combout(\ShiftRight0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~59 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N10
cycloneive_lcell_comb \ShiftRight0~58 (
// Equation(s):
// \ShiftRight0~58_combout  = (\Mux23~1_combout ) # ((\Mux25~1_combout ) # ((\Mux24~1_combout ) # (\Mux26~1_combout )))

	.dataa(Mux23),
	.datab(Mux25),
	.datac(Mux24),
	.datad(Mux26),
	.cin(gnd),
	.combout(\ShiftRight0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~58 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N18
cycloneive_lcell_comb \ShiftRight0~60 (
// Equation(s):
// \ShiftRight0~60_combout  = (\Mux31~1_combout ) # ((\ShiftRight0~57_combout ) # ((\ShiftRight0~59_combout ) # (\ShiftRight0~58_combout )))

	.dataa(Mux31),
	.datab(\ShiftRight0~57_combout ),
	.datac(\ShiftRight0~59_combout ),
	.datad(\ShiftRight0~58_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~60 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N24
cycloneive_lcell_comb \ShiftRight0~61 (
// Equation(s):
// \ShiftRight0~61_combout  = (\ShiftRight0~52_combout ) # ((\ShiftRight0~53_combout ) # ((\ShiftRight0~55_combout ) # (\ShiftRight0~60_combout )))

	.dataa(\ShiftRight0~52_combout ),
	.datab(\ShiftRight0~53_combout ),
	.datac(\ShiftRight0~55_combout ),
	.datad(\ShiftRight0~60_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~61 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y36_N16
cycloneive_lcell_comb \Selector30~2 (
// Equation(s):
// \Selector30~2_combout  = (\Selector30~1_combout  & (\Selector0~7_combout  & (!\ShiftRight0~61_combout  & !\Mux32~4_combout )))

	.dataa(\Selector30~1_combout ),
	.datab(\Selector0~7_combout ),
	.datac(\ShiftRight0~61_combout ),
	.datad(Mux32),
	.cin(gnd),
	.combout(\Selector30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector30~2 .lut_mask = 16'h0008;
defparam \Selector30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N2
cycloneive_lcell_comb \ShiftRight0~96 (
// Equation(s):
// \ShiftRight0~96_combout  = (\Mux36~4_combout  & (Mux0)) # (!\Mux36~4_combout  & ((Mux1)))

	.dataa(gnd),
	.datab(Mux0),
	.datac(Mux1),
	.datad(Mux36),
	.cin(gnd),
	.combout(\ShiftRight0~96_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~96 .lut_mask = 16'hCCF0;
defparam \ShiftRight0~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N20
cycloneive_lcell_comb \ShiftRight0~97 (
// Equation(s):
// \ShiftRight0~97_combout  = (\Mux36~4_combout  & ((Mux2))) # (!\Mux36~4_combout  & (Mux3))

	.dataa(gnd),
	.datab(Mux36),
	.datac(Mux3),
	.datad(Mux2),
	.cin(gnd),
	.combout(\ShiftRight0~97_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~97 .lut_mask = 16'hFC30;
defparam \ShiftRight0~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N30
cycloneive_lcell_comb \ShiftRight0~137 (
// Equation(s):
// \ShiftRight0~137_combout  = (\Mux35~3_combout  & (((\ShiftRight0~96_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & (\ShiftRight0~96_combout )) # (!\Mux35~2_combout  & ((\ShiftRight0~97_combout )))))

	.dataa(Mux351),
	.datab(Mux35),
	.datac(\ShiftRight0~96_combout ),
	.datad(\ShiftRight0~97_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~137_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~137 .lut_mask = 16'hF1E0;
defparam \ShiftRight0~137 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N14
cycloneive_lcell_comb \ShiftRight0~98 (
// Equation(s):
// \ShiftRight0~98_combout  = (\Mux36~4_combout  & ((Mux4))) # (!\Mux36~4_combout  & (Mux5))

	.dataa(gnd),
	.datab(Mux36),
	.datac(Mux52),
	.datad(Mux4),
	.cin(gnd),
	.combout(\ShiftRight0~98_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~98 .lut_mask = 16'hFC30;
defparam \ShiftRight0~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N16
cycloneive_lcell_comb \ShiftRight0~99 (
// Equation(s):
// \ShiftRight0~99_combout  = (\Mux36~4_combout  & (Mux6)) # (!\Mux36~4_combout  & ((Mux7)))

	.dataa(gnd),
	.datab(Mux36),
	.datac(Mux61),
	.datad(Mux71),
	.cin(gnd),
	.combout(\ShiftRight0~99_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~99 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N12
cycloneive_lcell_comb \ShiftRight0~138 (
// Equation(s):
// \ShiftRight0~138_combout  = (\Mux35~3_combout  & (\ShiftRight0~98_combout )) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & (\ShiftRight0~98_combout )) # (!\Mux35~2_combout  & ((\ShiftRight0~99_combout )))))

	.dataa(Mux351),
	.datab(\ShiftRight0~98_combout ),
	.datac(Mux35),
	.datad(\ShiftRight0~99_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~138_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~138 .lut_mask = 16'hCDC8;
defparam \ShiftRight0~138 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N28
cycloneive_lcell_comb \ShiftRight0~90 (
// Equation(s):
// \ShiftRight0~90_combout  = (\Mux36~4_combout  & (Mux16)) # (!\Mux36~4_combout  & ((Mux17)))

	.dataa(Mux161),
	.datab(gnd),
	.datac(Mux36),
	.datad(Mux171),
	.cin(gnd),
	.combout(\ShiftRight0~90_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~90 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N26
cycloneive_lcell_comb \ShiftRight0~91 (
// Equation(s):
// \ShiftRight0~91_combout  = (\Mux36~4_combout  & ((Mux18))) # (!\Mux36~4_combout  & (Mux19))

	.dataa(Mux191),
	.datab(gnd),
	.datac(Mux181),
	.datad(Mux36),
	.cin(gnd),
	.combout(\ShiftRight0~91_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~91 .lut_mask = 16'hF0AA;
defparam \ShiftRight0~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N6
cycloneive_lcell_comb \ShiftRight0~135 (
// Equation(s):
// \ShiftRight0~135_combout  = (\Mux35~2_combout  & (((\ShiftRight0~90_combout )))) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & (\ShiftRight0~90_combout )) # (!\Mux35~3_combout  & ((\ShiftRight0~91_combout )))))

	.dataa(Mux35),
	.datab(Mux351),
	.datac(\ShiftRight0~90_combout ),
	.datad(\ShiftRight0~91_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~135_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~135 .lut_mask = 16'hF1E0;
defparam \ShiftRight0~135 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N4
cycloneive_lcell_comb \ShiftRight0~93 (
// Equation(s):
// \ShiftRight0~93_combout  = (\Mux36~4_combout  & (Mux22)) # (!\Mux36~4_combout  & ((Mux23)))

	.dataa(gnd),
	.datab(Mux221),
	.datac(Mux36),
	.datad(Mux231),
	.cin(gnd),
	.combout(\ShiftRight0~93_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~93 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N4
cycloneive_lcell_comb \ShiftRight0~92 (
// Equation(s):
// \ShiftRight0~92_combout  = (\Mux36~4_combout  & (Mux20)) # (!\Mux36~4_combout  & ((Mux21)))

	.dataa(Mux36),
	.datab(gnd),
	.datac(Mux201),
	.datad(Mux211),
	.cin(gnd),
	.combout(\ShiftRight0~92_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~92 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N16
cycloneive_lcell_comb \ShiftRight0~136 (
// Equation(s):
// \ShiftRight0~136_combout  = (\Mux35~3_combout  & (((\ShiftRight0~92_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftRight0~92_combout ))) # (!\Mux35~2_combout  & (\ShiftRight0~93_combout ))))

	.dataa(Mux351),
	.datab(\ShiftRight0~93_combout ),
	.datac(\ShiftRight0~92_combout ),
	.datad(Mux35),
	.cin(gnd),
	.combout(\ShiftRight0~136_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~136 .lut_mask = 16'hF0E4;
defparam \ShiftRight0~136 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N2
cycloneive_lcell_comb \ShiftRight0~94 (
// Equation(s):
// \ShiftRight0~94_combout  = (\Mux34~3_combout  & (\ShiftRight0~135_combout )) # (!\Mux34~3_combout  & ((\ShiftRight0~136_combout )))

	.dataa(Mux34),
	.datab(gnd),
	.datac(\ShiftRight0~135_combout ),
	.datad(\ShiftRight0~136_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~94_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~94 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N26
cycloneive_lcell_comb \ShiftRight0~88 (
// Equation(s):
// \ShiftRight0~88_combout  = (\Mux36~4_combout  & ((Mux26))) # (!\Mux36~4_combout  & (Mux27))

	.dataa(gnd),
	.datab(Mux271),
	.datac(Mux261),
	.datad(Mux36),
	.cin(gnd),
	.combout(\ShiftRight0~88_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~88 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N28
cycloneive_lcell_comb \ShiftRight0~87 (
// Equation(s):
// \ShiftRight0~87_combout  = (\Mux36~4_combout  & ((Mux24))) # (!\Mux36~4_combout  & (Mux25))

	.dataa(Mux251),
	.datab(Mux36),
	.datac(gnd),
	.datad(Mux241),
	.cin(gnd),
	.combout(\ShiftRight0~87_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~87 .lut_mask = 16'hEE22;
defparam \ShiftRight0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N30
cycloneive_lcell_comb \ShiftRight0~134 (
// Equation(s):
// \ShiftRight0~134_combout  = (\Mux35~2_combout  & (((\ShiftRight0~87_combout )))) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & ((\ShiftRight0~87_combout ))) # (!\Mux35~3_combout  & (\ShiftRight0~88_combout ))))

	.dataa(Mux35),
	.datab(Mux351),
	.datac(\ShiftRight0~88_combout ),
	.datad(\ShiftRight0~87_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~134_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~134 .lut_mask = 16'hFE10;
defparam \ShiftRight0~134 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N20
cycloneive_lcell_comb \ShiftRight0~85 (
// Equation(s):
// \ShiftRight0~85_combout  = (\Mux36~4_combout  & (Mux28)) # (!\Mux36~4_combout  & ((Mux29)))

	.dataa(gnd),
	.datab(Mux281),
	.datac(Mux36),
	.datad(Mux291),
	.cin(gnd),
	.combout(\ShiftRight0~85_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~85 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N12
cycloneive_lcell_comb \ShiftRight0~84 (
// Equation(s):
// \ShiftRight0~84_combout  = (!\Mux35~4_combout  & ((\Mux36~4_combout  & ((Mux30))) # (!\Mux36~4_combout  & (Mux31))))

	.dataa(Mux36),
	.datab(Mux311),
	.datac(Mux301),
	.datad(Mux352),
	.cin(gnd),
	.combout(\ShiftRight0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~84 .lut_mask = 16'h00E4;
defparam \ShiftRight0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N26
cycloneive_lcell_comb \ShiftRight0~86 (
// Equation(s):
// \ShiftRight0~86_combout  = (!\Mux34~3_combout  & ((\ShiftRight0~84_combout ) # ((\Mux35~4_combout  & \ShiftRight0~85_combout ))))

	.dataa(Mux34),
	.datab(Mux352),
	.datac(\ShiftRight0~85_combout ),
	.datad(\ShiftRight0~84_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~86 .lut_mask = 16'h5540;
defparam \ShiftRight0~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N24
cycloneive_lcell_comb \ShiftRight0~89 (
// Equation(s):
// \ShiftRight0~89_combout  = (!\Mux33~3_combout  & ((\ShiftRight0~86_combout ) # ((\Mux34~3_combout  & \ShiftRight0~134_combout ))))

	.dataa(Mux34),
	.datab(Mux33),
	.datac(\ShiftRight0~134_combout ),
	.datad(\ShiftRight0~86_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~89_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~89 .lut_mask = 16'h3320;
defparam \ShiftRight0~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N28
cycloneive_lcell_comb \ShiftRight0~95 (
// Equation(s):
// \ShiftRight0~95_combout  = (!\Mux32~4_combout  & ((\ShiftRight0~89_combout ) # ((\ShiftRight0~94_combout  & \Mux33~3_combout ))))

	.dataa(Mux32),
	.datab(\ShiftRight0~94_combout ),
	.datac(Mux33),
	.datad(\ShiftRight0~89_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~95_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~95 .lut_mask = 16'h5540;
defparam \ShiftRight0~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N12
cycloneive_lcell_comb \ShiftRight0~102 (
// Equation(s):
// \ShiftRight0~102_combout  = (\Mux36~4_combout  & (Mux10)) # (!\Mux36~4_combout  & ((Mux11)))

	.dataa(Mux101),
	.datab(gnd),
	.datac(Mux36),
	.datad(Mux111),
	.cin(gnd),
	.combout(\ShiftRight0~102_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~102 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N28
cycloneive_lcell_comb \ShiftRight0~101 (
// Equation(s):
// \ShiftRight0~101_combout  = (\Mux36~4_combout  & (Mux8)) # (!\Mux36~4_combout  & ((Mux9)))

	.dataa(gnd),
	.datab(Mux81),
	.datac(Mux36),
	.datad(Mux91),
	.cin(gnd),
	.combout(\ShiftRight0~101_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~101 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N22
cycloneive_lcell_comb \ShiftRight0~139 (
// Equation(s):
// \ShiftRight0~139_combout  = (\Mux35~3_combout  & (((\ShiftRight0~101_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftRight0~101_combout ))) # (!\Mux35~2_combout  & (\ShiftRight0~102_combout ))))

	.dataa(Mux351),
	.datab(Mux35),
	.datac(\ShiftRight0~102_combout ),
	.datad(\ShiftRight0~101_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~139_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~139 .lut_mask = 16'hFE10;
defparam \ShiftRight0~139 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N18
cycloneive_lcell_comb \ShiftRight0~104 (
// Equation(s):
// \ShiftRight0~104_combout  = (\Mux36~4_combout  & ((Mux14))) # (!\Mux36~4_combout  & (Mux15))

	.dataa(gnd),
	.datab(Mux152),
	.datac(Mux36),
	.datad(Mux141),
	.cin(gnd),
	.combout(\ShiftRight0~104_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~104 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N12
cycloneive_lcell_comb \ShiftRight0~140 (
// Equation(s):
// \ShiftRight0~140_combout  = (\Mux35~2_combout  & (\ShiftRight0~103_combout )) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & (\ShiftRight0~103_combout )) # (!\Mux35~3_combout  & ((\ShiftRight0~104_combout )))))

	.dataa(\ShiftRight0~103_combout ),
	.datab(Mux35),
	.datac(Mux351),
	.datad(\ShiftRight0~104_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~140_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~140 .lut_mask = 16'hABA8;
defparam \ShiftRight0~140 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N18
cycloneive_lcell_comb \Selector23~0 (
// Equation(s):
// \Selector23~0_combout  = (\Mux34~3_combout  & (\ShiftRight0~139_combout )) # (!\Mux34~3_combout  & ((\ShiftRight0~140_combout )))

	.dataa(Mux34),
	.datab(\ShiftRight0~139_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~140_combout ),
	.cin(gnd),
	.combout(\Selector23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~0 .lut_mask = 16'hDD88;
defparam \Selector23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N8
cycloneive_lcell_comb \ShiftRight0~105 (
// Equation(s):
// \ShiftRight0~105_combout  = (\Mux33~3_combout  & ((ShiftRight0))) # (!\Mux33~3_combout  & (\Selector23~0_combout ))

	.dataa(gnd),
	.datab(\Selector23~0_combout ),
	.datac(Mux33),
	.datad(ShiftRight0),
	.cin(gnd),
	.combout(\ShiftRight0~105_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~105 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N14
cycloneive_lcell_comb \Selector31~0 (
// Equation(s):
// \Selector31~0_combout  = (\Selector24~0_combout  & ((\ShiftRight0~95_combout ) # ((\Mux32~4_combout  & \ShiftRight0~105_combout ))))

	.dataa(Mux32),
	.datab(\ShiftRight0~95_combout ),
	.datac(\ShiftRight0~105_combout ),
	.datad(\Selector24~0_combout ),
	.cin(gnd),
	.combout(\Selector31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~0 .lut_mask = 16'hEC00;
defparam \Selector31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N22
cycloneive_lcell_comb \Selector0~13 (
// Equation(s):
// \Selector0~13_combout  = (!cuifaluOp_0 & (!cuifaluOp_31 & (cuifaluOp_1 & cuifaluOp_2)))

	.dataa(cuifaluOp_0),
	.datab(cuifaluOp_3),
	.datac(cuifaluOp_1),
	.datad(cuifaluOp_2),
	.cin(gnd),
	.combout(\Selector0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~13 .lut_mask = 16'h1000;
defparam \Selector0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N24
cycloneive_lcell_comb \Selector31~1 (
// Equation(s):
// \Selector31~1_combout  = (\Add0~0_combout  & ((\Selector0~10_combout ) # (\Selector0~13_combout )))

	.dataa(gnd),
	.datab(\Selector0~10_combout ),
	.datac(\Selector0~13_combout ),
	.datad(\Add0~0_combout ),
	.cin(gnd),
	.combout(\Selector31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~1 .lut_mask = 16'hFC00;
defparam \Selector31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N0
cycloneive_lcell_comb \LessThan1~1 (
// Equation(s):
// \LessThan1~1_cout  = CARRY((\Mux36~4_combout  & !Mux31))

	.dataa(Mux36),
	.datab(Mux311),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan1~1_cout ));
// synopsys translate_off
defparam \LessThan1~1 .lut_mask = 16'h0022;
defparam \LessThan1~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N2
cycloneive_lcell_comb \LessThan1~3 (
// Equation(s):
// \LessThan1~3_cout  = CARRY((Mux30 & ((!\LessThan1~1_cout ) # (!\Mux35~4_combout ))) # (!Mux30 & (!\Mux35~4_combout  & !\LessThan1~1_cout )))

	.dataa(Mux301),
	.datab(Mux352),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~1_cout ),
	.combout(),
	.cout(\LessThan1~3_cout ));
// synopsys translate_off
defparam \LessThan1~3 .lut_mask = 16'h002B;
defparam \LessThan1~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N4
cycloneive_lcell_comb \LessThan1~5 (
// Equation(s):
// \LessThan1~5_cout  = CARRY((\Mux34~3_combout  & ((!\LessThan1~3_cout ) # (!Mux29))) # (!\Mux34~3_combout  & (!Mux29 & !\LessThan1~3_cout )))

	.dataa(Mux34),
	.datab(Mux291),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~3_cout ),
	.combout(),
	.cout(\LessThan1~5_cout ));
// synopsys translate_off
defparam \LessThan1~5 .lut_mask = 16'h002B;
defparam \LessThan1~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N6
cycloneive_lcell_comb \LessThan1~7 (
// Equation(s):
// \LessThan1~7_cout  = CARRY((\Mux33~3_combout  & (Mux28 & !\LessThan1~5_cout )) # (!\Mux33~3_combout  & ((Mux28) # (!\LessThan1~5_cout ))))

	.dataa(Mux33),
	.datab(Mux281),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~5_cout ),
	.combout(),
	.cout(\LessThan1~7_cout ));
// synopsys translate_off
defparam \LessThan1~7 .lut_mask = 16'h004D;
defparam \LessThan1~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N8
cycloneive_lcell_comb \LessThan1~9 (
// Equation(s):
// \LessThan1~9_cout  = CARRY((\Mux32~4_combout  & ((!\LessThan1~7_cout ) # (!Mux27))) # (!\Mux32~4_combout  & (!Mux27 & !\LessThan1~7_cout )))

	.dataa(Mux32),
	.datab(Mux271),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~7_cout ),
	.combout(),
	.cout(\LessThan1~9_cout ));
// synopsys translate_off
defparam \LessThan1~9 .lut_mask = 16'h002B;
defparam \LessThan1~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N10
cycloneive_lcell_comb \LessThan1~11 (
// Equation(s):
// \LessThan1~11_cout  = CARRY((\Mux31~1_combout  & (Mux26 & !\LessThan1~9_cout )) # (!\Mux31~1_combout  & ((Mux26) # (!\LessThan1~9_cout ))))

	.dataa(Mux31),
	.datab(Mux261),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~9_cout ),
	.combout(),
	.cout(\LessThan1~11_cout ));
// synopsys translate_off
defparam \LessThan1~11 .lut_mask = 16'h004D;
defparam \LessThan1~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N12
cycloneive_lcell_comb \LessThan1~13 (
// Equation(s):
// \LessThan1~13_cout  = CARRY((\Mux30~1_combout  & ((!\LessThan1~11_cout ) # (!Mux25))) # (!\Mux30~1_combout  & (!Mux25 & !\LessThan1~11_cout )))

	.dataa(Mux30),
	.datab(Mux251),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~11_cout ),
	.combout(),
	.cout(\LessThan1~13_cout ));
// synopsys translate_off
defparam \LessThan1~13 .lut_mask = 16'h002B;
defparam \LessThan1~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N14
cycloneive_lcell_comb \LessThan1~15 (
// Equation(s):
// \LessThan1~15_cout  = CARRY((\Mux29~1_combout  & (Mux24 & !\LessThan1~13_cout )) # (!\Mux29~1_combout  & ((Mux24) # (!\LessThan1~13_cout ))))

	.dataa(Mux29),
	.datab(Mux241),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~13_cout ),
	.combout(),
	.cout(\LessThan1~15_cout ));
// synopsys translate_off
defparam \LessThan1~15 .lut_mask = 16'h004D;
defparam \LessThan1~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N16
cycloneive_lcell_comb \LessThan1~17 (
// Equation(s):
// \LessThan1~17_cout  = CARRY((Mux23 & (\Mux28~1_combout  & !\LessThan1~15_cout )) # (!Mux23 & ((\Mux28~1_combout ) # (!\LessThan1~15_cout ))))

	.dataa(Mux231),
	.datab(Mux28),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~15_cout ),
	.combout(),
	.cout(\LessThan1~17_cout ));
// synopsys translate_off
defparam \LessThan1~17 .lut_mask = 16'h004D;
defparam \LessThan1~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N18
cycloneive_lcell_comb \LessThan1~19 (
// Equation(s):
// \LessThan1~19_cout  = CARRY((Mux22 & ((!\LessThan1~17_cout ) # (!\Mux27~1_combout ))) # (!Mux22 & (!\Mux27~1_combout  & !\LessThan1~17_cout )))

	.dataa(Mux221),
	.datab(Mux27),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~17_cout ),
	.combout(),
	.cout(\LessThan1~19_cout ));
// synopsys translate_off
defparam \LessThan1~19 .lut_mask = 16'h002B;
defparam \LessThan1~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N20
cycloneive_lcell_comb \LessThan1~21 (
// Equation(s):
// \LessThan1~21_cout  = CARRY((Mux21 & (\Mux26~1_combout  & !\LessThan1~19_cout )) # (!Mux21 & ((\Mux26~1_combout ) # (!\LessThan1~19_cout ))))

	.dataa(Mux211),
	.datab(Mux26),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~19_cout ),
	.combout(),
	.cout(\LessThan1~21_cout ));
// synopsys translate_off
defparam \LessThan1~21 .lut_mask = 16'h004D;
defparam \LessThan1~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N22
cycloneive_lcell_comb \LessThan1~23 (
// Equation(s):
// \LessThan1~23_cout  = CARRY((\Mux25~1_combout  & (Mux20 & !\LessThan1~21_cout )) # (!\Mux25~1_combout  & ((Mux20) # (!\LessThan1~21_cout ))))

	.dataa(Mux25),
	.datab(Mux201),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~21_cout ),
	.combout(),
	.cout(\LessThan1~23_cout ));
// synopsys translate_off
defparam \LessThan1~23 .lut_mask = 16'h004D;
defparam \LessThan1~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N24
cycloneive_lcell_comb \LessThan1~25 (
// Equation(s):
// \LessThan1~25_cout  = CARRY((Mux19 & (\Mux24~1_combout  & !\LessThan1~23_cout )) # (!Mux19 & ((\Mux24~1_combout ) # (!\LessThan1~23_cout ))))

	.dataa(Mux191),
	.datab(Mux24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~23_cout ),
	.combout(),
	.cout(\LessThan1~25_cout ));
// synopsys translate_off
defparam \LessThan1~25 .lut_mask = 16'h004D;
defparam \LessThan1~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N26
cycloneive_lcell_comb \LessThan1~27 (
// Equation(s):
// \LessThan1~27_cout  = CARRY((Mux18 & ((!\LessThan1~25_cout ) # (!\Mux23~1_combout ))) # (!Mux18 & (!\Mux23~1_combout  & !\LessThan1~25_cout )))

	.dataa(Mux181),
	.datab(Mux23),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~25_cout ),
	.combout(),
	.cout(\LessThan1~27_cout ));
// synopsys translate_off
defparam \LessThan1~27 .lut_mask = 16'h002B;
defparam \LessThan1~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N28
cycloneive_lcell_comb \LessThan1~29 (
// Equation(s):
// \LessThan1~29_cout  = CARRY((\Mux22~1_combout  & ((!\LessThan1~27_cout ) # (!Mux17))) # (!\Mux22~1_combout  & (!Mux17 & !\LessThan1~27_cout )))

	.dataa(Mux22),
	.datab(Mux171),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~27_cout ),
	.combout(),
	.cout(\LessThan1~29_cout ));
// synopsys translate_off
defparam \LessThan1~29 .lut_mask = 16'h002B;
defparam \LessThan1~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y43_N30
cycloneive_lcell_comb \LessThan1~31 (
// Equation(s):
// \LessThan1~31_cout  = CARRY((Mux16 & ((!\LessThan1~29_cout ) # (!\Mux21~1_combout ))) # (!Mux16 & (!\Mux21~1_combout  & !\LessThan1~29_cout )))

	.dataa(Mux161),
	.datab(Mux21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~29_cout ),
	.combout(),
	.cout(\LessThan1~31_cout ));
// synopsys translate_off
defparam \LessThan1~31 .lut_mask = 16'h002B;
defparam \LessThan1~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N0
cycloneive_lcell_comb \LessThan1~33 (
// Equation(s):
// \LessThan1~33_cout  = CARRY((\Mux20~1_combout  & ((!\LessThan1~31_cout ) # (!Mux15))) # (!\Mux20~1_combout  & (!Mux15 & !\LessThan1~31_cout )))

	.dataa(Mux20),
	.datab(Mux152),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~31_cout ),
	.combout(),
	.cout(\LessThan1~33_cout ));
// synopsys translate_off
defparam \LessThan1~33 .lut_mask = 16'h002B;
defparam \LessThan1~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N2
cycloneive_lcell_comb \LessThan1~35 (
// Equation(s):
// \LessThan1~35_cout  = CARRY((Mux14 & ((!\LessThan1~33_cout ) # (!\Mux19~1_combout ))) # (!Mux14 & (!\Mux19~1_combout  & !\LessThan1~33_cout )))

	.dataa(Mux141),
	.datab(Mux192),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~33_cout ),
	.combout(),
	.cout(\LessThan1~35_cout ));
// synopsys translate_off
defparam \LessThan1~35 .lut_mask = 16'h002B;
defparam \LessThan1~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N4
cycloneive_lcell_comb \LessThan1~37 (
// Equation(s):
// \LessThan1~37_cout  = CARRY((\Mux18~1_combout  & ((!\LessThan1~35_cout ) # (!Mux13))) # (!\Mux18~1_combout  & (!Mux13 & !\LessThan1~35_cout )))

	.dataa(Mux182),
	.datab(Mux131),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~35_cout ),
	.combout(),
	.cout(\LessThan1~37_cout ));
// synopsys translate_off
defparam \LessThan1~37 .lut_mask = 16'h002B;
defparam \LessThan1~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N6
cycloneive_lcell_comb \LessThan1~39 (
// Equation(s):
// \LessThan1~39_cout  = CARRY((\Mux17~1_combout  & (Mux12 & !\LessThan1~37_cout )) # (!\Mux17~1_combout  & ((Mux12) # (!\LessThan1~37_cout ))))

	.dataa(Mux172),
	.datab(Mux121),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~37_cout ),
	.combout(),
	.cout(\LessThan1~39_cout ));
// synopsys translate_off
defparam \LessThan1~39 .lut_mask = 16'h004D;
defparam \LessThan1~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N8
cycloneive_lcell_comb \LessThan1~41 (
// Equation(s):
// \LessThan1~41_cout  = CARRY((Mux11 & (\Mux16~1_combout  & !\LessThan1~39_cout )) # (!Mux11 & ((\Mux16~1_combout ) # (!\LessThan1~39_cout ))))

	.dataa(Mux111),
	.datab(Mux16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~39_cout ),
	.combout(),
	.cout(\LessThan1~41_cout ));
// synopsys translate_off
defparam \LessThan1~41 .lut_mask = 16'h004D;
defparam \LessThan1~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N10
cycloneive_lcell_comb \LessThan1~43 (
// Equation(s):
// \LessThan1~43_cout  = CARRY((\Mux15~1_combout  & (Mux10 & !\LessThan1~41_cout )) # (!\Mux15~1_combout  & ((Mux10) # (!\LessThan1~41_cout ))))

	.dataa(Mux151),
	.datab(Mux101),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~41_cout ),
	.combout(),
	.cout(\LessThan1~43_cout ));
// synopsys translate_off
defparam \LessThan1~43 .lut_mask = 16'h004D;
defparam \LessThan1~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N12
cycloneive_lcell_comb \LessThan1~45 (
// Equation(s):
// \LessThan1~45_cout  = CARRY((Mux9 & (\Mux14~1_combout  & !\LessThan1~43_cout )) # (!Mux9 & ((\Mux14~1_combout ) # (!\LessThan1~43_cout ))))

	.dataa(Mux91),
	.datab(Mux14),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~43_cout ),
	.combout(),
	.cout(\LessThan1~45_cout ));
// synopsys translate_off
defparam \LessThan1~45 .lut_mask = 16'h004D;
defparam \LessThan1~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N14
cycloneive_lcell_comb \LessThan1~47 (
// Equation(s):
// \LessThan1~47_cout  = CARRY((\Mux13~1_combout  & (Mux8 & !\LessThan1~45_cout )) # (!\Mux13~1_combout  & ((Mux8) # (!\LessThan1~45_cout ))))

	.dataa(Mux132),
	.datab(Mux81),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~45_cout ),
	.combout(),
	.cout(\LessThan1~47_cout ));
// synopsys translate_off
defparam \LessThan1~47 .lut_mask = 16'h004D;
defparam \LessThan1~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N16
cycloneive_lcell_comb \LessThan1~49 (
// Equation(s):
// \LessThan1~49_cout  = CARRY((\Mux12~1_combout  & ((!\LessThan1~47_cout ) # (!Mux7))) # (!\Mux12~1_combout  & (!Mux7 & !\LessThan1~47_cout )))

	.dataa(Mux12),
	.datab(Mux71),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~47_cout ),
	.combout(),
	.cout(\LessThan1~49_cout ));
// synopsys translate_off
defparam \LessThan1~49 .lut_mask = 16'h002B;
defparam \LessThan1~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N18
cycloneive_lcell_comb \LessThan1~51 (
// Equation(s):
// \LessThan1~51_cout  = CARRY((Mux6 & ((!\LessThan1~49_cout ) # (!\Mux11~1_combout ))) # (!Mux6 & (!\Mux11~1_combout  & !\LessThan1~49_cout )))

	.dataa(Mux61),
	.datab(Mux112),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~49_cout ),
	.combout(),
	.cout(\LessThan1~51_cout ));
// synopsys translate_off
defparam \LessThan1~51 .lut_mask = 16'h002B;
defparam \LessThan1~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N20
cycloneive_lcell_comb \LessThan1~53 (
// Equation(s):
// \LessThan1~53_cout  = CARRY((Mux5 & (\Mux10~1_combout  & !\LessThan1~51_cout )) # (!Mux5 & ((\Mux10~1_combout ) # (!\LessThan1~51_cout ))))

	.dataa(Mux52),
	.datab(Mux102),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~51_cout ),
	.combout(),
	.cout(\LessThan1~53_cout ));
// synopsys translate_off
defparam \LessThan1~53 .lut_mask = 16'h004D;
defparam \LessThan1~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N22
cycloneive_lcell_comb \LessThan1~55 (
// Equation(s):
// \LessThan1~55_cout  = CARRY((\Mux9~1_combout  & (Mux4 & !\LessThan1~53_cout )) # (!\Mux9~1_combout  & ((Mux4) # (!\LessThan1~53_cout ))))

	.dataa(Mux92),
	.datab(Mux4),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~53_cout ),
	.combout(),
	.cout(\LessThan1~55_cout ));
// synopsys translate_off
defparam \LessThan1~55 .lut_mask = 16'h004D;
defparam \LessThan1~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N24
cycloneive_lcell_comb \LessThan1~57 (
// Equation(s):
// \LessThan1~57_cout  = CARRY((\Mux8~1_combout  & ((!\LessThan1~55_cout ) # (!Mux3))) # (!\Mux8~1_combout  & (!Mux3 & !\LessThan1~55_cout )))

	.dataa(Mux82),
	.datab(Mux3),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~55_cout ),
	.combout(),
	.cout(\LessThan1~57_cout ));
// synopsys translate_off
defparam \LessThan1~57 .lut_mask = 16'h002B;
defparam \LessThan1~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N26
cycloneive_lcell_comb \LessThan1~59 (
// Equation(s):
// \LessThan1~59_cout  = CARRY((Mux2 & ((!\LessThan1~57_cout ) # (!\Mux7~1_combout ))) # (!Mux2 & (!\Mux7~1_combout  & !\LessThan1~57_cout )))

	.dataa(Mux2),
	.datab(Mux7),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~57_cout ),
	.combout(),
	.cout(\LessThan1~59_cout ));
// synopsys translate_off
defparam \LessThan1~59 .lut_mask = 16'h002B;
defparam \LessThan1~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N28
cycloneive_lcell_comb \LessThan1~61 (
// Equation(s):
// \LessThan1~61_cout  = CARRY((Mux1 & (\Mux6~1_combout  & !\LessThan1~59_cout )) # (!Mux1 & ((\Mux6~1_combout ) # (!\LessThan1~59_cout ))))

	.dataa(Mux1),
	.datab(Mux62),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~59_cout ),
	.combout(),
	.cout(\LessThan1~61_cout ));
// synopsys translate_off
defparam \LessThan1~61 .lut_mask = 16'h004D;
defparam \LessThan1~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y42_N30
cycloneive_lcell_comb \LessThan1~62 (
// Equation(s):
// \LessThan1~62_combout  = (Mux0 & (\LessThan1~61_cout  & \Mux5~6_combout )) # (!Mux0 & ((\LessThan1~61_cout ) # (\Mux5~6_combout )))

	.dataa(gnd),
	.datab(Mux0),
	.datac(gnd),
	.datad(Mux53),
	.cin(\LessThan1~61_cout ),
	.combout(\LessThan1~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan1~62 .lut_mask = 16'hF330;
defparam \LessThan1~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N0
cycloneive_lcell_comb \LessThan0~1 (
// Equation(s):
// \LessThan0~1_cout  = CARRY((\Mux36~4_combout  & !Mux31))

	.dataa(Mux36),
	.datab(Mux311),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan0~1_cout ));
// synopsys translate_off
defparam \LessThan0~1 .lut_mask = 16'h0022;
defparam \LessThan0~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N2
cycloneive_lcell_comb \LessThan0~3 (
// Equation(s):
// \LessThan0~3_cout  = CARRY((Mux30 & ((!\LessThan0~1_cout ) # (!\Mux35~4_combout ))) # (!Mux30 & (!\Mux35~4_combout  & !\LessThan0~1_cout )))

	.dataa(Mux301),
	.datab(Mux352),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~1_cout ),
	.combout(),
	.cout(\LessThan0~3_cout ));
// synopsys translate_off
defparam \LessThan0~3 .lut_mask = 16'h002B;
defparam \LessThan0~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N4
cycloneive_lcell_comb \LessThan0~5 (
// Equation(s):
// \LessThan0~5_cout  = CARRY((\Mux34~3_combout  & ((!\LessThan0~3_cout ) # (!Mux29))) # (!\Mux34~3_combout  & (!Mux29 & !\LessThan0~3_cout )))

	.dataa(Mux34),
	.datab(Mux291),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~3_cout ),
	.combout(),
	.cout(\LessThan0~5_cout ));
// synopsys translate_off
defparam \LessThan0~5 .lut_mask = 16'h002B;
defparam \LessThan0~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N6
cycloneive_lcell_comb \LessThan0~7 (
// Equation(s):
// \LessThan0~7_cout  = CARRY((\Mux33~3_combout  & (Mux28 & !\LessThan0~5_cout )) # (!\Mux33~3_combout  & ((Mux28) # (!\LessThan0~5_cout ))))

	.dataa(Mux33),
	.datab(Mux281),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~5_cout ),
	.combout(),
	.cout(\LessThan0~7_cout ));
// synopsys translate_off
defparam \LessThan0~7 .lut_mask = 16'h004D;
defparam \LessThan0~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N8
cycloneive_lcell_comb \LessThan0~9 (
// Equation(s):
// \LessThan0~9_cout  = CARRY((Mux27 & (\Mux32~4_combout  & !\LessThan0~7_cout )) # (!Mux27 & ((\Mux32~4_combout ) # (!\LessThan0~7_cout ))))

	.dataa(Mux271),
	.datab(Mux32),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~7_cout ),
	.combout(),
	.cout(\LessThan0~9_cout ));
// synopsys translate_off
defparam \LessThan0~9 .lut_mask = 16'h004D;
defparam \LessThan0~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N10
cycloneive_lcell_comb \LessThan0~11 (
// Equation(s):
// \LessThan0~11_cout  = CARRY((\Mux31~1_combout  & (Mux26 & !\LessThan0~9_cout )) # (!\Mux31~1_combout  & ((Mux26) # (!\LessThan0~9_cout ))))

	.dataa(Mux31),
	.datab(Mux261),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~9_cout ),
	.combout(),
	.cout(\LessThan0~11_cout ));
// synopsys translate_off
defparam \LessThan0~11 .lut_mask = 16'h004D;
defparam \LessThan0~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N12
cycloneive_lcell_comb \LessThan0~13 (
// Equation(s):
// \LessThan0~13_cout  = CARRY((\Mux30~1_combout  & ((!\LessThan0~11_cout ) # (!Mux25))) # (!\Mux30~1_combout  & (!Mux25 & !\LessThan0~11_cout )))

	.dataa(Mux30),
	.datab(Mux251),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~11_cout ),
	.combout(),
	.cout(\LessThan0~13_cout ));
// synopsys translate_off
defparam \LessThan0~13 .lut_mask = 16'h002B;
defparam \LessThan0~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N14
cycloneive_lcell_comb \LessThan0~15 (
// Equation(s):
// \LessThan0~15_cout  = CARRY((Mux24 & ((!\LessThan0~13_cout ) # (!\Mux29~1_combout ))) # (!Mux24 & (!\Mux29~1_combout  & !\LessThan0~13_cout )))

	.dataa(Mux241),
	.datab(Mux29),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~13_cout ),
	.combout(),
	.cout(\LessThan0~15_cout ));
// synopsys translate_off
defparam \LessThan0~15 .lut_mask = 16'h002B;
defparam \LessThan0~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N16
cycloneive_lcell_comb \LessThan0~17 (
// Equation(s):
// \LessThan0~17_cout  = CARRY((Mux23 & (\Mux28~1_combout  & !\LessThan0~15_cout )) # (!Mux23 & ((\Mux28~1_combout ) # (!\LessThan0~15_cout ))))

	.dataa(Mux231),
	.datab(Mux28),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~15_cout ),
	.combout(),
	.cout(\LessThan0~17_cout ));
// synopsys translate_off
defparam \LessThan0~17 .lut_mask = 16'h004D;
defparam \LessThan0~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N18
cycloneive_lcell_comb \LessThan0~19 (
// Equation(s):
// \LessThan0~19_cout  = CARRY((Mux22 & ((!\LessThan0~17_cout ) # (!\Mux27~1_combout ))) # (!Mux22 & (!\Mux27~1_combout  & !\LessThan0~17_cout )))

	.dataa(Mux221),
	.datab(Mux27),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~17_cout ),
	.combout(),
	.cout(\LessThan0~19_cout ));
// synopsys translate_off
defparam \LessThan0~19 .lut_mask = 16'h002B;
defparam \LessThan0~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N20
cycloneive_lcell_comb \LessThan0~21 (
// Equation(s):
// \LessThan0~21_cout  = CARRY((\Mux26~1_combout  & ((!\LessThan0~19_cout ) # (!Mux21))) # (!\Mux26~1_combout  & (!Mux21 & !\LessThan0~19_cout )))

	.dataa(Mux26),
	.datab(Mux211),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~19_cout ),
	.combout(),
	.cout(\LessThan0~21_cout ));
// synopsys translate_off
defparam \LessThan0~21 .lut_mask = 16'h002B;
defparam \LessThan0~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N22
cycloneive_lcell_comb \LessThan0~23 (
// Equation(s):
// \LessThan0~23_cout  = CARRY((\Mux25~1_combout  & (Mux20 & !\LessThan0~21_cout )) # (!\Mux25~1_combout  & ((Mux20) # (!\LessThan0~21_cout ))))

	.dataa(Mux25),
	.datab(Mux201),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~21_cout ),
	.combout(),
	.cout(\LessThan0~23_cout ));
// synopsys translate_off
defparam \LessThan0~23 .lut_mask = 16'h004D;
defparam \LessThan0~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N24
cycloneive_lcell_comb \LessThan0~25 (
// Equation(s):
// \LessThan0~25_cout  = CARRY((Mux19 & (\Mux24~1_combout  & !\LessThan0~23_cout )) # (!Mux19 & ((\Mux24~1_combout ) # (!\LessThan0~23_cout ))))

	.dataa(Mux191),
	.datab(Mux24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~23_cout ),
	.combout(),
	.cout(\LessThan0~25_cout ));
// synopsys translate_off
defparam \LessThan0~25 .lut_mask = 16'h004D;
defparam \LessThan0~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N26
cycloneive_lcell_comb \LessThan0~27 (
// Equation(s):
// \LessThan0~27_cout  = CARRY((\Mux23~1_combout  & (Mux18 & !\LessThan0~25_cout )) # (!\Mux23~1_combout  & ((Mux18) # (!\LessThan0~25_cout ))))

	.dataa(Mux23),
	.datab(Mux181),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~25_cout ),
	.combout(),
	.cout(\LessThan0~27_cout ));
// synopsys translate_off
defparam \LessThan0~27 .lut_mask = 16'h004D;
defparam \LessThan0~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N28
cycloneive_lcell_comb \LessThan0~29 (
// Equation(s):
// \LessThan0~29_cout  = CARRY((Mux17 & (\Mux22~1_combout  & !\LessThan0~27_cout )) # (!Mux17 & ((\Mux22~1_combout ) # (!\LessThan0~27_cout ))))

	.dataa(Mux171),
	.datab(Mux22),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~27_cout ),
	.combout(),
	.cout(\LessThan0~29_cout ));
// synopsys translate_off
defparam \LessThan0~29 .lut_mask = 16'h004D;
defparam \LessThan0~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y40_N30
cycloneive_lcell_comb \LessThan0~31 (
// Equation(s):
// \LessThan0~31_cout  = CARRY((Mux16 & ((!\LessThan0~29_cout ) # (!\Mux21~1_combout ))) # (!Mux16 & (!\Mux21~1_combout  & !\LessThan0~29_cout )))

	.dataa(Mux161),
	.datab(Mux21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~29_cout ),
	.combout(),
	.cout(\LessThan0~31_cout ));
// synopsys translate_off
defparam \LessThan0~31 .lut_mask = 16'h002B;
defparam \LessThan0~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N0
cycloneive_lcell_comb \LessThan0~33 (
// Equation(s):
// \LessThan0~33_cout  = CARRY((\Mux20~1_combout  & ((!\LessThan0~31_cout ) # (!Mux15))) # (!\Mux20~1_combout  & (!Mux15 & !\LessThan0~31_cout )))

	.dataa(Mux20),
	.datab(Mux152),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~31_cout ),
	.combout(),
	.cout(\LessThan0~33_cout ));
// synopsys translate_off
defparam \LessThan0~33 .lut_mask = 16'h002B;
defparam \LessThan0~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N2
cycloneive_lcell_comb \LessThan0~35 (
// Equation(s):
// \LessThan0~35_cout  = CARRY((\Mux19~1_combout  & (Mux14 & !\LessThan0~33_cout )) # (!\Mux19~1_combout  & ((Mux14) # (!\LessThan0~33_cout ))))

	.dataa(Mux192),
	.datab(Mux141),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~33_cout ),
	.combout(),
	.cout(\LessThan0~35_cout ));
// synopsys translate_off
defparam \LessThan0~35 .lut_mask = 16'h004D;
defparam \LessThan0~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N4
cycloneive_lcell_comb \LessThan0~37 (
// Equation(s):
// \LessThan0~37_cout  = CARRY((\Mux18~1_combout  & ((!\LessThan0~35_cout ) # (!Mux13))) # (!\Mux18~1_combout  & (!Mux13 & !\LessThan0~35_cout )))

	.dataa(Mux182),
	.datab(Mux131),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~35_cout ),
	.combout(),
	.cout(\LessThan0~37_cout ));
// synopsys translate_off
defparam \LessThan0~37 .lut_mask = 16'h002B;
defparam \LessThan0~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N6
cycloneive_lcell_comb \LessThan0~39 (
// Equation(s):
// \LessThan0~39_cout  = CARRY((Mux12 & ((!\LessThan0~37_cout ) # (!\Mux17~1_combout ))) # (!Mux12 & (!\Mux17~1_combout  & !\LessThan0~37_cout )))

	.dataa(Mux121),
	.datab(Mux172),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~37_cout ),
	.combout(),
	.cout(\LessThan0~39_cout ));
// synopsys translate_off
defparam \LessThan0~39 .lut_mask = 16'h002B;
defparam \LessThan0~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N8
cycloneive_lcell_comb \LessThan0~41 (
// Equation(s):
// \LessThan0~41_cout  = CARRY((\Mux16~1_combout  & ((!\LessThan0~39_cout ) # (!Mux11))) # (!\Mux16~1_combout  & (!Mux11 & !\LessThan0~39_cout )))

	.dataa(Mux16),
	.datab(Mux111),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~39_cout ),
	.combout(),
	.cout(\LessThan0~41_cout ));
// synopsys translate_off
defparam \LessThan0~41 .lut_mask = 16'h002B;
defparam \LessThan0~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N10
cycloneive_lcell_comb \LessThan0~43 (
// Equation(s):
// \LessThan0~43_cout  = CARRY((\Mux15~1_combout  & (Mux10 & !\LessThan0~41_cout )) # (!\Mux15~1_combout  & ((Mux10) # (!\LessThan0~41_cout ))))

	.dataa(Mux151),
	.datab(Mux101),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~41_cout ),
	.combout(),
	.cout(\LessThan0~43_cout ));
// synopsys translate_off
defparam \LessThan0~43 .lut_mask = 16'h004D;
defparam \LessThan0~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N12
cycloneive_lcell_comb \LessThan0~45 (
// Equation(s):
// \LessThan0~45_cout  = CARRY((\Mux14~1_combout  & ((!\LessThan0~43_cout ) # (!Mux9))) # (!\Mux14~1_combout  & (!Mux9 & !\LessThan0~43_cout )))

	.dataa(Mux14),
	.datab(Mux91),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~43_cout ),
	.combout(),
	.cout(\LessThan0~45_cout ));
// synopsys translate_off
defparam \LessThan0~45 .lut_mask = 16'h002B;
defparam \LessThan0~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N14
cycloneive_lcell_comb \LessThan0~47 (
// Equation(s):
// \LessThan0~47_cout  = CARRY((Mux8 & ((!\LessThan0~45_cout ) # (!\Mux13~1_combout ))) # (!Mux8 & (!\Mux13~1_combout  & !\LessThan0~45_cout )))

	.dataa(Mux81),
	.datab(Mux132),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~45_cout ),
	.combout(),
	.cout(\LessThan0~47_cout ));
// synopsys translate_off
defparam \LessThan0~47 .lut_mask = 16'h002B;
defparam \LessThan0~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N16
cycloneive_lcell_comb \LessThan0~49 (
// Equation(s):
// \LessThan0~49_cout  = CARRY((Mux7 & (\Mux12~1_combout  & !\LessThan0~47_cout )) # (!Mux7 & ((\Mux12~1_combout ) # (!\LessThan0~47_cout ))))

	.dataa(Mux71),
	.datab(Mux12),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~47_cout ),
	.combout(),
	.cout(\LessThan0~49_cout ));
// synopsys translate_off
defparam \LessThan0~49 .lut_mask = 16'h004D;
defparam \LessThan0~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N18
cycloneive_lcell_comb \LessThan0~51 (
// Equation(s):
// \LessThan0~51_cout  = CARRY((Mux6 & ((!\LessThan0~49_cout ) # (!\Mux11~1_combout ))) # (!Mux6 & (!\Mux11~1_combout  & !\LessThan0~49_cout )))

	.dataa(Mux61),
	.datab(Mux112),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~49_cout ),
	.combout(),
	.cout(\LessThan0~51_cout ));
// synopsys translate_off
defparam \LessThan0~51 .lut_mask = 16'h002B;
defparam \LessThan0~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N20
cycloneive_lcell_comb \LessThan0~53 (
// Equation(s):
// \LessThan0~53_cout  = CARRY((\Mux10~1_combout  & ((!\LessThan0~51_cout ) # (!Mux5))) # (!\Mux10~1_combout  & (!Mux5 & !\LessThan0~51_cout )))

	.dataa(Mux102),
	.datab(Mux52),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~51_cout ),
	.combout(),
	.cout(\LessThan0~53_cout ));
// synopsys translate_off
defparam \LessThan0~53 .lut_mask = 16'h002B;
defparam \LessThan0~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N22
cycloneive_lcell_comb \LessThan0~55 (
// Equation(s):
// \LessThan0~55_cout  = CARRY((Mux4 & ((!\LessThan0~53_cout ) # (!\Mux9~1_combout ))) # (!Mux4 & (!\Mux9~1_combout  & !\LessThan0~53_cout )))

	.dataa(Mux4),
	.datab(Mux92),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~53_cout ),
	.combout(),
	.cout(\LessThan0~55_cout ));
// synopsys translate_off
defparam \LessThan0~55 .lut_mask = 16'h002B;
defparam \LessThan0~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N24
cycloneive_lcell_comb \LessThan0~57 (
// Equation(s):
// \LessThan0~57_cout  = CARRY((Mux3 & (\Mux8~1_combout  & !\LessThan0~55_cout )) # (!Mux3 & ((\Mux8~1_combout ) # (!\LessThan0~55_cout ))))

	.dataa(Mux3),
	.datab(Mux82),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~55_cout ),
	.combout(),
	.cout(\LessThan0~57_cout ));
// synopsys translate_off
defparam \LessThan0~57 .lut_mask = 16'h004D;
defparam \LessThan0~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N26
cycloneive_lcell_comb \LessThan0~59 (
// Equation(s):
// \LessThan0~59_cout  = CARRY((\Mux7~1_combout  & (Mux2 & !\LessThan0~57_cout )) # (!\Mux7~1_combout  & ((Mux2) # (!\LessThan0~57_cout ))))

	.dataa(Mux7),
	.datab(Mux2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~57_cout ),
	.combout(),
	.cout(\LessThan0~59_cout ));
// synopsys translate_off
defparam \LessThan0~59 .lut_mask = 16'h004D;
defparam \LessThan0~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N28
cycloneive_lcell_comb \LessThan0~61 (
// Equation(s):
// \LessThan0~61_cout  = CARRY((Mux1 & (\Mux6~1_combout  & !\LessThan0~59_cout )) # (!Mux1 & ((\Mux6~1_combout ) # (!\LessThan0~59_cout ))))

	.dataa(Mux1),
	.datab(Mux62),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~59_cout ),
	.combout(),
	.cout(\LessThan0~61_cout ));
// synopsys translate_off
defparam \LessThan0~61 .lut_mask = 16'h004D;
defparam \LessThan0~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y39_N30
cycloneive_lcell_comb \LessThan0~62 (
// Equation(s):
// \LessThan0~62_combout  = (\Mux5~6_combout  & (\LessThan0~61_cout  & Mux0)) # (!\Mux5~6_combout  & ((\LessThan0~61_cout ) # (Mux0)))

	.dataa(gnd),
	.datab(Mux53),
	.datac(gnd),
	.datad(Mux0),
	.cin(\LessThan0~61_cout ),
	.combout(\LessThan0~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan0~62 .lut_mask = 16'hF330;
defparam \LessThan0~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N12
cycloneive_lcell_comb \Selector31~3 (
// Equation(s):
// \Selector31~3_combout  = (cuifaluOp_2 & ((cuifaluOp_0 & (\LessThan1~62_combout )) # (!cuifaluOp_0 & ((\LessThan0~62_combout )))))

	.dataa(cuifaluOp_0),
	.datab(cuifaluOp_2),
	.datac(\LessThan1~62_combout ),
	.datad(\LessThan0~62_combout ),
	.cin(gnd),
	.combout(\Selector31~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~3 .lut_mask = 16'hC480;
defparam \Selector31~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N18
cycloneive_lcell_comb \Selector31~4 (
// Equation(s):
// \Selector31~4_combout  = (\Selector31~2_combout ) # ((cuifaluOp_31 & (cuifaluOp_1 & \Selector31~3_combout )))

	.dataa(\Selector31~2_combout ),
	.datab(cuifaluOp_3),
	.datac(cuifaluOp_1),
	.datad(\Selector31~3_combout ),
	.cin(gnd),
	.combout(\Selector31~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~4 .lut_mask = 16'hEAAA;
defparam \Selector31~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N20
cycloneive_lcell_comb \Selector31~5 (
// Equation(s):
// \Selector31~5_combout  = (\Selector31~1_combout ) # ((\Selector31~4_combout ) # ((\Selector0~12_combout  & \Add1~0_combout )))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector31~1_combout ),
	.datac(\Add1~0_combout ),
	.datad(\Selector31~4_combout ),
	.cin(gnd),
	.combout(\Selector31~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~5 .lut_mask = 16'hFFEC;
defparam \Selector31~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N8
cycloneive_lcell_comb \ShiftRight0~106 (
// Equation(s):
// \ShiftRight0~106_combout  = (\Mux34~3_combout ) # ((\Mux35~4_combout ) # ((\Mux36~4_combout ) # (\Mux33~3_combout )))

	.dataa(Mux34),
	.datab(Mux352),
	.datac(Mux36),
	.datad(Mux33),
	.cin(gnd),
	.combout(\ShiftRight0~106_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~106 .lut_mask = 16'hFFFE;
defparam \ShiftRight0~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N6
cycloneive_lcell_comb \Selector31~7 (
// Equation(s):
// \Selector31~7_combout  = (!\Mux32~4_combout  & (!\ShiftRight0~106_combout  & (!\ShiftRight0~61_combout  & \Selector0~7_combout )))

	.dataa(Mux32),
	.datab(\ShiftRight0~106_combout ),
	.datac(\ShiftRight0~61_combout ),
	.datad(\Selector0~7_combout ),
	.cin(gnd),
	.combout(\Selector31~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector31~7 .lut_mask = 16'h0100;
defparam \Selector31~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N6
cycloneive_lcell_comb \ShiftRight0~109 (
// Equation(s):
// \ShiftRight0~109_combout  = (\Mux35~4_combout  & ((\Mux36~4_combout  & (Mux1)) # (!\Mux36~4_combout  & ((Mux2)))))

	.dataa(Mux36),
	.datab(Mux1),
	.datac(Mux2),
	.datad(Mux352),
	.cin(gnd),
	.combout(\ShiftRight0~109_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~109 .lut_mask = 16'hD800;
defparam \ShiftRight0~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N14
cycloneive_lcell_comb \ShiftRight0~145 (
// Equation(s):
// \ShiftRight0~145_combout  = (\ShiftRight0~109_combout ) # ((!\Mux35~3_combout  & (\ShiftRight0~76_combout  & !\Mux35~2_combout )))

	.dataa(Mux351),
	.datab(\ShiftRight0~76_combout ),
	.datac(Mux35),
	.datad(\ShiftRight0~109_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~145_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~145 .lut_mask = 16'hFF04;
defparam \ShiftRight0~145 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N18
cycloneive_lcell_comb \ShiftRight0~144 (
// Equation(s):
// \ShiftRight0~144_combout  = (!\Mux35~3_combout  & (!\Mux36~4_combout  & (!\Mux35~2_combout  & Mux0)))

	.dataa(Mux351),
	.datab(Mux36),
	.datac(Mux35),
	.datad(Mux0),
	.cin(gnd),
	.combout(\ShiftRight0~144_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~144 .lut_mask = 16'h0100;
defparam \ShiftRight0~144 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N4
cycloneive_lcell_comb \ShiftRight0~110 (
// Equation(s):
// \ShiftRight0~110_combout  = (\Mux34~3_combout  & ((\ShiftRight0~144_combout ))) # (!\Mux34~3_combout  & (\ShiftRight0~145_combout ))

	.dataa(Mux34),
	.datab(\ShiftRight0~145_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~144_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~110_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~110 .lut_mask = 16'hEE44;
defparam \ShiftRight0~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N24
cycloneive_lcell_comb \ShiftRight0~146 (
// Equation(s):
// \ShiftRight0~146_combout  = (\Mux35~3_combout  & (((\ShiftRight0~77_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftRight0~77_combout ))) # (!\Mux35~2_combout  & (\ShiftRight0~79_combout ))))

	.dataa(Mux351),
	.datab(Mux35),
	.datac(\ShiftRight0~79_combout ),
	.datad(\ShiftRight0~77_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~146_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~146 .lut_mask = 16'hFE10;
defparam \ShiftRight0~146 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N22
cycloneive_lcell_comb \ShiftRight0~81 (
// Equation(s):
// \ShiftRight0~81_combout  = (\Mux36~4_combout  & (Mux11)) # (!\Mux36~4_combout  & ((Mux12)))

	.dataa(Mux111),
	.datab(Mux121),
	.datac(Mux36),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~81 .lut_mask = 16'hACAC;
defparam \ShiftRight0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N10
cycloneive_lcell_comb \ShiftRight0~147 (
// Equation(s):
// \ShiftRight0~147_combout  = (\Mux35~3_combout  & (((\ShiftRight0~80_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftRight0~80_combout ))) # (!\Mux35~2_combout  & (\ShiftRight0~81_combout ))))

	.dataa(Mux351),
	.datab(Mux35),
	.datac(\ShiftRight0~81_combout ),
	.datad(\ShiftRight0~80_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~147_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~147 .lut_mask = 16'hFE10;
defparam \ShiftRight0~147 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N0
cycloneive_lcell_comb \Selector20~1 (
// Equation(s):
// \Selector20~1_combout  = (\Mux34~3_combout  & (\ShiftRight0~146_combout )) # (!\Mux34~3_combout  & ((\ShiftRight0~147_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~146_combout ),
	.datac(Mux34),
	.datad(\ShiftRight0~147_combout ),
	.cin(gnd),
	.combout(\Selector20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~1 .lut_mask = 16'hCFC0;
defparam \Selector20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N18
cycloneive_lcell_comb \ShiftRight0~111 (
// Equation(s):
// \ShiftRight0~111_combout  = (\Mux33~3_combout  & (\ShiftRight0~110_combout )) # (!\Mux33~3_combout  & ((\Selector20~1_combout )))

	.dataa(Mux33),
	.datab(gnd),
	.datac(\ShiftRight0~110_combout ),
	.datad(\Selector20~1_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~111_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~111 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~111 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N26
cycloneive_lcell_comb \ShiftLeft0~53 (
// Equation(s):
// \ShiftLeft0~53_combout  = (\Mux36~4_combout  & (Mux29)) # (!\Mux36~4_combout  & ((Mux28)))

	.dataa(gnd),
	.datab(Mux291),
	.datac(Mux36),
	.datad(Mux281),
	.cin(gnd),
	.combout(\ShiftLeft0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~53 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N2
cycloneive_lcell_comb \ShiftLeft0~106 (
// Equation(s):
// \ShiftLeft0~106_combout  = (\Mux35~3_combout  & (((\ShiftLeft0~52_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & (\ShiftLeft0~52_combout )) # (!\Mux35~2_combout  & ((\ShiftLeft0~53_combout )))))

	.dataa(Mux351),
	.datab(Mux35),
	.datac(\ShiftLeft0~52_combout ),
	.datad(\ShiftLeft0~53_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~106_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~106 .lut_mask = 16'hF1E0;
defparam \ShiftLeft0~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N30
cycloneive_lcell_comb \Selector0~14 (
// Equation(s):
// \Selector0~14_combout  = (!cuifaluOp_0 & (!cuifaluOp_1 & (!cuifaluOp_31 & cuifaluOp_2)))

	.dataa(cuifaluOp_0),
	.datab(cuifaluOp_1),
	.datac(cuifaluOp_3),
	.datad(cuifaluOp_2),
	.cin(gnd),
	.combout(\Selector0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~14 .lut_mask = 16'h0100;
defparam \Selector0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N4
cycloneive_lcell_comb \Selector16~0 (
// Equation(s):
// \Selector16~0_combout  = (!\Mux32~4_combout  & (\Selector0~14_combout  & !\ShiftRight0~61_combout ))

	.dataa(gnd),
	.datab(Mux32),
	.datac(\Selector0~14_combout ),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\Selector16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~0 .lut_mask = 16'h0030;
defparam \Selector16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N12
cycloneive_lcell_comb \Selector28~12 (
// Equation(s):
// \Selector28~12_combout  = (!\Mux34~3_combout  & (\ShiftLeft0~106_combout  & (\Selector16~0_combout  & !\Mux33~3_combout )))

	.dataa(Mux34),
	.datab(\ShiftLeft0~106_combout ),
	.datac(\Selector16~0_combout ),
	.datad(Mux33),
	.cin(gnd),
	.combout(\Selector28~12_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~12 .lut_mask = 16'h0040;
defparam \Selector28~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N24
cycloneive_lcell_comb \Selector0~21 (
// Equation(s):
// \Selector0~21_combout  = (!cuifaluOp_31 & (!cuifaluOp_1 & (cuifaluOp_2 & !\ShiftRight0~61_combout )))

	.dataa(cuifaluOp_3),
	.datab(cuifaluOp_1),
	.datac(cuifaluOp_2),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\Selector0~21_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~21 .lut_mask = 16'h0010;
defparam \Selector0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N30
cycloneive_lcell_comb \Selector20~0 (
// Equation(s):
// \Selector20~0_combout  = (cuifaluOp_0 & (\Mux32~4_combout  & \Selector0~21_combout ))

	.dataa(cuifaluOp_0),
	.datab(gnd),
	.datac(Mux32),
	.datad(\Selector0~21_combout ),
	.cin(gnd),
	.combout(\Selector20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~0 .lut_mask = 16'hA000;
defparam \Selector20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N22
cycloneive_lcell_comb \Selector2~2 (
// Equation(s):
// \Selector2~2_combout  = (cuifaluOp_31) # (((\Mux32~4_combout  & !\ShiftRight0~61_combout )) # (!cuifaluOp_2))

	.dataa(cuifaluOp_3),
	.datab(Mux32),
	.datac(cuifaluOp_2),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\Selector2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~2 .lut_mask = 16'hAFEF;
defparam \Selector2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N0
cycloneive_lcell_comb \Selector28~7 (
// Equation(s):
// \Selector28~7_combout  = (!cuifaluOp_1 & (cuifaluOp_0 & (!\Selector2~2_combout  & !\ShiftRight0~61_combout )))

	.dataa(cuifaluOp_1),
	.datab(cuifaluOp_0),
	.datac(\Selector2~2_combout ),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\Selector28~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~7 .lut_mask = 16'h0004;
defparam \Selector28~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N22
cycloneive_lcell_comb \Selector0~17 (
// Equation(s):
// \Selector0~17_combout  = (cuifaluOp_1 & (!cuifaluOp_31 & (!cuifaluOp_2 & !cuifaluOp_0)))

	.dataa(cuifaluOp_1),
	.datab(cuifaluOp_3),
	.datac(cuifaluOp_2),
	.datad(cuifaluOp_0),
	.cin(gnd),
	.combout(\Selector0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~17 .lut_mask = 16'h0002;
defparam \Selector0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N2
cycloneive_lcell_comb \Selector0~15 (
// Equation(s):
// \Selector0~15_combout  = (!cuifaluOp_1 & (!cuifaluOp_31 & (!cuifaluOp_2 & cuifaluOp_0)))

	.dataa(cuifaluOp_1),
	.datab(cuifaluOp_3),
	.datac(cuifaluOp_2),
	.datad(cuifaluOp_0),
	.cin(gnd),
	.combout(\Selector0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~15 .lut_mask = 16'h0100;
defparam \Selector0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N26
cycloneive_lcell_comb \Selector28~2 (
// Equation(s):
// \Selector28~2_combout  = (\Selector0~15_combout ) # ((\Selector0~16_combout  & Mux28))

	.dataa(\Selector0~16_combout ),
	.datab(gnd),
	.datac(Mux281),
	.datad(\Selector0~15_combout ),
	.cin(gnd),
	.combout(\Selector28~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~2 .lut_mask = 16'hFFA0;
defparam \Selector28~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N4
cycloneive_lcell_comb \Selector28~3 (
// Equation(s):
// \Selector28~3_combout  = (\Mux33~3_combout  & ((\Selector28~2_combout ) # ((\Selector0~17_combout  & !Mux28)))) # (!\Mux33~3_combout  & (\Selector0~17_combout  & ((Mux28))))

	.dataa(Mux33),
	.datab(\Selector0~17_combout ),
	.datac(\Selector28~2_combout ),
	.datad(Mux281),
	.cin(gnd),
	.combout(\Selector28~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~3 .lut_mask = 16'hE4A8;
defparam \Selector28~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N0
cycloneive_lcell_comb \ShiftRight0~107 (
// Equation(s):
// \ShiftRight0~107_combout  = (!\Mux34~3_combout  & !\Mux33~3_combout )

	.dataa(Mux34),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux33),
	.cin(gnd),
	.combout(\ShiftRight0~107_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~107 .lut_mask = 16'h0055;
defparam \ShiftRight0~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N18
cycloneive_lcell_comb \Selector2~14 (
// Equation(s):
// \Selector2~14_combout  = (\Mux33~3_combout ) # ((!\Mux34~3_combout  & ((\Mux35~3_combout ) # (\Mux35~2_combout ))))

	.dataa(Mux351),
	.datab(Mux35),
	.datac(Mux34),
	.datad(Mux33),
	.cin(gnd),
	.combout(\Selector2~14_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~14 .lut_mask = 16'hFF0E;
defparam \Selector2~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N8
cycloneive_lcell_comb \ShiftRight0~141 (
// Equation(s):
// \ShiftRight0~141_combout  = (\Mux35~3_combout  & (((\ShiftRight0~71_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & (\ShiftRight0~71_combout )) # (!\Mux35~2_combout  & ((\ShiftRight0~65_combout )))))

	.dataa(Mux351),
	.datab(Mux35),
	.datac(\ShiftRight0~71_combout ),
	.datad(\ShiftRight0~65_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~141_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~141 .lut_mask = 16'hF1E0;
defparam \ShiftRight0~141 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N20
cycloneive_lcell_comb \Selector28~8 (
// Equation(s):
// \Selector28~8_combout  = (\ShiftRight0~107_combout  & (\ShiftRight0~63_combout  & (!\Selector2~14_combout ))) # (!\ShiftRight0~107_combout  & (((\Selector2~14_combout ) # (\ShiftRight0~141_combout ))))

	.dataa(\ShiftRight0~63_combout ),
	.datab(\ShiftRight0~107_combout ),
	.datac(\Selector2~14_combout ),
	.datad(\ShiftRight0~141_combout ),
	.cin(gnd),
	.combout(\Selector28~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~8 .lut_mask = 16'h3B38;
defparam \Selector28~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N26
cycloneive_lcell_comb \ShiftRight0~142 (
// Equation(s):
// \ShiftRight0~142_combout  = (\Mux35~3_combout  & (((\ShiftRight0~82_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftRight0~82_combout ))) # (!\Mux35~2_combout  & (\ShiftRight0~68_combout ))))

	.dataa(Mux351),
	.datab(Mux35),
	.datac(\ShiftRight0~68_combout ),
	.datad(\ShiftRight0~82_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~142_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~142 .lut_mask = 16'hFE10;
defparam \ShiftRight0~142 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N20
cycloneive_lcell_comb \ShiftRight0~143 (
// Equation(s):
// \ShiftRight0~143_combout  = (\Mux35~2_combout  & (((\ShiftRight0~69_combout )))) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & ((\ShiftRight0~69_combout ))) # (!\Mux35~3_combout  & (\ShiftRight0~70_combout ))))

	.dataa(\ShiftRight0~70_combout ),
	.datab(Mux35),
	.datac(Mux351),
	.datad(\ShiftRight0~69_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~143_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~143 .lut_mask = 16'hFE02;
defparam \ShiftRight0~143 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N10
cycloneive_lcell_comb \ShiftRight0~108 (
// Equation(s):
// \ShiftRight0~108_combout  = (\Mux34~3_combout  & (\ShiftRight0~142_combout )) # (!\Mux34~3_combout  & ((\ShiftRight0~143_combout )))

	.dataa(Mux34),
	.datab(gnd),
	.datac(\ShiftRight0~142_combout ),
	.datad(\ShiftRight0~143_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~108_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~108 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N14
cycloneive_lcell_comb \Selector28~9 (
// Equation(s):
// \Selector28~9_combout  = (\Selector2~14_combout  & ((\Selector28~8_combout  & (\ShiftRight0~108_combout )) # (!\Selector28~8_combout  & ((\ShiftRight0~66_combout ))))) # (!\Selector2~14_combout  & (\Selector28~8_combout ))

	.dataa(\Selector2~14_combout ),
	.datab(\Selector28~8_combout ),
	.datac(\ShiftRight0~108_combout ),
	.datad(\ShiftRight0~66_combout ),
	.cin(gnd),
	.combout(\Selector28~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~9 .lut_mask = 16'hE6C4;
defparam \Selector28~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N18
cycloneive_lcell_comb \Selector0~18 (
// Equation(s):
// \Selector0~18_combout  = (cuifaluOp_0 & (!cuifaluOp_2 & (!cuifaluOp_31 & cuifaluOp_1)))

	.dataa(cuifaluOp_0),
	.datab(cuifaluOp_2),
	.datac(cuifaluOp_3),
	.datad(cuifaluOp_1),
	.cin(gnd),
	.combout(\Selector0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~18 .lut_mask = 16'h0200;
defparam \Selector0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N22
cycloneive_lcell_comb \Selector28~4 (
// Equation(s):
// \Selector28~4_combout  = (!\Mux33~3_combout  & (\Selector0~18_combout  & !Mux28))

	.dataa(Mux33),
	.datab(\Selector0~18_combout ),
	.datac(gnd),
	.datad(Mux281),
	.cin(gnd),
	.combout(\Selector28~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~4 .lut_mask = 16'h0044;
defparam \Selector28~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N0
cycloneive_lcell_comb \Selector0~20 (
// Equation(s):
// \Selector0~20_combout  = (!cuifaluOp_0 & (cuifaluOp_2 & (!cuifaluOp_31 & cuifaluOp_1)))

	.dataa(cuifaluOp_0),
	.datab(cuifaluOp_2),
	.datac(cuifaluOp_3),
	.datad(cuifaluOp_1),
	.cin(gnd),
	.combout(\Selector0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~20 .lut_mask = 16'h0400;
defparam \Selector0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N4
cycloneive_lcell_comb \Add0~4 (
// Equation(s):
// \Add0~4_combout  = ((Mux29 $ (\Mux34~3_combout  $ (!\Add0~3 )))) # (GND)
// \Add0~5  = CARRY((Mux29 & ((\Mux34~3_combout ) # (!\Add0~3 ))) # (!Mux29 & (\Mux34~3_combout  & !\Add0~3 )))

	.dataa(Mux291),
	.datab(Mux34),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
// synopsys translate_off
defparam \Add0~4 .lut_mask = 16'h698E;
defparam \Add0~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N6
cycloneive_lcell_comb \Add0~6 (
// Equation(s):
// \Add0~6_combout  = (\Mux33~3_combout  & ((Mux28 & (\Add0~5  & VCC)) # (!Mux28 & (!\Add0~5 )))) # (!\Mux33~3_combout  & ((Mux28 & (!\Add0~5 )) # (!Mux28 & ((\Add0~5 ) # (GND)))))
// \Add0~7  = CARRY((\Mux33~3_combout  & (!Mux28 & !\Add0~5 )) # (!\Mux33~3_combout  & ((!\Add0~5 ) # (!Mux28))))

	.dataa(Mux33),
	.datab(Mux281),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
// synopsys translate_off
defparam \Add0~6 .lut_mask = 16'h9617;
defparam \Add0~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N4
cycloneive_lcell_comb \Add1~4 (
// Equation(s):
// \Add1~4_combout  = ((\Mux34~3_combout  $ (Mux29 $ (\Add1~3 )))) # (GND)
// \Add1~5  = CARRY((\Mux34~3_combout  & (Mux29 & !\Add1~3 )) # (!\Mux34~3_combout  & ((Mux29) # (!\Add1~3 ))))

	.dataa(Mux34),
	.datab(Mux291),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'h964D;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N6
cycloneive_lcell_comb \Add1~6 (
// Equation(s):
// \Add1~6_combout  = (Mux28 & ((\Mux33~3_combout  & (!\Add1~5 )) # (!\Mux33~3_combout  & (\Add1~5  & VCC)))) # (!Mux28 & ((\Mux33~3_combout  & ((\Add1~5 ) # (GND))) # (!\Mux33~3_combout  & (!\Add1~5 ))))
// \Add1~7  = CARRY((Mux28 & (\Mux33~3_combout  & !\Add1~5 )) # (!Mux28 & ((\Mux33~3_combout ) # (!\Add1~5 ))))

	.dataa(Mux281),
	.datab(Mux33),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h694D;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N24
cycloneive_lcell_comb \Selector28~5 (
// Equation(s):
// \Selector28~5_combout  = (\Selector0~19_combout  & ((\Add1~6_combout ) # ((\Selector0~20_combout  & \Add0~6_combout )))) # (!\Selector0~19_combout  & (\Selector0~20_combout  & (\Add0~6_combout )))

	.dataa(\Selector0~19_combout ),
	.datab(\Selector0~20_combout ),
	.datac(\Add0~6_combout ),
	.datad(\Add1~6_combout ),
	.cin(gnd),
	.combout(\Selector28~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~5 .lut_mask = 16'hEAC0;
defparam \Selector28~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N6
cycloneive_lcell_comb \Selector28~6 (
// Equation(s):
// \Selector28~6_combout  = (\Selector28~4_combout ) # ((\Selector28~5_combout ) # ((\Selector0~15_combout  & Mux28)))

	.dataa(\Selector0~15_combout ),
	.datab(Mux281),
	.datac(\Selector28~4_combout ),
	.datad(\Selector28~5_combout ),
	.cin(gnd),
	.combout(\Selector28~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~6 .lut_mask = 16'hFFF8;
defparam \Selector28~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N12
cycloneive_lcell_comb \Selector28~10 (
// Equation(s):
// \Selector28~10_combout  = (\Selector28~3_combout ) # ((\Selector28~6_combout ) # ((\Selector28~7_combout  & \Selector28~9_combout )))

	.dataa(\Selector28~7_combout ),
	.datab(\Selector28~3_combout ),
	.datac(\Selector28~9_combout ),
	.datad(\Selector28~6_combout ),
	.cin(gnd),
	.combout(\Selector28~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector28~10 .lut_mask = 16'hFFEC;
defparam \Selector28~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N24
cycloneive_lcell_comb \ShiftLeft0~58 (
// Equation(s):
// \ShiftLeft0~58_combout  = (\Mux36~4_combout  & ((Mux27))) # (!\Mux36~4_combout  & (Mux26))

	.dataa(gnd),
	.datab(Mux261),
	.datac(Mux36),
	.datad(Mux271),
	.cin(gnd),
	.combout(\ShiftLeft0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~58 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N10
cycloneive_lcell_comb \ShiftLeft0~59 (
// Equation(s):
// \ShiftLeft0~59_combout  = (\Mux36~4_combout  & ((Mux25))) # (!\Mux36~4_combout  & (Mux24))

	.dataa(gnd),
	.datab(Mux36),
	.datac(Mux241),
	.datad(Mux251),
	.cin(gnd),
	.combout(\ShiftLeft0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~59 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N18
cycloneive_lcell_comb \ShiftLeft0~109 (
// Equation(s):
// \ShiftLeft0~109_combout  = (\Mux35~2_combout  & (\ShiftLeft0~58_combout )) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & (\ShiftLeft0~58_combout )) # (!\Mux35~3_combout  & ((\ShiftLeft0~59_combout )))))

	.dataa(Mux35),
	.datab(\ShiftLeft0~58_combout ),
	.datac(Mux351),
	.datad(\ShiftLeft0~59_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~109_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~109 .lut_mask = 16'hCDC8;
defparam \ShiftLeft0~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N2
cycloneive_lcell_comb \Selector0~23 (
// Equation(s):
// \Selector0~23_combout  = (\Mux5~6_combout  & (((\Selector0~15_combout )))) # (!\Mux5~6_combout  & (\Selector0~18_combout  & ((!Mux0))))

	.dataa(\Selector0~18_combout ),
	.datab(\Selector0~15_combout ),
	.datac(Mux53),
	.datad(Mux0),
	.cin(gnd),
	.combout(\Selector0~23_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~23 .lut_mask = 16'hC0CA;
defparam \Selector0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N4
cycloneive_lcell_comb \Selector0~16 (
// Equation(s):
// \Selector0~16_combout  = (!cuifaluOp_1 & (!cuifaluOp_31 & (!cuifaluOp_2 & !cuifaluOp_0)))

	.dataa(cuifaluOp_1),
	.datab(cuifaluOp_3),
	.datac(cuifaluOp_2),
	.datad(cuifaluOp_0),
	.cin(gnd),
	.combout(\Selector0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~16 .lut_mask = 16'h0001;
defparam \Selector0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N12
cycloneive_lcell_comb \Selector0~24 (
// Equation(s):
// \Selector0~24_combout  = (\Selector0~15_combout ) # ((\Selector0~16_combout  & ((\Mux5~4_combout ) # (\Mux5~1_combout ))))

	.dataa(Mux51),
	.datab(\Selector0~16_combout ),
	.datac(\Selector0~15_combout ),
	.datad(Mux5),
	.cin(gnd),
	.combout(\Selector0~24_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~24 .lut_mask = 16'hFCF8;
defparam \Selector0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N22
cycloneive_lcell_comb \Selector0~25 (
// Equation(s):
// \Selector0~25_combout  = (cuifaluOp_0 & (!cuifaluOp_1 & (!cuifaluOp_31 & cuifaluOp_2)))

	.dataa(cuifaluOp_0),
	.datab(cuifaluOp_1),
	.datac(cuifaluOp_3),
	.datad(cuifaluOp_2),
	.cin(gnd),
	.combout(\Selector0~25_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~25 .lut_mask = 16'h0200;
defparam \Selector0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N0
cycloneive_lcell_comb \Selector8~0 (
// Equation(s):
// \Selector8~0_combout  = (!\Mux32~4_combout  & (\Selector0~25_combout  & !\ShiftRight0~61_combout ))

	.dataa(gnd),
	.datab(Mux32),
	.datac(\Selector0~25_combout ),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~0 .lut_mask = 16'h0030;
defparam \Selector8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N18
cycloneive_lcell_comb \Selector0~26 (
// Equation(s):
// \Selector0~26_combout  = (Mux0 & ((\Selector0~24_combout ) # ((!\ShiftRight0~106_combout  & \Selector8~0_combout ))))

	.dataa(\ShiftRight0~106_combout ),
	.datab(Mux0),
	.datac(\Selector0~24_combout ),
	.datad(\Selector8~0_combout ),
	.cin(gnd),
	.combout(\Selector0~26_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~26 .lut_mask = 16'hC4C0;
defparam \Selector0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N28
cycloneive_lcell_comb \Selector0~22 (
// Equation(s):
// \Selector0~22_combout  = (\Selector0~17_combout  & (Mux0 $ (((\Mux5~1_combout ) # (\Mux5~4_combout )))))

	.dataa(Mux5),
	.datab(Mux51),
	.datac(\Selector0~17_combout ),
	.datad(Mux0),
	.cin(gnd),
	.combout(\Selector0~22_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~22 .lut_mask = 16'h10E0;
defparam \Selector0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N22
cycloneive_lcell_comb \ShiftLeft0~57 (
// Equation(s):
// \ShiftLeft0~57_combout  = (\Mux36~4_combout  & ((Mux9))) # (!\Mux36~4_combout  & (Mux8))

	.dataa(Mux81),
	.datab(gnd),
	.datac(Mux91),
	.datad(Mux36),
	.cin(gnd),
	.combout(\ShiftLeft0~57_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~57 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N30
cycloneive_lcell_comb \ShiftLeft0~56 (
// Equation(s):
// \ShiftLeft0~56_combout  = (\Mux36~4_combout  & ((Mux11))) # (!\Mux36~4_combout  & (Mux10))

	.dataa(gnd),
	.datab(Mux101),
	.datac(Mux111),
	.datad(Mux36),
	.cin(gnd),
	.combout(\ShiftLeft0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~56 .lut_mask = 16'hF0CC;
defparam \ShiftLeft0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N0
cycloneive_lcell_comb \ShiftLeft0~108 (
// Equation(s):
// \ShiftLeft0~108_combout  = (\Mux35~2_combout  & (((\ShiftLeft0~56_combout )))) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & ((\ShiftLeft0~56_combout ))) # (!\Mux35~3_combout  & (\ShiftLeft0~57_combout ))))

	.dataa(Mux35),
	.datab(Mux351),
	.datac(\ShiftLeft0~57_combout ),
	.datad(\ShiftLeft0~56_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~108_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~108 .lut_mask = 16'hFE10;
defparam \ShiftLeft0~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N0
cycloneive_lcell_comb \ShiftLeft0~55 (
// Equation(s):
// \ShiftLeft0~55_combout  = (\Mux36~4_combout  & (Mux13)) # (!\Mux36~4_combout  & ((Mux12)))

	.dataa(gnd),
	.datab(Mux131),
	.datac(Mux121),
	.datad(Mux36),
	.cin(gnd),
	.combout(\ShiftLeft0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~55 .lut_mask = 16'hCCF0;
defparam \ShiftLeft0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N20
cycloneive_lcell_comb \ShiftLeft0~54 (
// Equation(s):
// \ShiftLeft0~54_combout  = (\Mux36~4_combout  & (Mux15)) # (!\Mux36~4_combout  & ((Mux14)))

	.dataa(gnd),
	.datab(Mux152),
	.datac(Mux36),
	.datad(Mux141),
	.cin(gnd),
	.combout(\ShiftLeft0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~54 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N6
cycloneive_lcell_comb \ShiftLeft0~107 (
// Equation(s):
// \ShiftLeft0~107_combout  = (\Mux35~3_combout  & (((\ShiftLeft0~54_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftLeft0~54_combout ))) # (!\Mux35~2_combout  & (\ShiftLeft0~55_combout ))))

	.dataa(Mux351),
	.datab(\ShiftLeft0~55_combout ),
	.datac(\ShiftLeft0~54_combout ),
	.datad(Mux35),
	.cin(gnd),
	.combout(\ShiftLeft0~107_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~107 .lut_mask = 16'hF0E4;
defparam \ShiftLeft0~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N18
cycloneive_lcell_comb \Selector0~28 (
// Equation(s):
// \Selector0~28_combout  = (\Mux34~3_combout  & ((\ShiftLeft0~107_combout ))) # (!\Mux34~3_combout  & (\ShiftLeft0~108_combout ))

	.dataa(Mux34),
	.datab(gnd),
	.datac(\ShiftLeft0~108_combout ),
	.datad(\ShiftLeft0~107_combout ),
	.cin(gnd),
	.combout(\Selector0~28_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~28 .lut_mask = 16'hFA50;
defparam \Selector0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N20
cycloneive_lcell_comb \ShiftLeft0~68 (
// Equation(s):
// \ShiftLeft0~68_combout  = (\Mux36~4_combout  & ((Mux5))) # (!\Mux36~4_combout  & (Mux4))

	.dataa(Mux4),
	.datab(gnd),
	.datac(Mux52),
	.datad(Mux36),
	.cin(gnd),
	.combout(\ShiftLeft0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~68 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N22
cycloneive_lcell_comb \ShiftLeft0~67 (
// Equation(s):
// \ShiftLeft0~67_combout  = (\Mux36~4_combout  & ((Mux7))) # (!\Mux36~4_combout  & (Mux6))

	.dataa(Mux61),
	.datab(Mux36),
	.datac(gnd),
	.datad(Mux71),
	.cin(gnd),
	.combout(\ShiftLeft0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~67 .lut_mask = 16'hEE22;
defparam \ShiftLeft0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N18
cycloneive_lcell_comb \ShiftLeft0~112 (
// Equation(s):
// \ShiftLeft0~112_combout  = (\Mux35~2_combout  & (((\ShiftLeft0~67_combout )))) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & ((\ShiftLeft0~67_combout ))) # (!\Mux35~3_combout  & (\ShiftLeft0~68_combout ))))

	.dataa(Mux35),
	.datab(Mux351),
	.datac(\ShiftLeft0~68_combout ),
	.datad(\ShiftLeft0~67_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~112_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~112 .lut_mask = 16'hFE10;
defparam \ShiftLeft0~112 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N8
cycloneive_lcell_comb \Selector0~41 (
// Equation(s):
// \Selector0~41_combout  = (\Mux34~3_combout ) # ((!\Mux35~3_combout  & (\Mux36~4_combout  & !\Mux35~2_combout )))

	.dataa(Mux351),
	.datab(Mux34),
	.datac(Mux36),
	.datad(Mux35),
	.cin(gnd),
	.combout(\Selector0~41_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~41 .lut_mask = 16'hCCDC;
defparam \Selector0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N4
cycloneive_lcell_comb \Selector0~32 (
// Equation(s):
// \Selector0~32_combout  = (\Selector0~31_combout  & ((\ShiftLeft0~112_combout ) # ((!\Selector0~41_combout )))) # (!\Selector0~31_combout  & (((Mux1 & \Selector0~41_combout ))))

	.dataa(\Selector0~31_combout ),
	.datab(\ShiftLeft0~112_combout ),
	.datac(Mux1),
	.datad(\Selector0~41_combout ),
	.cin(gnd),
	.combout(\Selector0~32_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~32 .lut_mask = 16'hD8AA;
defparam \Selector0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N10
cycloneive_lcell_comb \Selector0~33 (
// Equation(s):
// \Selector0~33_combout  = (cuifaluOp_31) # ((!\ShiftRight0~61_combout  & ((\Mux32~4_combout ) # (\Mux33~3_combout ))))

	.dataa(Mux32),
	.datab(Mux33),
	.datac(cuifaluOp_3),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\Selector0~33_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~33 .lut_mask = 16'hF0FE;
defparam \Selector0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N0
cycloneive_lcell_comb \Selector16~1 (
// Equation(s):
// \Selector16~1_combout  = (!cuifaluOp_1 & (!\ShiftRight0~61_combout  & (cuifaluOp_2 & !\Selector0~33_combout )))

	.dataa(cuifaluOp_1),
	.datab(\ShiftRight0~61_combout ),
	.datac(cuifaluOp_2),
	.datad(\Selector0~33_combout ),
	.cin(gnd),
	.combout(\Selector16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~1 .lut_mask = 16'h0010;
defparam \Selector16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N14
cycloneive_lcell_comb \Selector0~34 (
// Equation(s):
// \Selector0~34_combout  = (!cuifaluOp_0 & (\Selector0~32_combout  & \Selector16~1_combout ))

	.dataa(cuifaluOp_0),
	.datab(\Selector0~32_combout ),
	.datac(\Selector16~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector0~34_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~34 .lut_mask = 16'h4040;
defparam \Selector0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N2
cycloneive_lcell_comb \ShiftLeft0~64 (
// Equation(s):
// \ShiftLeft0~64_combout  = (\Mux36~4_combout  & ((Mux17))) # (!\Mux36~4_combout  & (Mux16))

	.dataa(Mux161),
	.datab(gnd),
	.datac(Mux36),
	.datad(Mux171),
	.cin(gnd),
	.combout(\ShiftLeft0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~64 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N4
cycloneive_lcell_comb \ShiftLeft0~63 (
// Equation(s):
// \ShiftLeft0~63_combout  = (\Mux36~4_combout  & (Mux19)) # (!\Mux36~4_combout  & ((Mux18)))

	.dataa(gnd),
	.datab(Mux191),
	.datac(Mux36),
	.datad(Mux181),
	.cin(gnd),
	.combout(\ShiftLeft0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~63 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N24
cycloneive_lcell_comb \ShiftLeft0~111 (
// Equation(s):
// \ShiftLeft0~111_combout  = (\Mux35~2_combout  & (((\ShiftLeft0~63_combout )))) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & ((\ShiftLeft0~63_combout ))) # (!\Mux35~3_combout  & (\ShiftLeft0~64_combout ))))

	.dataa(Mux35),
	.datab(Mux351),
	.datac(\ShiftLeft0~64_combout ),
	.datad(\ShiftLeft0~63_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~111_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~111 .lut_mask = 16'hFE10;
defparam \ShiftLeft0~111 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N8
cycloneive_lcell_comb \Selector8~1 (
// Equation(s):
// \Selector8~1_combout  = (\Mux34~3_combout  & (\ShiftLeft0~110_combout )) # (!\Mux34~3_combout  & ((\ShiftLeft0~111_combout )))

	.dataa(\ShiftLeft0~110_combout ),
	.datab(gnd),
	.datac(Mux34),
	.datad(\ShiftLeft0~111_combout ),
	.cin(gnd),
	.combout(\Selector8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~1 .lut_mask = 16'hAFA0;
defparam \Selector8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N22
cycloneive_lcell_comb \ShiftLeft0~65 (
// Equation(s):
// \ShiftLeft0~65_combout  = (\Mux33~3_combout  & ((ShiftLeft0))) # (!\Mux33~3_combout  & (\Selector8~1_combout ))

	.dataa(gnd),
	.datab(Mux33),
	.datac(\Selector8~1_combout ),
	.datad(ShiftLeft0),
	.cin(gnd),
	.combout(\ShiftLeft0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~65 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N2
cycloneive_lcell_comb \Selector0~40 (
// Equation(s):
// \Selector0~40_combout  = (!cuifaluOp_0 & (\Mux32~4_combout  & (\ShiftLeft0~65_combout  & \Selector0~21_combout )))

	.dataa(cuifaluOp_0),
	.datab(Mux32),
	.datac(\ShiftLeft0~65_combout ),
	.datad(\Selector0~21_combout ),
	.cin(gnd),
	.combout(\Selector0~40_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~40 .lut_mask = 16'h4000;
defparam \Selector0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N28
cycloneive_lcell_comb \Selector0~35 (
// Equation(s):
// \Selector0~35_combout  = (\Selector0~34_combout ) # ((\Selector0~40_combout ) # ((\Selector0~27_combout  & \Selector0~28_combout )))

	.dataa(\Selector0~27_combout ),
	.datab(\Selector0~28_combout ),
	.datac(\Selector0~34_combout ),
	.datad(\Selector0~40_combout ),
	.cin(gnd),
	.combout(\Selector0~35_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~35 .lut_mask = 16'hFFF8;
defparam \Selector0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N10
cycloneive_lcell_comb \Selector0~36 (
// Equation(s):
// \Selector0~36_combout  = (\Selector0~23_combout ) # ((\Selector0~26_combout ) # ((\Selector0~22_combout ) # (\Selector0~35_combout )))

	.dataa(\Selector0~23_combout ),
	.datab(\Selector0~26_combout ),
	.datac(\Selector0~22_combout ),
	.datad(\Selector0~35_combout ),
	.cin(gnd),
	.combout(\Selector0~36_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~36 .lut_mask = 16'hFFFE;
defparam \Selector0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N20
cycloneive_lcell_comb \Selector0~19 (
// Equation(s):
// \Selector0~19_combout  = (!cuifaluOp_31 & (cuifaluOp_1 & (cuifaluOp_2 & cuifaluOp_0)))

	.dataa(cuifaluOp_3),
	.datab(cuifaluOp_1),
	.datac(cuifaluOp_2),
	.datad(cuifaluOp_0),
	.cin(gnd),
	.combout(\Selector0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~19 .lut_mask = 16'h4000;
defparam \Selector0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N8
cycloneive_lcell_comb \Add1~8 (
// Equation(s):
// \Add1~8_combout  = ((Mux27 $ (\Mux32~4_combout  $ (\Add1~7 )))) # (GND)
// \Add1~9  = CARRY((Mux27 & ((!\Add1~7 ) # (!\Mux32~4_combout ))) # (!Mux27 & (!\Mux32~4_combout  & !\Add1~7 )))

	.dataa(Mux271),
	.datab(Mux32),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'h962B;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N12
cycloneive_lcell_comb \Add1~12 (
// Equation(s):
// \Add1~12_combout  = ((\Mux30~1_combout  $ (Mux25 $ (\Add1~11 )))) # (GND)
// \Add1~13  = CARRY((\Mux30~1_combout  & (Mux25 & !\Add1~11 )) # (!\Mux30~1_combout  & ((Mux25) # (!\Add1~11 ))))

	.dataa(Mux30),
	.datab(Mux251),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout(\Add1~13 ));
// synopsys translate_off
defparam \Add1~12 .lut_mask = 16'h964D;
defparam \Add1~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N14
cycloneive_lcell_comb \Add1~14 (
// Equation(s):
// \Add1~14_combout  = (\Mux29~1_combout  & ((Mux24 & (!\Add1~13 )) # (!Mux24 & ((\Add1~13 ) # (GND))))) # (!\Mux29~1_combout  & ((Mux24 & (\Add1~13  & VCC)) # (!Mux24 & (!\Add1~13 ))))
// \Add1~15  = CARRY((\Mux29~1_combout  & ((!\Add1~13 ) # (!Mux24))) # (!\Mux29~1_combout  & (!Mux24 & !\Add1~13 )))

	.dataa(Mux29),
	.datab(Mux241),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~13 ),
	.combout(\Add1~14_combout ),
	.cout(\Add1~15 ));
// synopsys translate_off
defparam \Add1~14 .lut_mask = 16'h692B;
defparam \Add1~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N16
cycloneive_lcell_comb \Add1~16 (
// Equation(s):
// \Add1~16_combout  = ((Mux23 $ (\Mux28~1_combout  $ (\Add1~15 )))) # (GND)
// \Add1~17  = CARRY((Mux23 & ((!\Add1~15 ) # (!\Mux28~1_combout ))) # (!Mux23 & (!\Mux28~1_combout  & !\Add1~15 )))

	.dataa(Mux231),
	.datab(Mux28),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~15 ),
	.combout(\Add1~16_combout ),
	.cout(\Add1~17 ));
// synopsys translate_off
defparam \Add1~16 .lut_mask = 16'h962B;
defparam \Add1~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N18
cycloneive_lcell_comb \Add1~18 (
// Equation(s):
// \Add1~18_combout  = (\Mux27~1_combout  & ((Mux22 & (!\Add1~17 )) # (!Mux22 & ((\Add1~17 ) # (GND))))) # (!\Mux27~1_combout  & ((Mux22 & (\Add1~17  & VCC)) # (!Mux22 & (!\Add1~17 ))))
// \Add1~19  = CARRY((\Mux27~1_combout  & ((!\Add1~17 ) # (!Mux22))) # (!\Mux27~1_combout  & (!Mux22 & !\Add1~17 )))

	.dataa(Mux27),
	.datab(Mux221),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~17 ),
	.combout(\Add1~18_combout ),
	.cout(\Add1~19 ));
// synopsys translate_off
defparam \Add1~18 .lut_mask = 16'h692B;
defparam \Add1~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N22
cycloneive_lcell_comb \Add1~22 (
// Equation(s):
// \Add1~22_combout  = (Mux20 & ((\Mux25~1_combout  & (!\Add1~21 )) # (!\Mux25~1_combout  & (\Add1~21  & VCC)))) # (!Mux20 & ((\Mux25~1_combout  & ((\Add1~21 ) # (GND))) # (!\Mux25~1_combout  & (!\Add1~21 ))))
// \Add1~23  = CARRY((Mux20 & (\Mux25~1_combout  & !\Add1~21 )) # (!Mux20 & ((\Mux25~1_combout ) # (!\Add1~21 ))))

	.dataa(Mux201),
	.datab(Mux25),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~21 ),
	.combout(\Add1~22_combout ),
	.cout(\Add1~23 ));
// synopsys translate_off
defparam \Add1~22 .lut_mask = 16'h694D;
defparam \Add1~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N24
cycloneive_lcell_comb \Add1~24 (
// Equation(s):
// \Add1~24_combout  = ((Mux19 $ (\Mux24~1_combout  $ (\Add1~23 )))) # (GND)
// \Add1~25  = CARRY((Mux19 & ((!\Add1~23 ) # (!\Mux24~1_combout ))) # (!Mux19 & (!\Mux24~1_combout  & !\Add1~23 )))

	.dataa(Mux191),
	.datab(Mux24),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~23 ),
	.combout(\Add1~24_combout ),
	.cout(\Add1~25 ));
// synopsys translate_off
defparam \Add1~24 .lut_mask = 16'h962B;
defparam \Add1~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N26
cycloneive_lcell_comb \Add1~26 (
// Equation(s):
// \Add1~26_combout  = (Mux18 & ((\Mux23~1_combout  & (!\Add1~25 )) # (!\Mux23~1_combout  & (\Add1~25  & VCC)))) # (!Mux18 & ((\Mux23~1_combout  & ((\Add1~25 ) # (GND))) # (!\Mux23~1_combout  & (!\Add1~25 ))))
// \Add1~27  = CARRY((Mux18 & (\Mux23~1_combout  & !\Add1~25 )) # (!Mux18 & ((\Mux23~1_combout ) # (!\Add1~25 ))))

	.dataa(Mux181),
	.datab(Mux23),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~25 ),
	.combout(\Add1~26_combout ),
	.cout(\Add1~27 ));
// synopsys translate_off
defparam \Add1~26 .lut_mask = 16'h694D;
defparam \Add1~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N28
cycloneive_lcell_comb \Add1~28 (
// Equation(s):
// \Add1~28_combout  = ((Mux17 $ (\Mux22~1_combout  $ (\Add1~27 )))) # (GND)
// \Add1~29  = CARRY((Mux17 & ((!\Add1~27 ) # (!\Mux22~1_combout ))) # (!Mux17 & (!\Mux22~1_combout  & !\Add1~27 )))

	.dataa(Mux171),
	.datab(Mux22),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~27 ),
	.combout(\Add1~28_combout ),
	.cout(\Add1~29 ));
// synopsys translate_off
defparam \Add1~28 .lut_mask = 16'h962B;
defparam \Add1~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y39_N30
cycloneive_lcell_comb \Add1~30 (
// Equation(s):
// \Add1~30_combout  = (\Mux21~1_combout  & ((Mux16 & (!\Add1~29 )) # (!Mux16 & ((\Add1~29 ) # (GND))))) # (!\Mux21~1_combout  & ((Mux16 & (\Add1~29  & VCC)) # (!Mux16 & (!\Add1~29 ))))
// \Add1~31  = CARRY((\Mux21~1_combout  & ((!\Add1~29 ) # (!Mux16))) # (!\Mux21~1_combout  & (!Mux16 & !\Add1~29 )))

	.dataa(Mux21),
	.datab(Mux161),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~29 ),
	.combout(\Add1~30_combout ),
	.cout(\Add1~31 ));
// synopsys translate_off
defparam \Add1~30 .lut_mask = 16'h692B;
defparam \Add1~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N0
cycloneive_lcell_comb \Add1~32 (
// Equation(s):
// \Add1~32_combout  = ((Mux15 $ (\Mux20~1_combout  $ (\Add1~31 )))) # (GND)
// \Add1~33  = CARRY((Mux15 & ((!\Add1~31 ) # (!\Mux20~1_combout ))) # (!Mux15 & (!\Mux20~1_combout  & !\Add1~31 )))

	.dataa(Mux152),
	.datab(Mux20),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~31 ),
	.combout(\Add1~32_combout ),
	.cout(\Add1~33 ));
// synopsys translate_off
defparam \Add1~32 .lut_mask = 16'h962B;
defparam \Add1~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N6
cycloneive_lcell_comb \Add1~38 (
// Equation(s):
// \Add1~38_combout  = (Mux12 & ((\Mux17~1_combout  & (!\Add1~37 )) # (!\Mux17~1_combout  & (\Add1~37  & VCC)))) # (!Mux12 & ((\Mux17~1_combout  & ((\Add1~37 ) # (GND))) # (!\Mux17~1_combout  & (!\Add1~37 ))))
// \Add1~39  = CARRY((Mux12 & (\Mux17~1_combout  & !\Add1~37 )) # (!Mux12 & ((\Mux17~1_combout ) # (!\Add1~37 ))))

	.dataa(Mux121),
	.datab(Mux172),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~37 ),
	.combout(\Add1~38_combout ),
	.cout(\Add1~39 ));
// synopsys translate_off
defparam \Add1~38 .lut_mask = 16'h694D;
defparam \Add1~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N8
cycloneive_lcell_comb \Add1~40 (
// Equation(s):
// \Add1~40_combout  = ((\Mux16~1_combout  $ (Mux11 $ (\Add1~39 )))) # (GND)
// \Add1~41  = CARRY((\Mux16~1_combout  & (Mux11 & !\Add1~39 )) # (!\Mux16~1_combout  & ((Mux11) # (!\Add1~39 ))))

	.dataa(Mux16),
	.datab(Mux111),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~39 ),
	.combout(\Add1~40_combout ),
	.cout(\Add1~41 ));
// synopsys translate_off
defparam \Add1~40 .lut_mask = 16'h964D;
defparam \Add1~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N10
cycloneive_lcell_comb \Add1~42 (
// Equation(s):
// \Add1~42_combout  = (Mux10 & ((\Mux15~1_combout  & (!\Add1~41 )) # (!\Mux15~1_combout  & (\Add1~41  & VCC)))) # (!Mux10 & ((\Mux15~1_combout  & ((\Add1~41 ) # (GND))) # (!\Mux15~1_combout  & (!\Add1~41 ))))
// \Add1~43  = CARRY((Mux10 & (\Mux15~1_combout  & !\Add1~41 )) # (!Mux10 & ((\Mux15~1_combout ) # (!\Add1~41 ))))

	.dataa(Mux101),
	.datab(Mux151),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~41 ),
	.combout(\Add1~42_combout ),
	.cout(\Add1~43 ));
// synopsys translate_off
defparam \Add1~42 .lut_mask = 16'h694D;
defparam \Add1~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N12
cycloneive_lcell_comb \Add1~44 (
// Equation(s):
// \Add1~44_combout  = ((Mux9 $ (\Mux14~1_combout  $ (\Add1~43 )))) # (GND)
// \Add1~45  = CARRY((Mux9 & ((!\Add1~43 ) # (!\Mux14~1_combout ))) # (!Mux9 & (!\Mux14~1_combout  & !\Add1~43 )))

	.dataa(Mux91),
	.datab(Mux14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~43 ),
	.combout(\Add1~44_combout ),
	.cout(\Add1~45 ));
// synopsys translate_off
defparam \Add1~44 .lut_mask = 16'h962B;
defparam \Add1~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N14
cycloneive_lcell_comb \Add1~46 (
// Equation(s):
// \Add1~46_combout  = (\Mux13~1_combout  & ((Mux8 & (!\Add1~45 )) # (!Mux8 & ((\Add1~45 ) # (GND))))) # (!\Mux13~1_combout  & ((Mux8 & (\Add1~45  & VCC)) # (!Mux8 & (!\Add1~45 ))))
// \Add1~47  = CARRY((\Mux13~1_combout  & ((!\Add1~45 ) # (!Mux8))) # (!\Mux13~1_combout  & (!Mux8 & !\Add1~45 )))

	.dataa(Mux132),
	.datab(Mux81),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~45 ),
	.combout(\Add1~46_combout ),
	.cout(\Add1~47 ));
// synopsys translate_off
defparam \Add1~46 .lut_mask = 16'h692B;
defparam \Add1~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N16
cycloneive_lcell_comb \Add1~48 (
// Equation(s):
// \Add1~48_combout  = ((\Mux12~1_combout  $ (Mux7 $ (\Add1~47 )))) # (GND)
// \Add1~49  = CARRY((\Mux12~1_combout  & (Mux7 & !\Add1~47 )) # (!\Mux12~1_combout  & ((Mux7) # (!\Add1~47 ))))

	.dataa(Mux12),
	.datab(Mux71),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~47 ),
	.combout(\Add1~48_combout ),
	.cout(\Add1~49 ));
// synopsys translate_off
defparam \Add1~48 .lut_mask = 16'h964D;
defparam \Add1~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N18
cycloneive_lcell_comb \Add1~50 (
// Equation(s):
// \Add1~50_combout  = (\Mux11~1_combout  & ((Mux6 & (!\Add1~49 )) # (!Mux6 & ((\Add1~49 ) # (GND))))) # (!\Mux11~1_combout  & ((Mux6 & (\Add1~49  & VCC)) # (!Mux6 & (!\Add1~49 ))))
// \Add1~51  = CARRY((\Mux11~1_combout  & ((!\Add1~49 ) # (!Mux6))) # (!\Mux11~1_combout  & (!Mux6 & !\Add1~49 )))

	.dataa(Mux112),
	.datab(Mux61),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~49 ),
	.combout(\Add1~50_combout ),
	.cout(\Add1~51 ));
// synopsys translate_off
defparam \Add1~50 .lut_mask = 16'h692B;
defparam \Add1~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N20
cycloneive_lcell_comb \Add1~52 (
// Equation(s):
// \Add1~52_combout  = ((Mux5 $ (\Mux10~1_combout  $ (\Add1~51 )))) # (GND)
// \Add1~53  = CARRY((Mux5 & ((!\Add1~51 ) # (!\Mux10~1_combout ))) # (!Mux5 & (!\Mux10~1_combout  & !\Add1~51 )))

	.dataa(Mux52),
	.datab(Mux102),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~51 ),
	.combout(\Add1~52_combout ),
	.cout(\Add1~53 ));
// synopsys translate_off
defparam \Add1~52 .lut_mask = 16'h962B;
defparam \Add1~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N22
cycloneive_lcell_comb \Add1~54 (
// Equation(s):
// \Add1~54_combout  = (Mux4 & ((\Mux9~1_combout  & (!\Add1~53 )) # (!\Mux9~1_combout  & (\Add1~53  & VCC)))) # (!Mux4 & ((\Mux9~1_combout  & ((\Add1~53 ) # (GND))) # (!\Mux9~1_combout  & (!\Add1~53 ))))
// \Add1~55  = CARRY((Mux4 & (\Mux9~1_combout  & !\Add1~53 )) # (!Mux4 & ((\Mux9~1_combout ) # (!\Add1~53 ))))

	.dataa(Mux4),
	.datab(Mux92),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~53 ),
	.combout(\Add1~54_combout ),
	.cout(\Add1~55 ));
// synopsys translate_off
defparam \Add1~54 .lut_mask = 16'h694D;
defparam \Add1~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N24
cycloneive_lcell_comb \Add1~56 (
// Equation(s):
// \Add1~56_combout  = ((\Mux8~1_combout  $ (Mux3 $ (\Add1~55 )))) # (GND)
// \Add1~57  = CARRY((\Mux8~1_combout  & (Mux3 & !\Add1~55 )) # (!\Mux8~1_combout  & ((Mux3) # (!\Add1~55 ))))

	.dataa(Mux82),
	.datab(Mux3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~55 ),
	.combout(\Add1~56_combout ),
	.cout(\Add1~57 ));
// synopsys translate_off
defparam \Add1~56 .lut_mask = 16'h964D;
defparam \Add1~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N26
cycloneive_lcell_comb \Add1~58 (
// Equation(s):
// \Add1~58_combout  = (Mux2 & ((\Mux7~1_combout  & (!\Add1~57 )) # (!\Mux7~1_combout  & (\Add1~57  & VCC)))) # (!Mux2 & ((\Mux7~1_combout  & ((\Add1~57 ) # (GND))) # (!\Mux7~1_combout  & (!\Add1~57 ))))
// \Add1~59  = CARRY((Mux2 & (\Mux7~1_combout  & !\Add1~57 )) # (!Mux2 & ((\Mux7~1_combout ) # (!\Add1~57 ))))

	.dataa(Mux2),
	.datab(Mux7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~57 ),
	.combout(\Add1~58_combout ),
	.cout(\Add1~59 ));
// synopsys translate_off
defparam \Add1~58 .lut_mask = 16'h694D;
defparam \Add1~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N28
cycloneive_lcell_comb \Add1~60 (
// Equation(s):
// \Add1~60_combout  = ((\Mux6~1_combout  $ (Mux1 $ (\Add1~59 )))) # (GND)
// \Add1~61  = CARRY((\Mux6~1_combout  & (Mux1 & !\Add1~59 )) # (!\Mux6~1_combout  & ((Mux1) # (!\Add1~59 ))))

	.dataa(Mux62),
	.datab(Mux1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~59 ),
	.combout(\Add1~60_combout ),
	.cout(\Add1~61 ));
// synopsys translate_off
defparam \Add1~60 .lut_mask = 16'h964D;
defparam \Add1~60 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y38_N30
cycloneive_lcell_comb \Add1~62 (
// Equation(s):
// \Add1~62_combout  = Mux0 $ (\Add1~61  $ (!\Mux5~6_combout ))

	.dataa(Mux0),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux53),
	.cin(\Add1~61 ),
	.combout(\Add1~62_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~62 .lut_mask = 16'h5AA5;
defparam \Add1~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N16
cycloneive_lcell_comb \Selector0~37 (
// Equation(s):
// \Selector0~37_combout  = (\Selector0~19_combout  & \Add1~62_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Selector0~19_combout ),
	.datad(\Add1~62_combout ),
	.cin(gnd),
	.combout(\Selector0~37_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~37 .lut_mask = 16'hF000;
defparam \Selector0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N8
cycloneive_lcell_comb \Add0~8 (
// Equation(s):
// \Add0~8_combout  = ((\Mux32~4_combout  $ (Mux27 $ (!\Add0~7 )))) # (GND)
// \Add0~9  = CARRY((\Mux32~4_combout  & ((Mux27) # (!\Add0~7 ))) # (!\Mux32~4_combout  & (Mux27 & !\Add0~7 )))

	.dataa(Mux32),
	.datab(Mux271),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
// synopsys translate_off
defparam \Add0~8 .lut_mask = 16'h698E;
defparam \Add0~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N12
cycloneive_lcell_comb \Add0~12 (
// Equation(s):
// \Add0~12_combout  = ((Mux25 $ (\Mux30~1_combout  $ (!\Add0~11 )))) # (GND)
// \Add0~13  = CARRY((Mux25 & ((\Mux30~1_combout ) # (!\Add0~11 ))) # (!Mux25 & (\Mux30~1_combout  & !\Add0~11 )))

	.dataa(Mux251),
	.datab(Mux30),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
// synopsys translate_off
defparam \Add0~12 .lut_mask = 16'h698E;
defparam \Add0~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N16
cycloneive_lcell_comb \Add0~16 (
// Equation(s):
// \Add0~16_combout  = ((Mux23 $ (\Mux28~1_combout  $ (!\Add0~15 )))) # (GND)
// \Add0~17  = CARRY((Mux23 & ((\Mux28~1_combout ) # (!\Add0~15 ))) # (!Mux23 & (\Mux28~1_combout  & !\Add0~15 )))

	.dataa(Mux231),
	.datab(Mux28),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
// synopsys translate_off
defparam \Add0~16 .lut_mask = 16'h698E;
defparam \Add0~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N20
cycloneive_lcell_comb \Add0~20 (
// Equation(s):
// \Add0~20_combout  = ((\Mux26~1_combout  $ (Mux21 $ (!\Add0~19 )))) # (GND)
// \Add0~21  = CARRY((\Mux26~1_combout  & ((Mux21) # (!\Add0~19 ))) # (!\Mux26~1_combout  & (Mux21 & !\Add0~19 )))

	.dataa(Mux26),
	.datab(Mux211),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
// synopsys translate_off
defparam \Add0~20 .lut_mask = 16'h698E;
defparam \Add0~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N22
cycloneive_lcell_comb \Add0~22 (
// Equation(s):
// \Add0~22_combout  = (Mux20 & ((\Mux25~1_combout  & (\Add0~21  & VCC)) # (!\Mux25~1_combout  & (!\Add0~21 )))) # (!Mux20 & ((\Mux25~1_combout  & (!\Add0~21 )) # (!\Mux25~1_combout  & ((\Add0~21 ) # (GND)))))
// \Add0~23  = CARRY((Mux20 & (!\Mux25~1_combout  & !\Add0~21 )) # (!Mux20 & ((!\Add0~21 ) # (!\Mux25~1_combout ))))

	.dataa(Mux201),
	.datab(Mux25),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
// synopsys translate_off
defparam \Add0~22 .lut_mask = 16'h9617;
defparam \Add0~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N26
cycloneive_lcell_comb \Add0~26 (
// Equation(s):
// \Add0~26_combout  = (\Mux23~1_combout  & ((Mux18 & (\Add0~25  & VCC)) # (!Mux18 & (!\Add0~25 )))) # (!\Mux23~1_combout  & ((Mux18 & (!\Add0~25 )) # (!Mux18 & ((\Add0~25 ) # (GND)))))
// \Add0~27  = CARRY((\Mux23~1_combout  & (!Mux18 & !\Add0~25 )) # (!\Mux23~1_combout  & ((!\Add0~25 ) # (!Mux18))))

	.dataa(Mux23),
	.datab(Mux181),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout(\Add0~27 ));
// synopsys translate_off
defparam \Add0~26 .lut_mask = 16'h9617;
defparam \Add0~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N28
cycloneive_lcell_comb \Add0~28 (
// Equation(s):
// \Add0~28_combout  = ((Mux17 $ (\Mux22~1_combout  $ (!\Add0~27 )))) # (GND)
// \Add0~29  = CARRY((Mux17 & ((\Mux22~1_combout ) # (!\Add0~27 ))) # (!Mux17 & (\Mux22~1_combout  & !\Add0~27 )))

	.dataa(Mux171),
	.datab(Mux22),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~27 ),
	.combout(\Add0~28_combout ),
	.cout(\Add0~29 ));
// synopsys translate_off
defparam \Add0~28 .lut_mask = 16'h698E;
defparam \Add0~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y41_N30
cycloneive_lcell_comb \Add0~30 (
// Equation(s):
// \Add0~30_combout  = (\Mux21~1_combout  & ((Mux16 & (\Add0~29  & VCC)) # (!Mux16 & (!\Add0~29 )))) # (!\Mux21~1_combout  & ((Mux16 & (!\Add0~29 )) # (!Mux16 & ((\Add0~29 ) # (GND)))))
// \Add0~31  = CARRY((\Mux21~1_combout  & (!Mux16 & !\Add0~29 )) # (!\Mux21~1_combout  & ((!\Add0~29 ) # (!Mux16))))

	.dataa(Mux21),
	.datab(Mux161),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~29 ),
	.combout(\Add0~30_combout ),
	.cout(\Add0~31 ));
// synopsys translate_off
defparam \Add0~30 .lut_mask = 16'h9617;
defparam \Add0~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N2
cycloneive_lcell_comb \Add0~34 (
// Equation(s):
// \Add0~34_combout  = (\Mux19~1_combout  & ((Mux14 & (\Add0~33  & VCC)) # (!Mux14 & (!\Add0~33 )))) # (!\Mux19~1_combout  & ((Mux14 & (!\Add0~33 )) # (!Mux14 & ((\Add0~33 ) # (GND)))))
// \Add0~35  = CARRY((\Mux19~1_combout  & (!Mux14 & !\Add0~33 )) # (!\Mux19~1_combout  & ((!\Add0~33 ) # (!Mux14))))

	.dataa(Mux192),
	.datab(Mux141),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~33 ),
	.combout(\Add0~34_combout ),
	.cout(\Add0~35 ));
// synopsys translate_off
defparam \Add0~34 .lut_mask = 16'h9617;
defparam \Add0~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N4
cycloneive_lcell_comb \Add0~36 (
// Equation(s):
// \Add0~36_combout  = ((Mux13 $ (\Mux18~1_combout  $ (!\Add0~35 )))) # (GND)
// \Add0~37  = CARRY((Mux13 & ((\Mux18~1_combout ) # (!\Add0~35 ))) # (!Mux13 & (\Mux18~1_combout  & !\Add0~35 )))

	.dataa(Mux131),
	.datab(Mux182),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~35 ),
	.combout(\Add0~36_combout ),
	.cout(\Add0~37 ));
// synopsys translate_off
defparam \Add0~36 .lut_mask = 16'h698E;
defparam \Add0~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N6
cycloneive_lcell_comb \Add0~38 (
// Equation(s):
// \Add0~38_combout  = (Mux12 & ((\Mux17~1_combout  & (\Add0~37  & VCC)) # (!\Mux17~1_combout  & (!\Add0~37 )))) # (!Mux12 & ((\Mux17~1_combout  & (!\Add0~37 )) # (!\Mux17~1_combout  & ((\Add0~37 ) # (GND)))))
// \Add0~39  = CARRY((Mux12 & (!\Mux17~1_combout  & !\Add0~37 )) # (!Mux12 & ((!\Add0~37 ) # (!\Mux17~1_combout ))))

	.dataa(Mux121),
	.datab(Mux172),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~37 ),
	.combout(\Add0~38_combout ),
	.cout(\Add0~39 ));
// synopsys translate_off
defparam \Add0~38 .lut_mask = 16'h9617;
defparam \Add0~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N8
cycloneive_lcell_comb \Add0~40 (
// Equation(s):
// \Add0~40_combout  = ((Mux11 $ (\Mux16~1_combout  $ (!\Add0~39 )))) # (GND)
// \Add0~41  = CARRY((Mux11 & ((\Mux16~1_combout ) # (!\Add0~39 ))) # (!Mux11 & (\Mux16~1_combout  & !\Add0~39 )))

	.dataa(Mux111),
	.datab(Mux16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~39 ),
	.combout(\Add0~40_combout ),
	.cout(\Add0~41 ));
// synopsys translate_off
defparam \Add0~40 .lut_mask = 16'h698E;
defparam \Add0~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N10
cycloneive_lcell_comb \Add0~42 (
// Equation(s):
// \Add0~42_combout  = (\Mux15~1_combout  & ((Mux10 & (\Add0~41  & VCC)) # (!Mux10 & (!\Add0~41 )))) # (!\Mux15~1_combout  & ((Mux10 & (!\Add0~41 )) # (!Mux10 & ((\Add0~41 ) # (GND)))))
// \Add0~43  = CARRY((\Mux15~1_combout  & (!Mux10 & !\Add0~41 )) # (!\Mux15~1_combout  & ((!\Add0~41 ) # (!Mux10))))

	.dataa(Mux151),
	.datab(Mux101),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~41 ),
	.combout(\Add0~42_combout ),
	.cout(\Add0~43 ));
// synopsys translate_off
defparam \Add0~42 .lut_mask = 16'h9617;
defparam \Add0~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N14
cycloneive_lcell_comb \Add0~46 (
// Equation(s):
// \Add0~46_combout  = (\Mux13~1_combout  & ((Mux8 & (\Add0~45  & VCC)) # (!Mux8 & (!\Add0~45 )))) # (!\Mux13~1_combout  & ((Mux8 & (!\Add0~45 )) # (!Mux8 & ((\Add0~45 ) # (GND)))))
// \Add0~47  = CARRY((\Mux13~1_combout  & (!Mux8 & !\Add0~45 )) # (!\Mux13~1_combout  & ((!\Add0~45 ) # (!Mux8))))

	.dataa(Mux132),
	.datab(Mux81),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~45 ),
	.combout(\Add0~46_combout ),
	.cout(\Add0~47 ));
// synopsys translate_off
defparam \Add0~46 .lut_mask = 16'h9617;
defparam \Add0~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N16
cycloneive_lcell_comb \Add0~48 (
// Equation(s):
// \Add0~48_combout  = ((\Mux12~1_combout  $ (Mux7 $ (!\Add0~47 )))) # (GND)
// \Add0~49  = CARRY((\Mux12~1_combout  & ((Mux7) # (!\Add0~47 ))) # (!\Mux12~1_combout  & (Mux7 & !\Add0~47 )))

	.dataa(Mux12),
	.datab(Mux71),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~47 ),
	.combout(\Add0~48_combout ),
	.cout(\Add0~49 ));
// synopsys translate_off
defparam \Add0~48 .lut_mask = 16'h698E;
defparam \Add0~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N18
cycloneive_lcell_comb \Add0~50 (
// Equation(s):
// \Add0~50_combout  = (Mux6 & ((\Mux11~1_combout  & (\Add0~49  & VCC)) # (!\Mux11~1_combout  & (!\Add0~49 )))) # (!Mux6 & ((\Mux11~1_combout  & (!\Add0~49 )) # (!\Mux11~1_combout  & ((\Add0~49 ) # (GND)))))
// \Add0~51  = CARRY((Mux6 & (!\Mux11~1_combout  & !\Add0~49 )) # (!Mux6 & ((!\Add0~49 ) # (!\Mux11~1_combout ))))

	.dataa(Mux61),
	.datab(Mux112),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~49 ),
	.combout(\Add0~50_combout ),
	.cout(\Add0~51 ));
// synopsys translate_off
defparam \Add0~50 .lut_mask = 16'h9617;
defparam \Add0~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N20
cycloneive_lcell_comb \Add0~52 (
// Equation(s):
// \Add0~52_combout  = ((\Mux10~1_combout  $ (Mux5 $ (!\Add0~51 )))) # (GND)
// \Add0~53  = CARRY((\Mux10~1_combout  & ((Mux5) # (!\Add0~51 ))) # (!\Mux10~1_combout  & (Mux5 & !\Add0~51 )))

	.dataa(Mux102),
	.datab(Mux52),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~51 ),
	.combout(\Add0~52_combout ),
	.cout(\Add0~53 ));
// synopsys translate_off
defparam \Add0~52 .lut_mask = 16'h698E;
defparam \Add0~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N22
cycloneive_lcell_comb \Add0~54 (
// Equation(s):
// \Add0~54_combout  = (Mux4 & ((\Mux9~1_combout  & (\Add0~53  & VCC)) # (!\Mux9~1_combout  & (!\Add0~53 )))) # (!Mux4 & ((\Mux9~1_combout  & (!\Add0~53 )) # (!\Mux9~1_combout  & ((\Add0~53 ) # (GND)))))
// \Add0~55  = CARRY((Mux4 & (!\Mux9~1_combout  & !\Add0~53 )) # (!Mux4 & ((!\Add0~53 ) # (!\Mux9~1_combout ))))

	.dataa(Mux4),
	.datab(Mux92),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~53 ),
	.combout(\Add0~54_combout ),
	.cout(\Add0~55 ));
// synopsys translate_off
defparam \Add0~54 .lut_mask = 16'h9617;
defparam \Add0~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N24
cycloneive_lcell_comb \Add0~56 (
// Equation(s):
// \Add0~56_combout  = ((\Mux8~1_combout  $ (Mux3 $ (!\Add0~55 )))) # (GND)
// \Add0~57  = CARRY((\Mux8~1_combout  & ((Mux3) # (!\Add0~55 ))) # (!\Mux8~1_combout  & (Mux3 & !\Add0~55 )))

	.dataa(Mux82),
	.datab(Mux3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~55 ),
	.combout(\Add0~56_combout ),
	.cout(\Add0~57 ));
// synopsys translate_off
defparam \Add0~56 .lut_mask = 16'h698E;
defparam \Add0~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N26
cycloneive_lcell_comb \Add0~58 (
// Equation(s):
// \Add0~58_combout  = (\Mux7~1_combout  & ((Mux2 & (\Add0~57  & VCC)) # (!Mux2 & (!\Add0~57 )))) # (!\Mux7~1_combout  & ((Mux2 & (!\Add0~57 )) # (!Mux2 & ((\Add0~57 ) # (GND)))))
// \Add0~59  = CARRY((\Mux7~1_combout  & (!Mux2 & !\Add0~57 )) # (!\Mux7~1_combout  & ((!\Add0~57 ) # (!Mux2))))

	.dataa(Mux7),
	.datab(Mux2),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~57 ),
	.combout(\Add0~58_combout ),
	.cout(\Add0~59 ));
// synopsys translate_off
defparam \Add0~58 .lut_mask = 16'h9617;
defparam \Add0~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N28
cycloneive_lcell_comb \Add0~60 (
// Equation(s):
// \Add0~60_combout  = ((\Mux6~1_combout  $ (Mux1 $ (!\Add0~59 )))) # (GND)
// \Add0~61  = CARRY((\Mux6~1_combout  & ((Mux1) # (!\Add0~59 ))) # (!\Mux6~1_combout  & (Mux1 & !\Add0~59 )))

	.dataa(Mux62),
	.datab(Mux1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~59 ),
	.combout(\Add0~60_combout ),
	.cout(\Add0~61 ));
// synopsys translate_off
defparam \Add0~60 .lut_mask = 16'h698E;
defparam \Add0~60 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y40_N30
cycloneive_lcell_comb \Add0~62 (
// Equation(s):
// \Add0~62_combout  = Mux0 $ (\Add0~61  $ (\Mux5~6_combout ))

	.dataa(Mux0),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux53),
	.cin(\Add0~61 ),
	.combout(\Add0~62_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~62 .lut_mask = 16'hA55A;
defparam \Add0~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N12
cycloneive_lcell_comb \ShiftLeft0~113 (
// Equation(s):
// \ShiftLeft0~113_combout  = (\Mux35~3_combout  & (((\ShiftLeft0~53_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftLeft0~53_combout ))) # (!\Mux35~2_combout  & (\ShiftLeft0~58_combout ))))

	.dataa(Mux351),
	.datab(\ShiftLeft0~58_combout ),
	.datac(\ShiftLeft0~53_combout ),
	.datad(Mux35),
	.cin(gnd),
	.combout(\ShiftLeft0~113_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~113 .lut_mask = 16'hF0E4;
defparam \ShiftLeft0~113 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N10
cycloneive_lcell_comb \Selector2~12 (
// Equation(s):
// \Selector2~12_combout  = (!cuifaluOp_1 & (!cuifaluOp_0 & (!\Selector2~2_combout  & !\ShiftRight0~61_combout )))

	.dataa(cuifaluOp_1),
	.datab(cuifaluOp_0),
	.datac(\Selector2~2_combout ),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\Selector2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~12 .lut_mask = 16'h0001;
defparam \Selector2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N10
cycloneive_lcell_comb \Selector2~3 (
// Equation(s):
// \Selector2~3_combout  = (\Selector0~25_combout  & (\ShiftRight0~107_combout  & (!\Mux32~4_combout  & !\ShiftRight0~61_combout )))

	.dataa(\Selector0~25_combout ),
	.datab(\ShiftRight0~107_combout ),
	.datac(Mux32),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\Selector2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~3 .lut_mask = 16'h0008;
defparam \Selector2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N2
cycloneive_lcell_comb \ShiftLeft0~70 (
// Equation(s):
// \ShiftLeft0~70_combout  = (\Mux33~3_combout  & ((ShiftLeft01))) # (!\Mux33~3_combout  & (\Selector10~0_combout ))

	.dataa(\Selector10~0_combout ),
	.datab(gnd),
	.datac(Mux33),
	.datad(ShiftLeft01),
	.cin(gnd),
	.combout(\ShiftLeft0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~70 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N2
cycloneive_lcell_comb \Selector0~29 (
// Equation(s):
// \Selector0~29_combout  = (\Mux32~4_combout  & (!cuifaluOp_0 & \Selector0~21_combout ))

	.dataa(Mux32),
	.datab(gnd),
	.datac(cuifaluOp_0),
	.datad(\Selector0~21_combout ),
	.cin(gnd),
	.combout(\Selector0~29_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~29 .lut_mask = 16'h0A00;
defparam \Selector0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N20
cycloneive_lcell_comb \Selector2~4 (
// Equation(s):
// \Selector2~4_combout  = (\Selector2~3_combout  & ((\ShiftRight0~75_combout ) # ((\ShiftLeft0~70_combout  & \Selector0~29_combout )))) # (!\Selector2~3_combout  & (\ShiftLeft0~70_combout  & (\Selector0~29_combout )))

	.dataa(\Selector2~3_combout ),
	.datab(\ShiftLeft0~70_combout ),
	.datac(\Selector0~29_combout ),
	.datad(\ShiftRight0~75_combout ),
	.cin(gnd),
	.combout(\Selector2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~4 .lut_mask = 16'hEAC0;
defparam \Selector2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N24
cycloneive_lcell_comb \Selector2~5 (
// Equation(s):
// \Selector2~5_combout  = (Mux2 & ((\Mux7~1_combout  & (\Selector0~16_combout )) # (!\Mux7~1_combout  & ((\Selector0~17_combout ))))) # (!Mux2 & (((\Selector0~17_combout ) # (!\Mux7~1_combout ))))

	.dataa(Mux2),
	.datab(\Selector0~16_combout ),
	.datac(\Selector0~17_combout ),
	.datad(Mux7),
	.cin(gnd),
	.combout(\Selector2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~5 .lut_mask = 16'hD8F5;
defparam \Selector2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N12
cycloneive_lcell_comb \Selector2~7 (
// Equation(s):
// \Selector2~7_combout  = (\Selector2~6_combout  & ((\Selector0~15_combout ) # (\Selector2~5_combout )))

	.dataa(\Selector2~6_combout ),
	.datab(gnd),
	.datac(\Selector0~15_combout ),
	.datad(\Selector2~5_combout ),
	.cin(gnd),
	.combout(\Selector2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~7 .lut_mask = 16'hAAA0;
defparam \Selector2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N12
cycloneive_lcell_comb \Selector2~8 (
// Equation(s):
// \Selector2~8_combout  = (\Add1~58_combout  & \Selector0~19_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\Add1~58_combout ),
	.datad(\Selector0~19_combout ),
	.cin(gnd),
	.combout(\Selector2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~8 .lut_mask = 16'hF000;
defparam \Selector2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N14
cycloneive_lcell_comb \Selector2~9 (
// Equation(s):
// \Selector2~9_combout  = (\Selector2~7_combout ) # ((\Selector2~8_combout ) # ((\Selector0~20_combout  & \Add0~58_combout )))

	.dataa(\Selector2~7_combout ),
	.datab(\Selector0~20_combout ),
	.datac(\Add0~58_combout ),
	.datad(\Selector2~8_combout ),
	.cin(gnd),
	.combout(\Selector2~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~9 .lut_mask = 16'hFFEA;
defparam \Selector2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N22
cycloneive_lcell_comb \ShiftLeft0~118 (
// Equation(s):
// \ShiftLeft0~118_combout  = (\Mux35~3_combout  & (\ShiftLeft0~55_combout )) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & (\ShiftLeft0~55_combout )) # (!\Mux35~2_combout  & ((\ShiftLeft0~56_combout )))))

	.dataa(\ShiftLeft0~55_combout ),
	.datab(Mux351),
	.datac(Mux35),
	.datad(\ShiftLeft0~56_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~118_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~118 .lut_mask = 16'hABA8;
defparam \ShiftLeft0~118 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N24
cycloneive_lcell_comb \ShiftLeft0~117 (
// Equation(s):
// \ShiftLeft0~117_combout  = (\Mux35~2_combout  & (((\ShiftLeft0~64_combout )))) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & (\ShiftLeft0~64_combout )) # (!\Mux35~3_combout  & ((\ShiftLeft0~54_combout )))))

	.dataa(Mux35),
	.datab(Mux351),
	.datac(\ShiftLeft0~64_combout ),
	.datad(\ShiftLeft0~54_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~117_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~117 .lut_mask = 16'hF1E0;
defparam \ShiftLeft0~117 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N20
cycloneive_lcell_comb \ShiftLeft0~71 (
// Equation(s):
// \ShiftLeft0~71_combout  = (\Mux34~3_combout  & ((\ShiftLeft0~117_combout ))) # (!\Mux34~3_combout  & (\ShiftLeft0~118_combout ))

	.dataa(Mux34),
	.datab(gnd),
	.datac(\ShiftLeft0~118_combout ),
	.datad(\ShiftLeft0~117_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~71 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N8
cycloneive_lcell_comb \ShiftLeft0~116 (
// Equation(s):
// \ShiftLeft0~116_combout  = (\Mux35~2_combout  & (((\ShiftLeft0~57_combout )))) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & (\ShiftLeft0~57_combout )) # (!\Mux35~3_combout  & ((\ShiftLeft0~67_combout )))))

	.dataa(Mux35),
	.datab(Mux351),
	.datac(\ShiftLeft0~57_combout ),
	.datad(\ShiftLeft0~67_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~116_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~116 .lut_mask = 16'hF1E0;
defparam \ShiftLeft0~116 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N16
cycloneive_lcell_comb \ShiftLeft0~66 (
// Equation(s):
// \ShiftLeft0~66_combout  = (\Mux36~4_combout  & ((Mux3))) # (!\Mux36~4_combout  & (Mux2))

	.dataa(Mux2),
	.datab(Mux36),
	.datac(Mux3),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~66 .lut_mask = 16'hE2E2;
defparam \ShiftLeft0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N14
cycloneive_lcell_comb \Selector2~10 (
// Equation(s):
// \Selector2~10_combout  = (\ShiftRight0~107_combout  & (!\Selector2~14_combout  & ((\ShiftLeft0~66_combout )))) # (!\ShiftRight0~107_combout  & ((\Selector2~14_combout ) # ((\ShiftLeft0~116_combout ))))

	.dataa(\ShiftRight0~107_combout ),
	.datab(\Selector2~14_combout ),
	.datac(\ShiftLeft0~116_combout ),
	.datad(\ShiftLeft0~66_combout ),
	.cin(gnd),
	.combout(\Selector2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~10 .lut_mask = 16'h7654;
defparam \Selector2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N28
cycloneive_lcell_comb \Selector2~11 (
// Equation(s):
// \Selector2~11_combout  = (\Selector2~14_combout  & ((\Selector2~10_combout  & (\ShiftLeft0~71_combout )) # (!\Selector2~10_combout  & ((\ShiftLeft0~68_combout ))))) # (!\Selector2~14_combout  & (((\Selector2~10_combout ))))

	.dataa(\ShiftLeft0~71_combout ),
	.datab(\Selector2~14_combout ),
	.datac(\ShiftLeft0~68_combout ),
	.datad(\Selector2~10_combout ),
	.cin(gnd),
	.combout(\Selector2~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~11 .lut_mask = 16'hBBC0;
defparam \Selector2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N28
cycloneive_lcell_comb \ShiftLeft0~73 (
// Equation(s):
// \ShiftLeft0~73_combout  = (\ShiftLeft0~72_combout ) # ((\Mux36~4_combout  & (!\Mux35~4_combout  & Mux30)))

	.dataa(\ShiftLeft0~72_combout ),
	.datab(Mux36),
	.datac(Mux352),
	.datad(Mux301),
	.cin(gnd),
	.combout(\ShiftLeft0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~73 .lut_mask = 16'hAEAA;
defparam \ShiftLeft0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N18
cycloneive_lcell_comb \Selector29~11 (
// Equation(s):
// \Selector29~11_combout  = (!\Mux33~3_combout  & (!\Mux34~3_combout  & (\ShiftLeft0~73_combout  & \Selector16~0_combout )))

	.dataa(Mux33),
	.datab(Mux34),
	.datac(\ShiftLeft0~73_combout ),
	.datad(\Selector16~0_combout ),
	.cin(gnd),
	.combout(\Selector29~11_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~11 .lut_mask = 16'h1000;
defparam \Selector29~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N2
cycloneive_lcell_comb \ShiftRight0~152 (
// Equation(s):
// \ShiftRight0~152_combout  = (\Mux35~3_combout  & (((\ShiftRight0~99_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftRight0~99_combout ))) # (!\Mux35~2_combout  & (\ShiftRight0~101_combout ))))

	.dataa(Mux351),
	.datab(\ShiftRight0~101_combout ),
	.datac(Mux35),
	.datad(\ShiftRight0~99_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~152_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~152 .lut_mask = 16'hFE04;
defparam \ShiftRight0~152 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N18
cycloneive_lcell_comb \ShiftRight0~153 (
// Equation(s):
// \ShiftRight0~153_combout  = (\Mux35~2_combout  & (((\ShiftRight0~102_combout )))) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & ((\ShiftRight0~102_combout ))) # (!\Mux35~3_combout  & (\ShiftRight0~103_combout ))))

	.dataa(\ShiftRight0~103_combout ),
	.datab(Mux35),
	.datac(Mux351),
	.datad(\ShiftRight0~102_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~153_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~153 .lut_mask = 16'hFE02;
defparam \ShiftRight0~153 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N22
cycloneive_lcell_comb \Selector21~0 (
// Equation(s):
// \Selector21~0_combout  = (\Mux34~3_combout  & (\ShiftRight0~152_combout )) # (!\Mux34~3_combout  & ((\ShiftRight0~153_combout )))

	.dataa(Mux34),
	.datab(gnd),
	.datac(\ShiftRight0~152_combout ),
	.datad(\ShiftRight0~153_combout ),
	.cin(gnd),
	.combout(\Selector21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~0 .lut_mask = 16'hF5A0;
defparam \Selector21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N0
cycloneive_lcell_comb \ShiftRight0~151 (
// Equation(s):
// \ShiftRight0~151_combout  = (\Mux35~3_combout  & (((\ShiftRight0~97_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftRight0~97_combout ))) # (!\Mux35~2_combout  & (\ShiftRight0~98_combout ))))

	.dataa(Mux351),
	.datab(\ShiftRight0~98_combout ),
	.datac(Mux35),
	.datad(\ShiftRight0~97_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~151_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~151 .lut_mask = 16'hFE04;
defparam \ShiftRight0~151 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N22
cycloneive_lcell_comb \ShiftRight0~113 (
// Equation(s):
// \ShiftRight0~113_combout  = (\Mux34~3_combout  & (\ShiftRight0~96_combout  & (!\Mux35~4_combout ))) # (!\Mux34~3_combout  & (((\ShiftRight0~151_combout ))))

	.dataa(Mux34),
	.datab(\ShiftRight0~96_combout ),
	.datac(Mux352),
	.datad(\ShiftRight0~151_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~113_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~113 .lut_mask = 16'h5D08;
defparam \ShiftRight0~113 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N8
cycloneive_lcell_comb \ShiftRight0~114 (
// Equation(s):
// \ShiftRight0~114_combout  = (\Mux33~3_combout  & ((\ShiftRight0~113_combout ))) # (!\Mux33~3_combout  & (\Selector21~0_combout ))

	.dataa(Mux33),
	.datab(gnd),
	.datac(\Selector21~0_combout ),
	.datad(\ShiftRight0~113_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~114_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~114 .lut_mask = 16'hFA50;
defparam \ShiftRight0~114 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N8
cycloneive_lcell_comb \Selector29~3 (
// Equation(s):
// \Selector29~3_combout  = (\Mux34~3_combout  & ((\Selector29~2_combout ) # ((\Selector0~17_combout  & !Mux29)))) # (!\Mux34~3_combout  & (((\Selector0~17_combout  & Mux29))))

	.dataa(\Selector29~2_combout ),
	.datab(\Selector0~17_combout ),
	.datac(Mux34),
	.datad(Mux291),
	.cin(gnd),
	.combout(\Selector29~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~3 .lut_mask = 16'hACE0;
defparam \Selector29~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N30
cycloneive_lcell_comb \ShiftRight0~150 (
// Equation(s):
// \ShiftRight0~150_combout  = (\Mux35~2_combout  & (((\ShiftRight0~91_combout )))) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & ((\ShiftRight0~91_combout ))) # (!\Mux35~3_combout  & (\ShiftRight0~92_combout ))))

	.dataa(Mux35),
	.datab(\ShiftRight0~92_combout ),
	.datac(\ShiftRight0~91_combout ),
	.datad(Mux351),
	.cin(gnd),
	.combout(\ShiftRight0~150_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~150 .lut_mask = 16'hF0E4;
defparam \ShiftRight0~150 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N30
cycloneive_lcell_comb \ShiftRight0~149 (
// Equation(s):
// \ShiftRight0~149_combout  = (\Mux35~3_combout  & (\ShiftRight0~104_combout )) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & (\ShiftRight0~104_combout )) # (!\Mux35~2_combout  & ((\ShiftRight0~90_combout )))))

	.dataa(Mux351),
	.datab(\ShiftRight0~104_combout ),
	.datac(Mux35),
	.datad(\ShiftRight0~90_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~149_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~149 .lut_mask = 16'hCDC8;
defparam \ShiftRight0~149 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N20
cycloneive_lcell_comb \ShiftRight0~112 (
// Equation(s):
// \ShiftRight0~112_combout  = (\Mux34~3_combout  & ((\ShiftRight0~149_combout ))) # (!\Mux34~3_combout  & (\ShiftRight0~150_combout ))

	.dataa(Mux34),
	.datab(gnd),
	.datac(\ShiftRight0~150_combout ),
	.datad(\ShiftRight0~149_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~112_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~112 .lut_mask = 16'hFA50;
defparam \ShiftRight0~112 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N6
cycloneive_lcell_comb \ShiftRight0~148 (
// Equation(s):
// \ShiftRight0~148_combout  = (\Mux35~2_combout  & (((\ShiftRight0~93_combout )))) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & (\ShiftRight0~93_combout )) # (!\Mux35~3_combout  & ((\ShiftRight0~87_combout )))))

	.dataa(Mux35),
	.datab(Mux351),
	.datac(\ShiftRight0~93_combout ),
	.datad(\ShiftRight0~87_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~148_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~148 .lut_mask = 16'hF1E0;
defparam \ShiftRight0~148 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N24
cycloneive_lcell_comb \Selector29~7 (
// Equation(s):
// \Selector29~7_combout  = (\ShiftRight0~107_combout  & (!\Selector2~14_combout  & (\ShiftRight0~85_combout ))) # (!\ShiftRight0~107_combout  & ((\Selector2~14_combout ) # ((\ShiftRight0~148_combout ))))

	.dataa(\ShiftRight0~107_combout ),
	.datab(\Selector2~14_combout ),
	.datac(\ShiftRight0~85_combout ),
	.datad(\ShiftRight0~148_combout ),
	.cin(gnd),
	.combout(\Selector29~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~7 .lut_mask = 16'h7564;
defparam \Selector29~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N10
cycloneive_lcell_comb \Selector29~8 (
// Equation(s):
// \Selector29~8_combout  = (\Selector2~14_combout  & ((\Selector29~7_combout  & ((\ShiftRight0~112_combout ))) # (!\Selector29~7_combout  & (\ShiftRight0~88_combout )))) # (!\Selector2~14_combout  & (((\Selector29~7_combout ))))

	.dataa(\ShiftRight0~88_combout ),
	.datab(\Selector2~14_combout ),
	.datac(\ShiftRight0~112_combout ),
	.datad(\Selector29~7_combout ),
	.cin(gnd),
	.combout(\Selector29~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~8 .lut_mask = 16'hF388;
defparam \Selector29~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N30
cycloneive_lcell_comb \Selector29~4 (
// Equation(s):
// \Selector29~4_combout  = (\Selector0~18_combout  & (!\Mux34~3_combout  & !Mux29))

	.dataa(gnd),
	.datab(\Selector0~18_combout ),
	.datac(Mux34),
	.datad(Mux291),
	.cin(gnd),
	.combout(\Selector29~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~4 .lut_mask = 16'h000C;
defparam \Selector29~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N28
cycloneive_lcell_comb \Selector29~5 (
// Equation(s):
// \Selector29~5_combout  = (\Selector0~19_combout  & ((\Add1~4_combout ) # ((\Selector0~20_combout  & \Add0~4_combout )))) # (!\Selector0~19_combout  & (((\Selector0~20_combout  & \Add0~4_combout ))))

	.dataa(\Selector0~19_combout ),
	.datab(\Add1~4_combout ),
	.datac(\Selector0~20_combout ),
	.datad(\Add0~4_combout ),
	.cin(gnd),
	.combout(\Selector29~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~5 .lut_mask = 16'hF888;
defparam \Selector29~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N18
cycloneive_lcell_comb \Selector29~6 (
// Equation(s):
// \Selector29~6_combout  = (\Selector29~4_combout ) # ((\Selector29~5_combout ) # ((\Selector0~15_combout  & Mux29)))

	.dataa(\Selector0~15_combout ),
	.datab(Mux291),
	.datac(\Selector29~4_combout ),
	.datad(\Selector29~5_combout ),
	.cin(gnd),
	.combout(\Selector29~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~6 .lut_mask = 16'hFFF8;
defparam \Selector29~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N0
cycloneive_lcell_comb \Selector29~9 (
// Equation(s):
// \Selector29~9_combout  = (\Selector29~3_combout ) # ((\Selector29~6_combout ) # ((\Selector28~7_combout  & \Selector29~8_combout )))

	.dataa(\Selector28~7_combout ),
	.datab(\Selector29~3_combout ),
	.datac(\Selector29~8_combout ),
	.datad(\Selector29~6_combout ),
	.cin(gnd),
	.combout(\Selector29~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector29~9 .lut_mask = 16'hFFEC;
defparam \Selector29~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N6
cycloneive_lcell_comb \Selector5~6 (
// Equation(s):
// \Selector5~6_combout  = (Mux5 & ((\Selector0~8_combout ) # ((\Mux10~1_combout  & \Selector0~9_combout ))))

	.dataa(Mux102),
	.datab(\Selector0~8_combout ),
	.datac(\Selector0~9_combout ),
	.datad(Mux52),
	.cin(gnd),
	.combout(\Selector5~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~6 .lut_mask = 16'hEC00;
defparam \Selector5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N28
cycloneive_lcell_comb \Selector5~7 (
// Equation(s):
// \Selector5~7_combout  = (\Selector0~10_combout  & (Mux5 $ (((\Mux5~1_combout ) # (\Mux10~0_combout )))))

	.dataa(Mux5),
	.datab(Mux52),
	.datac(Mux10),
	.datad(\Selector0~10_combout ),
	.cin(gnd),
	.combout(\Selector5~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~7 .lut_mask = 16'h3600;
defparam \Selector5~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N14
cycloneive_lcell_comb \Selector5~8 (
// Equation(s):
// \Selector5~8_combout  = (\Mux10~1_combout  & (\Selector0~8_combout )) # (!\Mux10~1_combout  & (((\Selector0~11_combout  & !Mux5))))

	.dataa(Mux102),
	.datab(\Selector0~8_combout ),
	.datac(\Selector0~11_combout ),
	.datad(Mux52),
	.cin(gnd),
	.combout(\Selector5~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~8 .lut_mask = 16'h88D8;
defparam \Selector5~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N0
cycloneive_lcell_comb \Selector5~5 (
// Equation(s):
// \Selector5~5_combout  = (\Selector0~12_combout  & ((\Add1~52_combout ) # ((\Selector0~13_combout  & \Add0~52_combout )))) # (!\Selector0~12_combout  & (\Selector0~13_combout  & (\Add0~52_combout )))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector0~13_combout ),
	.datac(\Add0~52_combout ),
	.datad(\Add1~52_combout ),
	.cin(gnd),
	.combout(\Selector5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~5 .lut_mask = 16'hEAC0;
defparam \Selector5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N4
cycloneive_lcell_comb \Selector5~9 (
// Equation(s):
// \Selector5~9_combout  = (\Selector5~6_combout ) # ((\Selector5~7_combout ) # ((\Selector5~8_combout ) # (\Selector5~5_combout )))

	.dataa(\Selector5~6_combout ),
	.datab(\Selector5~7_combout ),
	.datac(\Selector5~8_combout ),
	.datad(\Selector5~5_combout ),
	.cin(gnd),
	.combout(\Selector5~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~9 .lut_mask = 16'hFFFE;
defparam \Selector5~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N24
cycloneive_lcell_comb \Selector5~0 (
// Equation(s):
// \Selector5~0_combout  = (\Mux32~4_combout ) # ((\Mux34~3_combout  & !\Mux33~3_combout ))

	.dataa(Mux34),
	.datab(gnd),
	.datac(Mux32),
	.datad(Mux33),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~0 .lut_mask = 16'hF0FA;
defparam \Selector5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N22
cycloneive_lcell_comb \Selector5~1 (
// Equation(s):
// \Selector5~1_combout  = (\Mux32~4_combout ) # (\Mux33~3_combout )

	.dataa(Mux32),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux33),
	.cin(gnd),
	.combout(\Selector5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~1 .lut_mask = 16'hFFAA;
defparam \Selector5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N20
cycloneive_lcell_comb \ShiftLeft0~76 (
// Equation(s):
// \ShiftLeft0~76_combout  = (\Mux36~4_combout  & (Mux20)) # (!\Mux36~4_combout  & ((Mux19)))

	.dataa(gnd),
	.datab(Mux36),
	.datac(Mux201),
	.datad(Mux191),
	.cin(gnd),
	.combout(\ShiftLeft0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~76 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N10
cycloneive_lcell_comb \ShiftLeft0~77 (
// Equation(s):
// \ShiftLeft0~77_combout  = (\Mux36~4_combout  & ((Mux18))) # (!\Mux36~4_combout  & (Mux17))

	.dataa(gnd),
	.datab(Mux171),
	.datac(Mux36),
	.datad(Mux181),
	.cin(gnd),
	.combout(\ShiftLeft0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~77 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N28
cycloneive_lcell_comb \ShiftLeft0~120 (
// Equation(s):
// \ShiftLeft0~120_combout  = (\Mux35~3_combout  & (\ShiftLeft0~76_combout )) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & (\ShiftLeft0~76_combout )) # (!\Mux35~2_combout  & ((\ShiftLeft0~77_combout )))))

	.dataa(Mux351),
	.datab(\ShiftLeft0~76_combout ),
	.datac(\ShiftLeft0~77_combout ),
	.datad(Mux35),
	.cin(gnd),
	.combout(\ShiftLeft0~120_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~120 .lut_mask = 16'hCCD8;
defparam \ShiftLeft0~120 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N22
cycloneive_lcell_comb \ShiftLeft0~78 (
// Equation(s):
// \ShiftLeft0~78_combout  = (\Mux36~4_combout  & ((Mux16))) # (!\Mux36~4_combout  & (Mux15))

	.dataa(gnd),
	.datab(Mux152),
	.datac(Mux36),
	.datad(Mux161),
	.cin(gnd),
	.combout(\ShiftLeft0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~78 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N0
cycloneive_lcell_comb \ShiftLeft0~79 (
// Equation(s):
// \ShiftLeft0~79_combout  = (\Mux36~4_combout  & ((Mux14))) # (!\Mux36~4_combout  & (Mux13))

	.dataa(gnd),
	.datab(Mux131),
	.datac(Mux36),
	.datad(Mux141),
	.cin(gnd),
	.combout(\ShiftLeft0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~79 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N20
cycloneive_lcell_comb \ShiftLeft0~121 (
// Equation(s):
// \ShiftLeft0~121_combout  = (\Mux35~3_combout  & (((\ShiftLeft0~78_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & (\ShiftLeft0~78_combout )) # (!\Mux35~2_combout  & ((\ShiftLeft0~79_combout )))))

	.dataa(Mux351),
	.datab(Mux35),
	.datac(\ShiftLeft0~78_combout ),
	.datad(\ShiftLeft0~79_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~121_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~121 .lut_mask = 16'hF1E0;
defparam \ShiftLeft0~121 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N28
cycloneive_lcell_comb \ShiftLeft0~80 (
// Equation(s):
// \ShiftLeft0~80_combout  = (\Mux34~3_combout  & (\ShiftLeft0~120_combout )) # (!\Mux34~3_combout  & ((\ShiftLeft0~121_combout )))

	.dataa(gnd),
	.datab(Mux34),
	.datac(\ShiftLeft0~120_combout ),
	.datad(\ShiftLeft0~121_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~80 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N10
cycloneive_lcell_comb \Selector5~2 (
// Equation(s):
// \Selector5~2_combout  = (\Selector5~0_combout  & (((\Selector5~1_combout )))) # (!\Selector5~0_combout  & ((\Selector5~1_combout  & ((\ShiftLeft0~80_combout ))) # (!\Selector5~1_combout  & (\ShiftLeft0~122_combout ))))

	.dataa(\ShiftLeft0~122_combout ),
	.datab(\Selector5~0_combout ),
	.datac(\Selector5~1_combout ),
	.datad(\ShiftLeft0~80_combout ),
	.cin(gnd),
	.combout(\Selector5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~2 .lut_mask = 16'hF2C2;
defparam \Selector5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N30
cycloneive_lcell_comb \ShiftLeft0~84 (
// Equation(s):
// \ShiftLeft0~84_combout  = (\Mux36~4_combout  & ((Mux26))) # (!\Mux36~4_combout  & (Mux25))

	.dataa(gnd),
	.datab(Mux251),
	.datac(Mux36),
	.datad(Mux261),
	.cin(gnd),
	.combout(\ShiftLeft0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~84 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N20
cycloneive_lcell_comb \ShiftLeft0~123 (
// Equation(s):
// \ShiftLeft0~123_combout  = (\Mux35~2_combout  & (\ShiftLeft0~83_combout )) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & (\ShiftLeft0~83_combout )) # (!\Mux35~3_combout  & ((\ShiftLeft0~84_combout )))))

	.dataa(\ShiftLeft0~83_combout ),
	.datab(Mux35),
	.datac(\ShiftLeft0~84_combout ),
	.datad(Mux351),
	.cin(gnd),
	.combout(\ShiftLeft0~123_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~123 .lut_mask = 16'hAAB8;
defparam \ShiftLeft0~123 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N2
cycloneive_lcell_comb \ShiftLeft0~87 (
// Equation(s):
// \ShiftLeft0~87_combout  = (!\Mux33~3_combout  & ((\Mux34~3_combout  & ((\ShiftLeft0~123_combout ))) # (!\Mux34~3_combout  & (\ShiftLeft0~124_combout ))))

	.dataa(\ShiftLeft0~124_combout ),
	.datab(Mux33),
	.datac(Mux34),
	.datad(\ShiftLeft0~123_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~87_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~87 .lut_mask = 16'h3202;
defparam \ShiftLeft0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N0
cycloneive_lcell_comb \ShiftLeft0~88 (
// Equation(s):
// \ShiftLeft0~88_combout  = (\ShiftLeft0~87_combout ) # ((\Mux33~3_combout  & (\ShiftLeft0~73_combout  & !\Mux34~3_combout )))

	.dataa(Mux33),
	.datab(\ShiftLeft0~73_combout ),
	.datac(Mux34),
	.datad(\ShiftLeft0~87_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~88_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~88 .lut_mask = 16'hFF08;
defparam \ShiftLeft0~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N18
cycloneive_lcell_comb \Selector5~3 (
// Equation(s):
// \Selector5~3_combout  = (\Selector5~0_combout  & ((\Selector5~2_combout  & ((\ShiftLeft0~88_combout ))) # (!\Selector5~2_combout  & (\ShiftLeft0~119_combout )))) # (!\Selector5~0_combout  & (((\Selector5~2_combout ))))

	.dataa(\ShiftLeft0~119_combout ),
	.datab(\Selector5~0_combout ),
	.datac(\Selector5~2_combout ),
	.datad(\ShiftLeft0~88_combout ),
	.cin(gnd),
	.combout(\Selector5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~3 .lut_mask = 16'hF838;
defparam \Selector5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N2
cycloneive_lcell_comb \Selector5~4 (
// Equation(s):
// \Selector5~4_combout  = (!\ShiftRight0~61_combout  & (\Selector0~7_combout  & \Selector5~3_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~61_combout ),
	.datac(\Selector0~7_combout ),
	.datad(\Selector5~3_combout ),
	.cin(gnd),
	.combout(\Selector5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector5~4 .lut_mask = 16'h3000;
defparam \Selector5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N22
cycloneive_lcell_comb \ShiftLeft0~125 (
// Equation(s):
// \ShiftLeft0~125_combout  = (!\Mux35~2_combout  & (Mux31 & (!\Mux36~4_combout  & !\Mux35~3_combout )))

	.dataa(Mux35),
	.datab(Mux311),
	.datac(Mux36),
	.datad(Mux351),
	.cin(gnd),
	.combout(\ShiftLeft0~125_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~125 .lut_mask = 16'h0004;
defparam \ShiftLeft0~125 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N2
cycloneive_lcell_comb \ShiftLeft0~89 (
// Equation(s):
// \ShiftLeft0~89_combout  = (\Mux35~4_combout  & ((\Mux36~4_combout  & (Mux30)) # (!\Mux36~4_combout  & ((Mux29)))))

	.dataa(Mux301),
	.datab(Mux36),
	.datac(Mux291),
	.datad(Mux352),
	.cin(gnd),
	.combout(\ShiftLeft0~89_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~89 .lut_mask = 16'hB800;
defparam \ShiftLeft0~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N30
cycloneive_lcell_comb \ShiftLeft0~83 (
// Equation(s):
// \ShiftLeft0~83_combout  = (\Mux36~4_combout  & (Mux28)) # (!\Mux36~4_combout  & ((Mux27)))

	.dataa(gnd),
	.datab(Mux281),
	.datac(Mux36),
	.datad(Mux271),
	.cin(gnd),
	.combout(\ShiftLeft0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~83 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N0
cycloneive_lcell_comb \ShiftLeft0~126 (
// Equation(s):
// \ShiftLeft0~126_combout  = (\ShiftLeft0~89_combout ) # ((!\Mux35~3_combout  & (\ShiftLeft0~83_combout  & !\Mux35~2_combout )))

	.dataa(Mux351),
	.datab(\ShiftLeft0~89_combout ),
	.datac(\ShiftLeft0~83_combout ),
	.datad(Mux35),
	.cin(gnd),
	.combout(\ShiftLeft0~126_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~126 .lut_mask = 16'hCCDC;
defparam \ShiftLeft0~126 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N4
cycloneive_lcell_comb \ShiftLeft0~82 (
// Equation(s):
// \ShiftLeft0~82_combout  = (\Mux36~4_combout  & (Mux6)) # (!\Mux36~4_combout  & ((Mux5)))

	.dataa(gnd),
	.datab(Mux36),
	.datac(Mux61),
	.datad(Mux52),
	.cin(gnd),
	.combout(\ShiftLeft0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~82 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N2
cycloneive_lcell_comb \ShiftLeft0~81 (
// Equation(s):
// \ShiftLeft0~81_combout  = (\Mux36~4_combout  & ((Mux8))) # (!\Mux36~4_combout  & (Mux7))

	.dataa(Mux71),
	.datab(gnd),
	.datac(Mux36),
	.datad(Mux81),
	.cin(gnd),
	.combout(\ShiftLeft0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~81 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N30
cycloneive_lcell_comb \ShiftLeft0~75 (
// Equation(s):
// \ShiftLeft0~75_combout  = (\Mux36~4_combout  & ((Mux10))) # (!\Mux36~4_combout  & (Mux9))

	.dataa(Mux36),
	.datab(gnd),
	.datac(Mux91),
	.datad(Mux101),
	.cin(gnd),
	.combout(\ShiftLeft0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~75 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N26
cycloneive_lcell_comb \ShiftLeft0~129 (
// Equation(s):
// \ShiftLeft0~129_combout  = (\Mux35~3_combout  & (((\ShiftLeft0~75_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftLeft0~75_combout ))) # (!\Mux35~2_combout  & (\ShiftLeft0~81_combout ))))

	.dataa(Mux351),
	.datab(\ShiftLeft0~81_combout ),
	.datac(\ShiftLeft0~75_combout ),
	.datad(Mux35),
	.cin(gnd),
	.combout(\ShiftLeft0~129_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~129 .lut_mask = 16'hF0E4;
defparam \ShiftLeft0~129 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N0
cycloneive_lcell_comb \ShiftLeft0~92 (
// Equation(s):
// \ShiftLeft0~92_combout  = (\Mux36~4_combout  & (Mux4)) # (!\Mux36~4_combout  & ((Mux3)))

	.dataa(Mux4),
	.datab(gnd),
	.datac(Mux36),
	.datad(Mux3),
	.cin(gnd),
	.combout(\ShiftLeft0~92_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~92 .lut_mask = 16'hAFA0;
defparam \ShiftLeft0~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N22
cycloneive_lcell_comb \Selector3~6 (
// Equation(s):
// \Selector3~6_combout  = (\Selector2~14_combout  & (!\ShiftRight0~107_combout )) # (!\Selector2~14_combout  & ((\ShiftRight0~107_combout  & ((\ShiftLeft0~92_combout ))) # (!\ShiftRight0~107_combout  & (\ShiftLeft0~129_combout ))))

	.dataa(\Selector2~14_combout ),
	.datab(\ShiftRight0~107_combout ),
	.datac(\ShiftLeft0~129_combout ),
	.datad(\ShiftLeft0~92_combout ),
	.cin(gnd),
	.combout(\Selector3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~6 .lut_mask = 16'h7632;
defparam \Selector3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N30
cycloneive_lcell_comb \ShiftLeft0~130 (
// Equation(s):
// \ShiftLeft0~130_combout  = (\Mux35~3_combout  & (((\ShiftLeft0~77_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftLeft0~77_combout ))) # (!\Mux35~2_combout  & (\ShiftLeft0~78_combout ))))

	.dataa(Mux351),
	.datab(Mux35),
	.datac(\ShiftLeft0~78_combout ),
	.datad(\ShiftLeft0~77_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~130_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~130 .lut_mask = 16'hFE10;
defparam \ShiftLeft0~130 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N4
cycloneive_lcell_comb \ShiftLeft0~74 (
// Equation(s):
// \ShiftLeft0~74_combout  = (\Mux36~4_combout  & (Mux12)) # (!\Mux36~4_combout  & ((Mux11)))

	.dataa(Mux36),
	.datab(gnd),
	.datac(Mux121),
	.datad(Mux111),
	.cin(gnd),
	.combout(\ShiftLeft0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~74 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N0
cycloneive_lcell_comb \ShiftLeft0~131 (
// Equation(s):
// \ShiftLeft0~131_combout  = (\Mux35~3_combout  & (((\ShiftLeft0~79_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftLeft0~79_combout ))) # (!\Mux35~2_combout  & (\ShiftLeft0~74_combout ))))

	.dataa(Mux351),
	.datab(\ShiftLeft0~74_combout ),
	.datac(\ShiftLeft0~79_combout ),
	.datad(Mux35),
	.cin(gnd),
	.combout(\ShiftLeft0~131_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~131 .lut_mask = 16'hF0E4;
defparam \ShiftLeft0~131 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N12
cycloneive_lcell_comb \ShiftLeft0~93 (
// Equation(s):
// \ShiftLeft0~93_combout  = (\Mux34~3_combout  & (\ShiftLeft0~130_combout )) # (!\Mux34~3_combout  & ((\ShiftLeft0~131_combout )))

	.dataa(gnd),
	.datab(Mux34),
	.datac(\ShiftLeft0~130_combout ),
	.datad(\ShiftLeft0~131_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~93_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~93 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N26
cycloneive_lcell_comb \Selector3~7 (
// Equation(s):
// \Selector3~7_combout  = (\Selector2~14_combout  & ((\Selector3~6_combout  & ((\ShiftLeft0~93_combout ))) # (!\Selector3~6_combout  & (\ShiftLeft0~82_combout )))) # (!\Selector2~14_combout  & (((\Selector3~6_combout ))))

	.dataa(\Selector2~14_combout ),
	.datab(\ShiftLeft0~82_combout ),
	.datac(\Selector3~6_combout ),
	.datad(\ShiftLeft0~93_combout ),
	.cin(gnd),
	.combout(\Selector3~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~7 .lut_mask = 16'hF858;
defparam \Selector3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N16
cycloneive_lcell_comb \ShiftLeft0~86 (
// Equation(s):
// \ShiftLeft0~86_combout  = (\Mux36~4_combout  & ((Mux22))) # (!\Mux36~4_combout  & (Mux21))

	.dataa(gnd),
	.datab(Mux211),
	.datac(Mux36),
	.datad(Mux221),
	.cin(gnd),
	.combout(\ShiftLeft0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~86 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N16
cycloneive_lcell_comb \ShiftLeft0~128 (
// Equation(s):
// \ShiftLeft0~128_combout  = (\Mux35~3_combout  & (((\ShiftLeft0~86_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftLeft0~86_combout ))) # (!\Mux35~2_combout  & (\ShiftLeft0~76_combout ))))

	.dataa(Mux351),
	.datab(\ShiftLeft0~76_combout ),
	.datac(\ShiftLeft0~86_combout ),
	.datad(Mux35),
	.cin(gnd),
	.combout(\ShiftLeft0~128_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~128 .lut_mask = 16'hF0E4;
defparam \ShiftLeft0~128 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N6
cycloneive_lcell_comb \ShiftLeft0~85 (
// Equation(s):
// \ShiftLeft0~85_combout  = (\Mux36~4_combout  & ((Mux24))) # (!\Mux36~4_combout  & (Mux23))

	.dataa(gnd),
	.datab(Mux36),
	.datac(Mux231),
	.datad(Mux241),
	.cin(gnd),
	.combout(\ShiftLeft0~85_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~85 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N10
cycloneive_lcell_comb \ShiftLeft0~127 (
// Equation(s):
// \ShiftLeft0~127_combout  = (\Mux35~3_combout  & (((\ShiftLeft0~84_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftLeft0~84_combout ))) # (!\Mux35~2_combout  & (\ShiftLeft0~85_combout ))))

	.dataa(Mux351),
	.datab(Mux35),
	.datac(\ShiftLeft0~85_combout ),
	.datad(\ShiftLeft0~84_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~127_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~127 .lut_mask = 16'hFE10;
defparam \ShiftLeft0~127 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N6
cycloneive_lcell_comb \Selector11~0 (
// Equation(s):
// \Selector11~0_combout  = (\Mux34~3_combout  & ((\ShiftLeft0~127_combout ))) # (!\Mux34~3_combout  & (\ShiftLeft0~128_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~128_combout ),
	.datac(Mux34),
	.datad(\ShiftLeft0~127_combout ),
	.cin(gnd),
	.combout(\Selector11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~0 .lut_mask = 16'hFC0C;
defparam \Selector11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N26
cycloneive_lcell_comb \ShiftLeft0~91 (
// Equation(s):
// \ShiftLeft0~91_combout  = (\Mux33~3_combout  & ((ShiftLeft02))) # (!\Mux33~3_combout  & (\Selector11~0_combout ))

	.dataa(gnd),
	.datab(Mux33),
	.datac(\Selector11~0_combout ),
	.datad(ShiftLeft02),
	.cin(gnd),
	.combout(\ShiftLeft0~91_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~91 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N8
cycloneive_lcell_comb \Selector3~0 (
// Equation(s):
// \Selector3~0_combout  = (\ShiftRight0~137_combout  & ((\Selector2~3_combout ) # ((\Selector0~29_combout  & \ShiftLeft0~91_combout )))) # (!\ShiftRight0~137_combout  & (\Selector0~29_combout  & ((\ShiftLeft0~91_combout ))))

	.dataa(\ShiftRight0~137_combout ),
	.datab(\Selector0~29_combout ),
	.datac(\Selector2~3_combout ),
	.datad(\ShiftLeft0~91_combout ),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~0 .lut_mask = 16'hECA0;
defparam \Selector3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N12
cycloneive_lcell_comb \Selector3~4 (
// Equation(s):
// \Selector3~4_combout  = (\Mux8~1_combout  & (((\Selector0~15_combout )))) # (!\Mux8~1_combout  & (\Selector0~18_combout  & ((!Mux3))))

	.dataa(\Selector0~18_combout ),
	.datab(\Selector0~15_combout ),
	.datac(Mux3),
	.datad(Mux82),
	.cin(gnd),
	.combout(\Selector3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~4 .lut_mask = 16'hCC0A;
defparam \Selector3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N16
cycloneive_lcell_comb \Selector3~2 (
// Equation(s):
// \Selector3~2_combout  = (Mux3 & ((\Selector0~15_combout ) # ((\Selector0~16_combout  & \Mux8~1_combout ))))

	.dataa(\Selector0~16_combout ),
	.datab(\Selector0~15_combout ),
	.datac(Mux3),
	.datad(Mux82),
	.cin(gnd),
	.combout(\Selector3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~2 .lut_mask = 16'hE0C0;
defparam \Selector3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N22
cycloneive_lcell_comb \Selector3~3 (
// Equation(s):
// \Selector3~3_combout  = (\Selector0~17_combout  & (Mux3 $ (((\Mux5~1_combout ) # (\Mux8~0_combout )))))

	.dataa(\Selector0~17_combout ),
	.datab(Mux3),
	.datac(Mux5),
	.datad(Mux8),
	.cin(gnd),
	.combout(\Selector3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~3 .lut_mask = 16'h2228;
defparam \Selector3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N18
cycloneive_lcell_comb \Selector3~1 (
// Equation(s):
// \Selector3~1_combout  = (\Selector0~20_combout  & ((\Add0~56_combout ) # ((\Add1~56_combout  & \Selector0~19_combout )))) # (!\Selector0~20_combout  & (\Add1~56_combout  & (\Selector0~19_combout )))

	.dataa(\Selector0~20_combout ),
	.datab(\Add1~56_combout ),
	.datac(\Selector0~19_combout ),
	.datad(\Add0~56_combout ),
	.cin(gnd),
	.combout(\Selector3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~1 .lut_mask = 16'hEAC0;
defparam \Selector3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N10
cycloneive_lcell_comb \Selector3~5 (
// Equation(s):
// \Selector3~5_combout  = (\Selector3~4_combout ) # ((\Selector3~2_combout ) # ((\Selector3~3_combout ) # (\Selector3~1_combout )))

	.dataa(\Selector3~4_combout ),
	.datab(\Selector3~2_combout ),
	.datac(\Selector3~3_combout ),
	.datad(\Selector3~1_combout ),
	.cin(gnd),
	.combout(\Selector3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~5 .lut_mask = 16'hFFFE;
defparam \Selector3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N2
cycloneive_lcell_comb \Selector0~30 (
// Equation(s):
// \Selector0~30_combout  = (\Mux35~3_combout ) # ((\Mux35~2_combout ) # (\Mux34~3_combout ))

	.dataa(Mux351),
	.datab(gnd),
	.datac(Mux35),
	.datad(Mux34),
	.cin(gnd),
	.combout(\Selector0~30_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~30 .lut_mask = 16'hFFFA;
defparam \Selector0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N26
cycloneive_lcell_comb \Selector1~0 (
// Equation(s):
// \Selector1~0_combout  = (!\Selector0~30_combout  & (!\Mux33~3_combout  & (\ShiftRight0~96_combout  & \Selector8~0_combout )))

	.dataa(\Selector0~30_combout ),
	.datab(Mux33),
	.datac(\ShiftRight0~96_combout ),
	.datad(\Selector8~0_combout ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~0 .lut_mask = 16'h1000;
defparam \Selector1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N12
cycloneive_lcell_comb \Selector1~9 (
// Equation(s):
// \Selector1~9_combout  = (Mux1 & ((\Selector0~15_combout ) # ((\Selector0~16_combout  & \Mux6~1_combout ))))

	.dataa(\Selector0~15_combout ),
	.datab(\Selector0~16_combout ),
	.datac(Mux1),
	.datad(Mux62),
	.cin(gnd),
	.combout(\Selector1~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~9 .lut_mask = 16'hE0A0;
defparam \Selector1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N8
cycloneive_lcell_comb \Selector1~2 (
// Equation(s):
// \Selector1~2_combout  = (\Mux6~1_combout  & (((\Selector0~15_combout )))) # (!\Mux6~1_combout  & (\Selector0~18_combout  & (!Mux1)))

	.dataa(\Selector0~18_combout ),
	.datab(Mux1),
	.datac(\Selector0~15_combout ),
	.datad(Mux62),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~2 .lut_mask = 16'hF022;
defparam \Selector1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N30
cycloneive_lcell_comb \ShiftLeft0~122 (
// Equation(s):
// \ShiftLeft0~122_combout  = (\Mux35~3_combout  & (\ShiftLeft0~81_combout )) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & (\ShiftLeft0~81_combout )) # (!\Mux35~2_combout  & ((\ShiftLeft0~82_combout )))))

	.dataa(Mux351),
	.datab(\ShiftLeft0~81_combout ),
	.datac(\ShiftLeft0~82_combout ),
	.datad(Mux35),
	.cin(gnd),
	.combout(\ShiftLeft0~122_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~122 .lut_mask = 16'hCCD8;
defparam \ShiftLeft0~122 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N20
cycloneive_lcell_comb \Selector1~3 (
// Equation(s):
// \Selector1~3_combout  = (\Selector0~30_combout  & ((\ShiftLeft0~92_combout ) # ((\Selector0~41_combout )))) # (!\Selector0~30_combout  & (((!\Selector0~41_combout  & Mux1))))

	.dataa(\Selector0~30_combout ),
	.datab(\ShiftLeft0~92_combout ),
	.datac(\Selector0~41_combout ),
	.datad(Mux1),
	.cin(gnd),
	.combout(\Selector1~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~3 .lut_mask = 16'hADA8;
defparam \Selector1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N18
cycloneive_lcell_comb \Selector1~4 (
// Equation(s):
// \Selector1~4_combout  = (\Selector0~41_combout  & ((\Selector1~3_combout  & ((\ShiftLeft0~122_combout ))) # (!\Selector1~3_combout  & (Mux2)))) # (!\Selector0~41_combout  & (((\Selector1~3_combout ))))

	.dataa(Mux2),
	.datab(\Selector0~41_combout ),
	.datac(\ShiftLeft0~122_combout ),
	.datad(\Selector1~3_combout ),
	.cin(gnd),
	.combout(\Selector1~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~4 .lut_mask = 16'hF388;
defparam \Selector1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N16
cycloneive_lcell_comb \Selector1~5 (
// Equation(s):
// \Selector1~5_combout  = (!cuifaluOp_0 & (\Selector16~1_combout  & \Selector1~4_combout ))

	.dataa(gnd),
	.datab(cuifaluOp_0),
	.datac(\Selector16~1_combout ),
	.datad(\Selector1~4_combout ),
	.cin(gnd),
	.combout(\Selector1~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~5 .lut_mask = 16'h3000;
defparam \Selector1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y43_N10
cycloneive_lcell_comb \ShiftLeft0~119 (
// Equation(s):
// \ShiftLeft0~119_combout  = (\Mux35~3_combout  & (\ShiftLeft0~74_combout )) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & (\ShiftLeft0~74_combout )) # (!\Mux35~2_combout  & ((\ShiftLeft0~75_combout )))))

	.dataa(Mux351),
	.datab(\ShiftLeft0~74_combout ),
	.datac(\ShiftLeft0~75_combout ),
	.datad(Mux35),
	.cin(gnd),
	.combout(\ShiftLeft0~119_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~119 .lut_mask = 16'hCCD8;
defparam \ShiftLeft0~119 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N8
cycloneive_lcell_comb \Selector1~6 (
// Equation(s):
// \Selector1~6_combout  = (\Mux34~3_combout  & ((\ShiftLeft0~121_combout ))) # (!\Mux34~3_combout  & (\ShiftLeft0~119_combout ))

	.dataa(Mux34),
	.datab(gnd),
	.datac(\ShiftLeft0~119_combout ),
	.datad(\ShiftLeft0~121_combout ),
	.cin(gnd),
	.combout(\Selector1~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~6 .lut_mask = 16'hFA50;
defparam \Selector1~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N20
cycloneive_lcell_comb \Selector0~27 (
// Equation(s):
// \Selector0~27_combout  = (!\Mux32~4_combout  & (\Mux33~3_combout  & (!cuifaluOp_0 & \Selector0~21_combout )))

	.dataa(Mux32),
	.datab(Mux33),
	.datac(cuifaluOp_0),
	.datad(\Selector0~21_combout ),
	.cin(gnd),
	.combout(\Selector0~27_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~27 .lut_mask = 16'h0400;
defparam \Selector0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N4
cycloneive_lcell_comb \Selector1~7 (
// Equation(s):
// \Selector1~7_combout  = (\ShiftLeft0~95_combout  & ((\Selector0~29_combout ) # ((\Selector1~6_combout  & \Selector0~27_combout )))) # (!\ShiftLeft0~95_combout  & (\Selector1~6_combout  & (\Selector0~27_combout )))

	.dataa(\ShiftLeft0~95_combout ),
	.datab(\Selector1~6_combout ),
	.datac(\Selector0~27_combout ),
	.datad(\Selector0~29_combout ),
	.cin(gnd),
	.combout(\Selector1~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~7 .lut_mask = 16'hEAC0;
defparam \Selector1~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N18
cycloneive_lcell_comb \Selector1~8 (
// Equation(s):
// \Selector1~8_combout  = (\Selector1~1_combout ) # ((\Selector1~2_combout ) # ((\Selector1~5_combout ) # (\Selector1~7_combout )))

	.dataa(\Selector1~1_combout ),
	.datab(\Selector1~2_combout ),
	.datac(\Selector1~5_combout ),
	.datad(\Selector1~7_combout ),
	.cin(gnd),
	.combout(\Selector1~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~8 .lut_mask = 16'hFFFE;
defparam \Selector1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N14
cycloneive_lcell_comb \Selector1~10 (
// Equation(s):
// \Selector1~10_combout  = (\Selector1~9_combout ) # ((\Selector1~8_combout ) # ((\Selector0~19_combout  & \Add1~60_combout )))

	.dataa(\Selector1~9_combout ),
	.datab(\Selector0~19_combout ),
	.datac(\Add1~60_combout ),
	.datad(\Selector1~8_combout ),
	.cin(gnd),
	.combout(\Selector1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector1~10 .lut_mask = 16'hFFEA;
defparam \Selector1~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N8
cycloneive_lcell_comb \ShiftLeft0~96 (
// Equation(s):
// \ShiftLeft0~96_combout  = (\Mux34~3_combout  & (\ShiftLeft0~111_combout )) # (!\Mux34~3_combout  & ((\ShiftLeft0~107_combout )))

	.dataa(Mux34),
	.datab(\ShiftLeft0~111_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~107_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~96_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~96 .lut_mask = 16'hDD88;
defparam \ShiftLeft0~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N16
cycloneive_lcell_comb \ShiftLeft0~61 (
// Equation(s):
// \ShiftLeft0~61_combout  = (\Mux36~4_combout  & ((Mux23))) # (!\Mux36~4_combout  & (Mux22))

	.dataa(Mux221),
	.datab(gnd),
	.datac(Mux36),
	.datad(Mux231),
	.cin(gnd),
	.combout(\ShiftLeft0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~61 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N18
cycloneive_lcell_comb \ShiftLeft0~62 (
// Equation(s):
// \ShiftLeft0~62_combout  = (\Mux36~4_combout  & (Mux21)) # (!\Mux36~4_combout  & ((Mux20)))

	.dataa(gnd),
	.datab(Mux36),
	.datac(Mux211),
	.datad(Mux201),
	.cin(gnd),
	.combout(\ShiftLeft0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~62 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N26
cycloneive_lcell_comb \ShiftLeft0~110 (
// Equation(s):
// \ShiftLeft0~110_combout  = (\Mux35~3_combout  & (((\ShiftLeft0~61_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & (\ShiftLeft0~61_combout )) # (!\Mux35~2_combout  & ((\ShiftLeft0~62_combout )))))

	.dataa(Mux351),
	.datab(Mux35),
	.datac(\ShiftLeft0~61_combout ),
	.datad(\ShiftLeft0~62_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~110_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~110 .lut_mask = 16'hF1E0;
defparam \ShiftLeft0~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N8
cycloneive_lcell_comb \ShiftLeft0~97 (
// Equation(s):
// \ShiftLeft0~97_combout  = (!\Mux33~3_combout  & ((\Mux34~3_combout  & ((\ShiftLeft0~109_combout ))) # (!\Mux34~3_combout  & (\ShiftLeft0~110_combout ))))

	.dataa(Mux33),
	.datab(Mux34),
	.datac(\ShiftLeft0~110_combout ),
	.datad(\ShiftLeft0~109_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~97_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~97 .lut_mask = 16'h5410;
defparam \ShiftLeft0~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N6
cycloneive_lcell_comb \ShiftLeft0~98 (
// Equation(s):
// \ShiftLeft0~98_combout  = (\ShiftLeft0~97_combout ) # ((\Mux33~3_combout  & (!\Mux34~3_combout  & \ShiftLeft0~106_combout )))

	.dataa(Mux33),
	.datab(Mux34),
	.datac(\ShiftLeft0~97_combout ),
	.datad(\ShiftLeft0~106_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~98_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~98 .lut_mask = 16'hF2F0;
defparam \ShiftLeft0~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N2
cycloneive_lcell_comb \Selector4~2 (
// Equation(s):
// \Selector4~2_combout  = (\Selector4~1_combout  & (((\ShiftLeft0~98_combout )) # (!\Selector5~1_combout ))) # (!\Selector4~1_combout  & (\Selector5~1_combout  & (\ShiftLeft0~96_combout )))

	.dataa(\Selector4~1_combout ),
	.datab(\Selector5~1_combout ),
	.datac(\ShiftLeft0~96_combout ),
	.datad(\ShiftLeft0~98_combout ),
	.cin(gnd),
	.combout(\Selector4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~2 .lut_mask = 16'hEA62;
defparam \Selector4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y40_N16
cycloneive_lcell_comb \Selector4~3 (
// Equation(s):
// \Selector4~3_combout  = (!\ShiftRight0~61_combout  & (\Selector0~7_combout  & \Selector4~2_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~61_combout ),
	.datac(\Selector0~7_combout ),
	.datad(\Selector4~2_combout ),
	.cin(gnd),
	.combout(\Selector4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~3 .lut_mask = 16'h3000;
defparam \Selector4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N30
cycloneive_lcell_comb \Selector4~7 (
// Equation(s):
// \Selector4~7_combout  = (\Mux9~1_combout  & (((\Selector0~8_combout )))) # (!\Mux9~1_combout  & (!Mux4 & ((\Selector0~11_combout ))))

	.dataa(Mux4),
	.datab(\Selector0~8_combout ),
	.datac(\Selector0~11_combout ),
	.datad(Mux92),
	.cin(gnd),
	.combout(\Selector4~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~7 .lut_mask = 16'hCC50;
defparam \Selector4~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N24
cycloneive_lcell_comb \Selector4~6 (
// Equation(s):
// \Selector4~6_combout  = (\Selector0~10_combout  & (Mux4 $ (((\Mux5~1_combout ) # (\Mux9~0_combout )))))

	.dataa(Mux5),
	.datab(\Selector0~10_combout ),
	.datac(Mux4),
	.datad(Mux9),
	.cin(gnd),
	.combout(\Selector4~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~6 .lut_mask = 16'h0C48;
defparam \Selector4~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N0
cycloneive_lcell_comb \Selector4~5 (
// Equation(s):
// \Selector4~5_combout  = (Mux4 & ((\Selector0~8_combout ) # ((\Mux9~1_combout  & \Selector0~9_combout ))))

	.dataa(Mux92),
	.datab(\Selector0~8_combout ),
	.datac(\Selector0~9_combout ),
	.datad(Mux4),
	.cin(gnd),
	.combout(\Selector4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~5 .lut_mask = 16'hEC00;
defparam \Selector4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N10
cycloneive_lcell_comb \Selector4~4 (
// Equation(s):
// \Selector4~4_combout  = (\Selector0~13_combout  & ((\Add0~54_combout ) # ((\Selector0~12_combout  & \Add1~54_combout )))) # (!\Selector0~13_combout  & (\Selector0~12_combout  & (\Add1~54_combout )))

	.dataa(\Selector0~13_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Add1~54_combout ),
	.datad(\Add0~54_combout ),
	.cin(gnd),
	.combout(\Selector4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~4 .lut_mask = 16'hEAC0;
defparam \Selector4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N12
cycloneive_lcell_comb \Selector4~8 (
// Equation(s):
// \Selector4~8_combout  = (\Selector4~7_combout ) # ((\Selector4~6_combout ) # ((\Selector4~5_combout ) # (\Selector4~4_combout )))

	.dataa(\Selector4~7_combout ),
	.datab(\Selector4~6_combout ),
	.datac(\Selector4~5_combout ),
	.datad(\Selector4~4_combout ),
	.cin(gnd),
	.combout(\Selector4~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector4~8 .lut_mask = 16'hFFFE;
defparam \Selector4~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N26
cycloneive_lcell_comb \ShiftLeft0~115 (
// Equation(s):
// \ShiftLeft0~115_combout  = (\Mux35~2_combout  & (((\ShiftLeft0~62_combout )))) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & ((\ShiftLeft0~62_combout ))) # (!\Mux35~3_combout  & (\ShiftLeft0~63_combout ))))

	.dataa(Mux35),
	.datab(Mux351),
	.datac(\ShiftLeft0~63_combout ),
	.datad(\ShiftLeft0~62_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~115_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~115 .lut_mask = 16'hFE10;
defparam \ShiftLeft0~115 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N6
cycloneive_lcell_comb \ShiftLeft0~114 (
// Equation(s):
// \ShiftLeft0~114_combout  = (\Mux35~2_combout  & (((\ShiftLeft0~59_combout )))) # (!\Mux35~2_combout  & ((\Mux35~3_combout  & ((\ShiftLeft0~59_combout ))) # (!\Mux35~3_combout  & (\ShiftLeft0~61_combout ))))

	.dataa(Mux35),
	.datab(\ShiftLeft0~61_combout ),
	.datac(Mux351),
	.datad(\ShiftLeft0~59_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~114_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~114 .lut_mask = 16'hFE04;
defparam \ShiftLeft0~114 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N12
cycloneive_lcell_comb \Selector10~0 (
// Equation(s):
// \Selector10~0_combout  = (\Mux34~3_combout  & ((\ShiftLeft0~114_combout ))) # (!\Mux34~3_combout  & (\ShiftLeft0~115_combout ))

	.dataa(Mux34),
	.datab(gnd),
	.datac(\ShiftLeft0~115_combout ),
	.datad(\ShiftLeft0~114_combout ),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~0 .lut_mask = 16'hFA50;
defparam \Selector10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N0
cycloneive_lcell_comb \Selector10~1 (
// Equation(s):
// \Selector10~1_combout  = (!cuifaluOp_0 & (\Selector16~1_combout  & \ShiftLeft0~71_combout ))

	.dataa(cuifaluOp_0),
	.datab(gnd),
	.datac(\Selector16~1_combout ),
	.datad(\ShiftLeft0~71_combout ),
	.cin(gnd),
	.combout(\Selector10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~1 .lut_mask = 16'h5000;
defparam \Selector10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N4
cycloneive_lcell_comb \Selector10~5 (
// Equation(s):
// \Selector10~5_combout  = (\Selector0~15_combout ) # ((\Selector0~16_combout  & ((\Mux15~0_combout ) # (\Mux5~1_combout ))))

	.dataa(Mux15),
	.datab(Mux5),
	.datac(\Selector0~15_combout ),
	.datad(\Selector0~16_combout ),
	.cin(gnd),
	.combout(\Selector10~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~5 .lut_mask = 16'hFEF0;
defparam \Selector10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N0
cycloneive_lcell_comb \Selector10~3 (
// Equation(s):
// \Selector10~3_combout  = (\Mux15~1_combout  & (((\Selector0~15_combout )))) # (!\Mux15~1_combout  & (\Selector0~18_combout  & ((!Mux10))))

	.dataa(\Selector0~18_combout ),
	.datab(\Selector0~15_combout ),
	.datac(Mux151),
	.datad(Mux101),
	.cin(gnd),
	.combout(\Selector10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~3 .lut_mask = 16'hC0CA;
defparam \Selector10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N2
cycloneive_lcell_comb \Selector10~4 (
// Equation(s):
// \Selector10~4_combout  = (\Selector10~3_combout ) # ((\Selector0~17_combout  & (Mux10 $ (\Mux15~1_combout ))))

	.dataa(Mux101),
	.datab(\Selector0~17_combout ),
	.datac(Mux151),
	.datad(\Selector10~3_combout ),
	.cin(gnd),
	.combout(\Selector10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~4 .lut_mask = 16'hFF48;
defparam \Selector10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N18
cycloneive_lcell_comb \Selector10~6 (
// Equation(s):
// \Selector10~6_combout  = (\Selector10~4_combout ) # ((Mux10 & \Selector10~5_combout ))

	.dataa(Mux101),
	.datab(gnd),
	.datac(\Selector10~5_combout ),
	.datad(\Selector10~4_combout ),
	.cin(gnd),
	.combout(\Selector10~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~6 .lut_mask = 16'hFFA0;
defparam \Selector10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N26
cycloneive_lcell_comb \Selector10~2 (
// Equation(s):
// \Selector10~2_combout  = (\Selector0~19_combout  & ((\Add1~42_combout ) # ((\Selector0~20_combout  & \Add0~42_combout )))) # (!\Selector0~19_combout  & (\Selector0~20_combout  & (\Add0~42_combout )))

	.dataa(\Selector0~19_combout ),
	.datab(\Selector0~20_combout ),
	.datac(\Add0~42_combout ),
	.datad(\Add1~42_combout ),
	.cin(gnd),
	.combout(\Selector10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~2 .lut_mask = 16'hEAC0;
defparam \Selector10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N6
cycloneive_lcell_comb \Selector10~7 (
// Equation(s):
// \Selector10~7_combout  = (\Selector10~6_combout ) # ((\Selector10~2_combout ) # ((\ShiftRight0~116_combout  & \Selector8~0_combout )))

	.dataa(\ShiftRight0~116_combout ),
	.datab(\Selector10~6_combout ),
	.datac(\Selector8~0_combout ),
	.datad(\Selector10~2_combout ),
	.cin(gnd),
	.combout(\Selector10~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~7 .lut_mask = 16'hFFEC;
defparam \Selector10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N20
cycloneive_lcell_comb \Selector10~8 (
// Equation(s):
// \Selector10~8_combout  = (\Selector10~1_combout ) # ((\Selector10~7_combout ) # ((\Selector10~0_combout  & \Selector0~27_combout )))

	.dataa(\Selector10~0_combout ),
	.datab(\Selector10~1_combout ),
	.datac(\Selector0~27_combout ),
	.datad(\Selector10~7_combout ),
	.cin(gnd),
	.combout(\Selector10~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector10~8 .lut_mask = 16'hFFEC;
defparam \Selector10~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N14
cycloneive_lcell_comb \ShiftLeft0~100 (
// Equation(s):
// \ShiftLeft0~100_combout  = (!\Selector0~30_combout  & ((\Mux36~4_combout  & (Mux31)) # (!\Mux36~4_combout  & ((Mux30)))))

	.dataa(Mux36),
	.datab(Mux311),
	.datac(\Selector0~30_combout ),
	.datad(Mux301),
	.cin(gnd),
	.combout(\ShiftLeft0~100_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~100 .lut_mask = 16'h0D08;
defparam \ShiftLeft0~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N28
cycloneive_lcell_comb \ShiftLeft0~101 (
// Equation(s):
// \ShiftLeft0~101_combout  = (\Mux33~3_combout  & (((\ShiftLeft0~100_combout )))) # (!\Mux33~3_combout  & (!\Mux34~3_combout  & ((\ShiftLeft0~114_combout ))))

	.dataa(Mux34),
	.datab(\ShiftLeft0~100_combout ),
	.datac(Mux33),
	.datad(\ShiftLeft0~114_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~101_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~101 .lut_mask = 16'hC5C0;
defparam \ShiftLeft0~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N18
cycloneive_lcell_comb \ShiftLeft0~102 (
// Equation(s):
// \ShiftLeft0~102_combout  = (\ShiftLeft0~101_combout ) # ((\Mux34~3_combout  & (\ShiftLeft0~113_combout  & !\Mux33~3_combout )))

	.dataa(Mux34),
	.datab(\ShiftLeft0~113_combout ),
	.datac(Mux33),
	.datad(\ShiftLeft0~101_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~102_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~102 .lut_mask = 16'hFF08;
defparam \ShiftLeft0~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N8
cycloneive_lcell_comb \Selector6~0 (
// Equation(s):
// \Selector6~0_combout  = (\Selector5~1_combout  & (((\Selector5~0_combout )))) # (!\Selector5~1_combout  & ((\Selector5~0_combout  & ((\ShiftLeft0~118_combout ))) # (!\Selector5~0_combout  & (\ShiftLeft0~116_combout ))))

	.dataa(\Selector5~1_combout ),
	.datab(\ShiftLeft0~116_combout ),
	.datac(\ShiftLeft0~118_combout ),
	.datad(\Selector5~0_combout ),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~0 .lut_mask = 16'hFA44;
defparam \Selector6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N10
cycloneive_lcell_comb \ShiftLeft0~99 (
// Equation(s):
// \ShiftLeft0~99_combout  = (\Mux34~3_combout  & (\ShiftLeft0~115_combout )) # (!\Mux34~3_combout  & ((\ShiftLeft0~117_combout )))

	.dataa(Mux34),
	.datab(gnd),
	.datac(\ShiftLeft0~115_combout ),
	.datad(\ShiftLeft0~117_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~99_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~99 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N4
cycloneive_lcell_comb \Selector6~1 (
// Equation(s):
// \Selector6~1_combout  = (\Selector5~1_combout  & ((\Selector6~0_combout  & (\ShiftLeft0~102_combout )) # (!\Selector6~0_combout  & ((\ShiftLeft0~99_combout ))))) # (!\Selector5~1_combout  & (((\Selector6~0_combout ))))

	.dataa(\Selector5~1_combout ),
	.datab(\ShiftLeft0~102_combout ),
	.datac(\Selector6~0_combout ),
	.datad(\ShiftLeft0~99_combout ),
	.cin(gnd),
	.combout(\Selector6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~1 .lut_mask = 16'hDAD0;
defparam \Selector6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N2
cycloneive_lcell_comb \Selector6~2 (
// Equation(s):
// \Selector6~2_combout  = (\Selector0~7_combout  & (!\ShiftRight0~61_combout  & \Selector6~1_combout ))

	.dataa(\Selector0~7_combout ),
	.datab(gnd),
	.datac(\ShiftRight0~61_combout ),
	.datad(\Selector6~1_combout ),
	.cin(gnd),
	.combout(\Selector6~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~2 .lut_mask = 16'h0A00;
defparam \Selector6~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N10
cycloneive_lcell_comb \Selector6~6 (
// Equation(s):
// \Selector6~6_combout  = (\Selector0~8_combout ) # ((\Selector0~9_combout  & ((\Mux5~1_combout ) # (\Mux11~0_combout ))))

	.dataa(Mux5),
	.datab(\Selector0~8_combout ),
	.datac(\Selector0~9_combout ),
	.datad(Mux11),
	.cin(gnd),
	.combout(\Selector6~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~6 .lut_mask = 16'hFCEC;
defparam \Selector6~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N22
cycloneive_lcell_comb \Selector6~4 (
// Equation(s):
// \Selector6~4_combout  = (\Mux11~1_combout  & (\Selector0~8_combout )) # (!\Mux11~1_combout  & (((!Mux6 & \Selector0~11_combout ))))

	.dataa(Mux112),
	.datab(\Selector0~8_combout ),
	.datac(Mux61),
	.datad(\Selector0~11_combout ),
	.cin(gnd),
	.combout(\Selector6~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~4 .lut_mask = 16'h8D88;
defparam \Selector6~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N8
cycloneive_lcell_comb \Selector6~5 (
// Equation(s):
// \Selector6~5_combout  = (\Selector6~4_combout ) # ((\Selector0~10_combout  & (\Mux11~1_combout  $ (Mux6))))

	.dataa(Mux112),
	.datab(Mux61),
	.datac(\Selector6~4_combout ),
	.datad(\Selector0~10_combout ),
	.cin(gnd),
	.combout(\Selector6~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~5 .lut_mask = 16'hF6F0;
defparam \Selector6~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N20
cycloneive_lcell_comb \Selector6~3 (
// Equation(s):
// \Selector6~3_combout  = (\Selector0~12_combout  & ((\Add1~50_combout ) # ((\Selector0~13_combout  & \Add0~50_combout )))) # (!\Selector0~12_combout  & (\Selector0~13_combout  & ((\Add0~50_combout ))))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector0~13_combout ),
	.datac(\Add1~50_combout ),
	.datad(\Add0~50_combout ),
	.cin(gnd),
	.combout(\Selector6~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~3 .lut_mask = 16'hECA0;
defparam \Selector6~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N16
cycloneive_lcell_comb \Selector6~7 (
// Equation(s):
// \Selector6~7_combout  = (\Selector6~5_combout ) # ((\Selector6~3_combout ) # ((\Selector6~6_combout  & Mux6)))

	.dataa(\Selector6~6_combout ),
	.datab(Mux61),
	.datac(\Selector6~5_combout ),
	.datad(\Selector6~3_combout ),
	.cin(gnd),
	.combout(\Selector6~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector6~7 .lut_mask = 16'hFFF8;
defparam \Selector6~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N24
cycloneive_lcell_comb \Selector7~5 (
// Equation(s):
// \Selector7~5_combout  = (\Mux12~1_combout  & (((\Selector0~8_combout )))) # (!\Mux12~1_combout  & (!Mux7 & (\Selector0~11_combout )))

	.dataa(Mux12),
	.datab(Mux71),
	.datac(\Selector0~11_combout ),
	.datad(\Selector0~8_combout ),
	.cin(gnd),
	.combout(\Selector7~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~5 .lut_mask = 16'hBA10;
defparam \Selector7~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N22
cycloneive_lcell_comb \Selector7~6 (
// Equation(s):
// \Selector7~6_combout  = (\Selector7~5_combout ) # ((\Selector0~10_combout  & (Mux7 $ (\Mux12~1_combout ))))

	.dataa(\Selector0~10_combout ),
	.datab(Mux71),
	.datac(Mux12),
	.datad(\Selector7~5_combout ),
	.cin(gnd),
	.combout(\Selector7~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~6 .lut_mask = 16'hFF28;
defparam \Selector7~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N4
cycloneive_lcell_comb \Selector7~4 (
// Equation(s):
// \Selector7~4_combout  = (Mux7 & ((\Selector0~8_combout ) # ((\Mux12~1_combout  & \Selector0~9_combout ))))

	.dataa(\Selector0~8_combout ),
	.datab(Mux12),
	.datac(\Selector0~9_combout ),
	.datad(Mux71),
	.cin(gnd),
	.combout(\Selector7~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~4 .lut_mask = 16'hEA00;
defparam \Selector7~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y38_N26
cycloneive_lcell_comb \Selector7~3 (
// Equation(s):
// \Selector7~3_combout  = (\Selector0~12_combout  & ((\Add1~48_combout ) # ((\Selector0~13_combout  & \Add0~48_combout )))) # (!\Selector0~12_combout  & (\Selector0~13_combout  & ((\Add0~48_combout ))))

	.dataa(\Selector0~12_combout ),
	.datab(\Selector0~13_combout ),
	.datac(\Add1~48_combout ),
	.datad(\Add0~48_combout ),
	.cin(gnd),
	.combout(\Selector7~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~3 .lut_mask = 16'hECA0;
defparam \Selector7~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N8
cycloneive_lcell_comb \ShiftLeft0~104 (
// Equation(s):
// \ShiftLeft0~104_combout  = (!\Mux34~3_combout  & ((\Mux33~3_combout  & (\ShiftLeft0~125_combout )) # (!\Mux33~3_combout  & ((\ShiftLeft0~127_combout )))))

	.dataa(Mux34),
	.datab(Mux33),
	.datac(\ShiftLeft0~125_combout ),
	.datad(\ShiftLeft0~127_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~104_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~104 .lut_mask = 16'h5140;
defparam \ShiftLeft0~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N30
cycloneive_lcell_comb \ShiftLeft0~105 (
// Equation(s):
// \ShiftLeft0~105_combout  = (\ShiftLeft0~104_combout ) # ((\Mux34~3_combout  & (!\Mux33~3_combout  & \ShiftLeft0~126_combout )))

	.dataa(Mux34),
	.datab(Mux33),
	.datac(\ShiftLeft0~104_combout ),
	.datad(\ShiftLeft0~126_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~105_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~105 .lut_mask = 16'hF2F0;
defparam \ShiftLeft0~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N12
cycloneive_lcell_comb \ShiftLeft0~103 (
// Equation(s):
// \ShiftLeft0~103_combout  = (\Mux34~3_combout  & ((\ShiftLeft0~128_combout ))) # (!\Mux34~3_combout  & (\ShiftLeft0~130_combout ))

	.dataa(gnd),
	.datab(Mux34),
	.datac(\ShiftLeft0~130_combout ),
	.datad(\ShiftLeft0~128_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~103_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~103 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N18
cycloneive_lcell_comb \Selector7~0 (
// Equation(s):
// \Selector7~0_combout  = (\Selector5~1_combout  & (((\Selector5~0_combout ) # (\ShiftLeft0~103_combout )))) # (!\Selector5~1_combout  & (\ShiftLeft0~129_combout  & (!\Selector5~0_combout )))

	.dataa(\ShiftLeft0~129_combout ),
	.datab(\Selector5~1_combout ),
	.datac(\Selector5~0_combout ),
	.datad(\ShiftLeft0~103_combout ),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~0 .lut_mask = 16'hCEC2;
defparam \Selector7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y42_N24
cycloneive_lcell_comb \Selector7~1 (
// Equation(s):
// \Selector7~1_combout  = (\Selector5~0_combout  & ((\Selector7~0_combout  & ((\ShiftLeft0~105_combout ))) # (!\Selector7~0_combout  & (\ShiftLeft0~131_combout )))) # (!\Selector5~0_combout  & (((\Selector7~0_combout ))))

	.dataa(\Selector5~0_combout ),
	.datab(\ShiftLeft0~131_combout ),
	.datac(\ShiftLeft0~105_combout ),
	.datad(\Selector7~0_combout ),
	.cin(gnd),
	.combout(\Selector7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~1 .lut_mask = 16'hF588;
defparam \Selector7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N10
cycloneive_lcell_comb \Selector7~2 (
// Equation(s):
// \Selector7~2_combout  = (\Selector0~7_combout  & (!\ShiftRight0~61_combout  & \Selector7~1_combout ))

	.dataa(\Selector0~7_combout ),
	.datab(gnd),
	.datac(\ShiftRight0~61_combout ),
	.datad(\Selector7~1_combout ),
	.cin(gnd),
	.combout(\Selector7~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector7~2 .lut_mask = 16'h0A00;
defparam \Selector7~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N8
cycloneive_lcell_comb \Selector11~1 (
// Equation(s):
// \Selector11~1_combout  = (!cuifaluOp_0 & (\ShiftLeft0~93_combout  & \Selector16~1_combout ))

	.dataa(cuifaluOp_0),
	.datab(gnd),
	.datac(\ShiftLeft0~93_combout ),
	.datad(\Selector16~1_combout ),
	.cin(gnd),
	.combout(\Selector11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~1 .lut_mask = 16'h5000;
defparam \Selector11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N30
cycloneive_lcell_comb \Selector11~4 (
// Equation(s):
// \Selector11~4_combout  = (Mux11 & ((\Selector0~15_combout ) # ((\Mux16~1_combout  & \Selector0~16_combout ))))

	.dataa(\Selector0~15_combout ),
	.datab(Mux16),
	.datac(\Selector0~16_combout ),
	.datad(Mux111),
	.cin(gnd),
	.combout(\Selector11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~4 .lut_mask = 16'hEA00;
defparam \Selector11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N18
cycloneive_lcell_comb \ShiftRight0~117 (
// Equation(s):
// \ShiftRight0~117_combout  = (!\Mux33~3_combout  & ((\Mux34~3_combout  & ((\ShiftRight0~138_combout ))) # (!\Mux34~3_combout  & (\ShiftRight0~139_combout ))))

	.dataa(Mux34),
	.datab(Mux33),
	.datac(\ShiftRight0~139_combout ),
	.datad(\ShiftRight0~138_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~117_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~117 .lut_mask = 16'h3210;
defparam \ShiftRight0~117 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N24
cycloneive_lcell_comb \ShiftRight0~118 (
// Equation(s):
// \ShiftRight0~118_combout  = (\ShiftRight0~117_combout ) # ((!\Mux34~3_combout  & (\Mux33~3_combout  & \ShiftRight0~137_combout )))

	.dataa(Mux34),
	.datab(Mux33),
	.datac(\ShiftRight0~137_combout ),
	.datad(\ShiftRight0~117_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~118_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~118 .lut_mask = 16'hFF40;
defparam \ShiftRight0~118 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N6
cycloneive_lcell_comb \Selector11~2 (
// Equation(s):
// \Selector11~2_combout  = (\Selector0~25_combout  & (!\Mux32~4_combout  & (\ShiftRight0~118_combout  & !\ShiftRight0~61_combout )))

	.dataa(\Selector0~25_combout ),
	.datab(Mux32),
	.datac(\ShiftRight0~118_combout ),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\Selector11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~2 .lut_mask = 16'h0020;
defparam \Selector11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N20
cycloneive_lcell_comb \Selector11~3 (
// Equation(s):
// \Selector11~3_combout  = (\Selector0~20_combout  & ((\Add0~40_combout ) # ((\Selector0~19_combout  & \Add1~40_combout )))) # (!\Selector0~20_combout  & (\Selector0~19_combout  & (\Add1~40_combout )))

	.dataa(\Selector0~20_combout ),
	.datab(\Selector0~19_combout ),
	.datac(\Add1~40_combout ),
	.datad(\Add0~40_combout ),
	.cin(gnd),
	.combout(\Selector11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~3 .lut_mask = 16'hEAC0;
defparam \Selector11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N16
cycloneive_lcell_comb \Selector11~7 (
// Equation(s):
// \Selector11~7_combout  = (\Selector11~6_combout ) # ((\Selector11~4_combout ) # ((\Selector11~2_combout ) # (\Selector11~3_combout )))

	.dataa(\Selector11~6_combout ),
	.datab(\Selector11~4_combout ),
	.datac(\Selector11~2_combout ),
	.datad(\Selector11~3_combout ),
	.cin(gnd),
	.combout(\Selector11~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~7 .lut_mask = 16'hFFFE;
defparam \Selector11~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N18
cycloneive_lcell_comb \Selector11~8 (
// Equation(s):
// \Selector11~8_combout  = (\Selector11~1_combout ) # ((\Selector11~7_combout ) # ((\Selector11~0_combout  & \Selector0~27_combout )))

	.dataa(\Selector11~0_combout ),
	.datab(\Selector11~1_combout ),
	.datac(\Selector0~27_combout ),
	.datad(\Selector11~7_combout ),
	.cin(gnd),
	.combout(\Selector11~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector11~8 .lut_mask = 16'hFFEC;
defparam \Selector11~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N2
cycloneive_lcell_comb \Selector24~2 (
// Equation(s):
// \Selector24~2_combout  = (\Add0~14_combout  & ((\Selector0~13_combout ) # ((\Selector0~12_combout  & \Add1~14_combout )))) # (!\Add0~14_combout  & (\Selector0~12_combout  & ((\Add1~14_combout ))))

	.dataa(\Add0~14_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Selector0~13_combout ),
	.datad(\Add1~14_combout ),
	.cin(gnd),
	.combout(\Selector24~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~2 .lut_mask = 16'hECA0;
defparam \Selector24~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N0
cycloneive_lcell_comb \Selector24~3 (
// Equation(s):
// \Selector24~3_combout  = (\Selector24~2_combout ) # ((!\Mux29~1_combout  & (\Selector0~11_combout  & !Mux24)))

	.dataa(Mux29),
	.datab(\Selector0~11_combout ),
	.datac(Mux241),
	.datad(\Selector24~2_combout ),
	.cin(gnd),
	.combout(\Selector24~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~3 .lut_mask = 16'hFF04;
defparam \Selector24~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N6
cycloneive_lcell_comb \Selector24~4 (
// Equation(s):
// \Selector24~4_combout  = (\Selector24~3_combout ) # ((\Selector0~10_combout  & (\Mux29~1_combout  $ (Mux24))))

	.dataa(Mux29),
	.datab(\Selector0~10_combout ),
	.datac(Mux241),
	.datad(\Selector24~3_combout ),
	.cin(gnd),
	.combout(\Selector24~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~4 .lut_mask = 16'hFF48;
defparam \Selector24~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N28
cycloneive_lcell_comb \Selector24~1 (
// Equation(s):
// \Selector24~1_combout  = (\Mux29~1_combout  & ((\Selector0~8_combout ) # ((Mux24 & \Selector0~9_combout )))) # (!\Mux29~1_combout  & (Mux24 & (\Selector0~8_combout )))

	.dataa(Mux29),
	.datab(Mux241),
	.datac(\Selector0~8_combout ),
	.datad(\Selector0~9_combout ),
	.cin(gnd),
	.combout(\Selector24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~1 .lut_mask = 16'hE8E0;
defparam \Selector24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N12
cycloneive_lcell_comb \ShiftRight0~119 (
// Equation(s):
// \ShiftRight0~119_combout  = (\Mux34~3_combout  & ((\ShiftRight0~147_combout ))) # (!\Mux34~3_combout  & (\ShiftRight0~142_combout ))

	.dataa(Mux34),
	.datab(gnd),
	.datac(\ShiftRight0~142_combout ),
	.datad(\ShiftRight0~147_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~119_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~119 .lut_mask = 16'hFA50;
defparam \ShiftRight0~119 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N30
cycloneive_lcell_comb \Selector24~5 (
// Equation(s):
// \Selector24~5_combout  = (\Selector5~0_combout  & ((\Selector5~1_combout ) # ((\ShiftRight0~143_combout )))) # (!\Selector5~0_combout  & (!\Selector5~1_combout  & (\ShiftRight0~141_combout )))

	.dataa(\Selector5~0_combout ),
	.datab(\Selector5~1_combout ),
	.datac(\ShiftRight0~141_combout ),
	.datad(\ShiftRight0~143_combout ),
	.cin(gnd),
	.combout(\Selector24~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~5 .lut_mask = 16'hBA98;
defparam \Selector24~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N14
cycloneive_lcell_comb \ShiftRight0~120 (
// Equation(s):
// \ShiftRight0~120_combout  = (!\Mux34~3_combout  & ((\Mux33~3_combout  & ((\ShiftRight0~144_combout ))) # (!\Mux33~3_combout  & (\ShiftRight0~146_combout ))))

	.dataa(Mux33),
	.datab(Mux34),
	.datac(\ShiftRight0~146_combout ),
	.datad(\ShiftRight0~144_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~120_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~120 .lut_mask = 16'h3210;
defparam \ShiftRight0~120 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N12
cycloneive_lcell_comb \ShiftRight0~121 (
// Equation(s):
// \ShiftRight0~121_combout  = (\ShiftRight0~120_combout ) # ((!\Mux33~3_combout  & (\Mux34~3_combout  & \ShiftRight0~145_combout )))

	.dataa(Mux33),
	.datab(Mux34),
	.datac(\ShiftRight0~120_combout ),
	.datad(\ShiftRight0~145_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~121_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~121 .lut_mask = 16'hF4F0;
defparam \ShiftRight0~121 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N4
cycloneive_lcell_comb \Selector24~6 (
// Equation(s):
// \Selector24~6_combout  = (\Selector5~1_combout  & ((\Selector24~5_combout  & ((\ShiftRight0~121_combout ))) # (!\Selector24~5_combout  & (\ShiftRight0~119_combout )))) # (!\Selector5~1_combout  & (((\Selector24~5_combout ))))

	.dataa(\ShiftRight0~119_combout ),
	.datab(\Selector5~1_combout ),
	.datac(\Selector24~5_combout ),
	.datad(\ShiftRight0~121_combout ),
	.cin(gnd),
	.combout(\Selector24~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector24~6 .lut_mask = 16'hF838;
defparam \Selector24~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N8
cycloneive_lcell_comb \ShiftRight0~124 (
// Equation(s):
// \ShiftRight0~124_combout  = (\Mux33~3_combout  & (\ShiftRight0~123_combout )) # (!\Mux33~3_combout  & (((!\Mux34~3_combout  & \ShiftRight0~152_combout ))))

	.dataa(\ShiftRight0~123_combout ),
	.datab(Mux33),
	.datac(Mux34),
	.datad(\ShiftRight0~152_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~124_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~124 .lut_mask = 16'h8B88;
defparam \ShiftRight0~124 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N26
cycloneive_lcell_comb \ShiftRight0~125 (
// Equation(s):
// \ShiftRight0~125_combout  = (\ShiftRight0~124_combout ) # ((\Mux34~3_combout  & (!\Mux33~3_combout  & \ShiftRight0~151_combout )))

	.dataa(Mux34),
	.datab(Mux33),
	.datac(\ShiftRight0~124_combout ),
	.datad(\ShiftRight0~151_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~125_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~125 .lut_mask = 16'hF2F0;
defparam \ShiftRight0~125 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N26
cycloneive_lcell_comb \ShiftRight0~122 (
// Equation(s):
// \ShiftRight0~122_combout  = (\Mux34~3_combout  & ((\ShiftRight0~153_combout ))) # (!\Mux34~3_combout  & (\ShiftRight0~149_combout ))

	.dataa(Mux34),
	.datab(gnd),
	.datac(\ShiftRight0~149_combout ),
	.datad(\ShiftRight0~153_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~122_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~122 .lut_mask = 16'hFA50;
defparam \ShiftRight0~122 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N6
cycloneive_lcell_comb \Selector25~4 (
// Equation(s):
// \Selector25~4_combout  = (\Selector5~1_combout  & (((\Selector5~0_combout ) # (\ShiftRight0~122_combout )))) # (!\Selector5~1_combout  & (\ShiftRight0~148_combout  & (!\Selector5~0_combout )))

	.dataa(\Selector5~1_combout ),
	.datab(\ShiftRight0~148_combout ),
	.datac(\Selector5~0_combout ),
	.datad(\ShiftRight0~122_combout ),
	.cin(gnd),
	.combout(\Selector25~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~4 .lut_mask = 16'hAEA4;
defparam \Selector25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N0
cycloneive_lcell_comb \Selector25~5 (
// Equation(s):
// \Selector25~5_combout  = (\Selector5~0_combout  & ((\Selector25~4_combout  & (\ShiftRight0~125_combout )) # (!\Selector25~4_combout  & ((\ShiftRight0~150_combout ))))) # (!\Selector5~0_combout  & (((\Selector25~4_combout ))))

	.dataa(\Selector5~0_combout ),
	.datab(\ShiftRight0~125_combout ),
	.datac(\ShiftRight0~150_combout ),
	.datad(\Selector25~4_combout ),
	.cin(gnd),
	.combout(\Selector25~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~5 .lut_mask = 16'hDDA0;
defparam \Selector25~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N14
cycloneive_lcell_comb \Selector25~0 (
// Equation(s):
// \Selector25~0_combout  = (Mux25 & ((\Selector0~8_combout ) # ((\Mux30~1_combout  & \Selector0~9_combout )))) # (!Mux25 & (\Mux30~1_combout  & (\Selector0~8_combout )))

	.dataa(Mux251),
	.datab(Mux30),
	.datac(\Selector0~8_combout ),
	.datad(\Selector0~9_combout ),
	.cin(gnd),
	.combout(\Selector25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~0 .lut_mask = 16'hE8E0;
defparam \Selector25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N0
cycloneive_lcell_comb \Selector25~1 (
// Equation(s):
// \Selector25~1_combout  = (\Selector0~13_combout  & ((\Add0~12_combout ) # ((\Selector0~12_combout  & \Add1~12_combout )))) # (!\Selector0~13_combout  & (\Selector0~12_combout  & ((\Add1~12_combout ))))

	.dataa(\Selector0~13_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Add0~12_combout ),
	.datad(\Add1~12_combout ),
	.cin(gnd),
	.combout(\Selector25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~1 .lut_mask = 16'hECA0;
defparam \Selector25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N2
cycloneive_lcell_comb \Selector25~2 (
// Equation(s):
// \Selector25~2_combout  = (\Selector25~1_combout ) # ((!Mux25 & (\Selector0~11_combout  & !\Mux30~1_combout )))

	.dataa(Mux251),
	.datab(\Selector0~11_combout ),
	.datac(Mux30),
	.datad(\Selector25~1_combout ),
	.cin(gnd),
	.combout(\Selector25~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~2 .lut_mask = 16'hFF04;
defparam \Selector25~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N4
cycloneive_lcell_comb \Selector25~3 (
// Equation(s):
// \Selector25~3_combout  = (\Selector25~2_combout ) # ((\Selector0~10_combout  & (Mux25 $ (\Mux30~1_combout ))))

	.dataa(Mux251),
	.datab(\Selector0~10_combout ),
	.datac(Mux30),
	.datad(\Selector25~2_combout ),
	.cin(gnd),
	.combout(\Selector25~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector25~3 .lut_mask = 16'hFF48;
defparam \Selector25~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N4
cycloneive_lcell_comb \Selector13~3 (
// Equation(s):
// \Selector13~3_combout  = (\Selector0~17_combout  & (Mux13 $ (((\Mux5~1_combout ) # (\Mux18~0_combout )))))

	.dataa(\Selector0~17_combout ),
	.datab(Mux5),
	.datac(Mux131),
	.datad(Mux18),
	.cin(gnd),
	.combout(\Selector13~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~3 .lut_mask = 16'h0A28;
defparam \Selector13~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N14
cycloneive_lcell_comb \Selector13~2 (
// Equation(s):
// \Selector13~2_combout  = (Mux13 & ((\Selector0~15_combout ) # ((\Selector0~16_combout  & \Mux18~1_combout ))))

	.dataa(\Selector0~16_combout ),
	.datab(\Selector0~15_combout ),
	.datac(Mux131),
	.datad(Mux182),
	.cin(gnd),
	.combout(\Selector13~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~2 .lut_mask = 16'hE0C0;
defparam \Selector13~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N28
cycloneive_lcell_comb \Selector13~1 (
// Equation(s):
// \Selector13~1_combout  = (\Add1~36_combout  & ((\Selector0~19_combout ) # ((\Selector0~20_combout  & \Add0~36_combout )))) # (!\Add1~36_combout  & (((\Selector0~20_combout  & \Add0~36_combout ))))

	.dataa(\Add1~36_combout ),
	.datab(\Selector0~19_combout ),
	.datac(\Selector0~20_combout ),
	.datad(\Add0~36_combout ),
	.cin(gnd),
	.combout(\Selector13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~1 .lut_mask = 16'hF888;
defparam \Selector13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N24
cycloneive_lcell_comb \Selector13~5 (
// Equation(s):
// \Selector13~5_combout  = (\Selector13~4_combout ) # ((\Selector13~3_combout ) # ((\Selector13~2_combout ) # (\Selector13~1_combout )))

	.dataa(\Selector13~4_combout ),
	.datab(\Selector13~3_combout ),
	.datac(\Selector13~2_combout ),
	.datad(\Selector13~1_combout ),
	.cin(gnd),
	.combout(\Selector13~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~5 .lut_mask = 16'hFFFE;
defparam \Selector13~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N10
cycloneive_lcell_comb \ShiftLeft0~124 (
// Equation(s):
// \ShiftLeft0~124_combout  = (\Mux35~3_combout  & (((\ShiftLeft0~85_combout )))) # (!\Mux35~3_combout  & ((\Mux35~2_combout  & ((\ShiftLeft0~85_combout ))) # (!\Mux35~2_combout  & (\ShiftLeft0~86_combout ))))

	.dataa(Mux351),
	.datab(\ShiftLeft0~86_combout ),
	.datac(Mux35),
	.datad(\ShiftLeft0~85_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~124_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~124 .lut_mask = 16'hFE04;
defparam \ShiftLeft0~124 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N14
cycloneive_lcell_comb \Selector13~0 (
// Equation(s):
// \Selector13~0_combout  = (\Selector0~27_combout  & ((\Mux34~3_combout  & (\ShiftLeft0~123_combout )) # (!\Mux34~3_combout  & ((\ShiftLeft0~124_combout )))))

	.dataa(Mux34),
	.datab(\ShiftLeft0~123_combout ),
	.datac(\Selector0~27_combout ),
	.datad(\ShiftLeft0~124_combout ),
	.cin(gnd),
	.combout(\Selector13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~0 .lut_mask = 16'hD080;
defparam \Selector13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N24
cycloneive_lcell_comb \Selector13~6 (
// Equation(s):
// \Selector13~6_combout  = (\Selector13~5_combout ) # ((\Selector13~0_combout ) # ((\Selector8~0_combout  & \ShiftRight0~114_combout )))

	.dataa(\Selector8~0_combout ),
	.datab(\ShiftRight0~114_combout ),
	.datac(\Selector13~5_combout ),
	.datad(\Selector13~0_combout ),
	.cin(gnd),
	.combout(\Selector13~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~6 .lut_mask = 16'hFFF8;
defparam \Selector13~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N26
cycloneive_lcell_comb \Selector13~7 (
// Equation(s):
// \Selector13~7_combout  = (\Selector13~6_combout ) # ((\Selector16~1_combout  & (!cuifaluOp_0 & \ShiftLeft0~80_combout )))

	.dataa(\Selector16~1_combout ),
	.datab(cuifaluOp_0),
	.datac(\ShiftLeft0~80_combout ),
	.datad(\Selector13~6_combout ),
	.cin(gnd),
	.combout(\Selector13~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector13~7 .lut_mask = 16'hFF20;
defparam \Selector13~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N28
cycloneive_lcell_comb \Selector12~2 (
// Equation(s):
// \Selector12~2_combout  = (Mux12 & ((\Selector0~15_combout ) # ((\Selector0~16_combout  & \Mux17~1_combout ))))

	.dataa(\Selector0~16_combout ),
	.datab(Mux172),
	.datac(Mux121),
	.datad(\Selector0~15_combout ),
	.cin(gnd),
	.combout(\Selector12~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~2 .lut_mask = 16'hF080;
defparam \Selector12~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N4
cycloneive_lcell_comb \Selector12~4 (
// Equation(s):
// \Selector12~4_combout  = (\Mux17~1_combout  & (\Selector0~15_combout )) # (!\Mux17~1_combout  & (((!Mux12 & \Selector0~18_combout ))))

	.dataa(\Selector0~15_combout ),
	.datab(Mux121),
	.datac(\Selector0~18_combout ),
	.datad(Mux172),
	.cin(gnd),
	.combout(\Selector12~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~4 .lut_mask = 16'hAA30;
defparam \Selector12~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N2
cycloneive_lcell_comb \Selector12~1 (
// Equation(s):
// \Selector12~1_combout  = (\Selector0~19_combout  & ((\Add1~38_combout ) # ((\Selector0~20_combout  & \Add0~38_combout )))) # (!\Selector0~19_combout  & (\Selector0~20_combout  & (\Add0~38_combout )))

	.dataa(\Selector0~19_combout ),
	.datab(\Selector0~20_combout ),
	.datac(\Add0~38_combout ),
	.datad(\Add1~38_combout ),
	.cin(gnd),
	.combout(\Selector12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~1 .lut_mask = 16'hEAC0;
defparam \Selector12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N14
cycloneive_lcell_comb \Selector12~5 (
// Equation(s):
// \Selector12~5_combout  = (\Selector12~3_combout ) # ((\Selector12~2_combout ) # ((\Selector12~4_combout ) # (\Selector12~1_combout )))

	.dataa(\Selector12~3_combout ),
	.datab(\Selector12~2_combout ),
	.datac(\Selector12~4_combout ),
	.datad(\Selector12~1_combout ),
	.cin(gnd),
	.combout(\Selector12~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~5 .lut_mask = 16'hFFFE;
defparam \Selector12~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N20
cycloneive_lcell_comb \Selector12~0 (
// Equation(s):
// \Selector12~0_combout  = (\Selector0~27_combout  & ((\Mux34~3_combout  & ((\ShiftLeft0~109_combout ))) # (!\Mux34~3_combout  & (\ShiftLeft0~110_combout ))))

	.dataa(\ShiftLeft0~110_combout ),
	.datab(\ShiftLeft0~109_combout ),
	.datac(\Selector0~27_combout ),
	.datad(Mux34),
	.cin(gnd),
	.combout(\Selector12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~0 .lut_mask = 16'hC0A0;
defparam \Selector12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N24
cycloneive_lcell_comb \Selector12~6 (
// Equation(s):
// \Selector12~6_combout  = (\Selector12~5_combout ) # ((\Selector12~0_combout ) # ((\ShiftRight0~111_combout  & \Selector8~0_combout )))

	.dataa(\ShiftRight0~111_combout ),
	.datab(\Selector8~0_combout ),
	.datac(\Selector12~5_combout ),
	.datad(\Selector12~0_combout ),
	.cin(gnd),
	.combout(\Selector12~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~6 .lut_mask = 16'hFFF8;
defparam \Selector12~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N14
cycloneive_lcell_comb \Selector12~7 (
// Equation(s):
// \Selector12~7_combout  = (\Selector12~6_combout ) # ((\Selector16~1_combout  & (\ShiftLeft0~96_combout  & !cuifaluOp_0)))

	.dataa(\Selector16~1_combout ),
	.datab(\ShiftLeft0~96_combout ),
	.datac(cuifaluOp_0),
	.datad(\Selector12~6_combout ),
	.cin(gnd),
	.combout(\Selector12~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector12~7 .lut_mask = 16'hFF08;
defparam \Selector12~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N8
cycloneive_lcell_comb \Selector26~0 (
// Equation(s):
// \Selector26~0_combout  = (\Selector0~8_combout  & (((\Mux31~1_combout ) # (Mux26)))) # (!\Selector0~8_combout  & (\Selector0~9_combout  & (\Mux31~1_combout  & Mux26)))

	.dataa(\Selector0~8_combout ),
	.datab(\Selector0~9_combout ),
	.datac(Mux31),
	.datad(Mux261),
	.cin(gnd),
	.combout(\Selector26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~0 .lut_mask = 16'hEAA0;
defparam \Selector26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N28
cycloneive_lcell_comb \Selector26~2 (
// Equation(s):
// \Selector26~2_combout  = (\Selector26~1_combout ) # ((\Selector0~11_combout  & (!\Mux31~1_combout  & !Mux26)))

	.dataa(\Selector26~1_combout ),
	.datab(\Selector0~11_combout ),
	.datac(Mux31),
	.datad(Mux261),
	.cin(gnd),
	.combout(\Selector26~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~2 .lut_mask = 16'hAAAE;
defparam \Selector26~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N26
cycloneive_lcell_comb \Selector26~3 (
// Equation(s):
// \Selector26~3_combout  = (\Selector26~2_combout ) # ((\Selector0~10_combout  & (Mux26 $ (\Mux31~1_combout ))))

	.dataa(Mux261),
	.datab(\Selector0~10_combout ),
	.datac(Mux31),
	.datad(\Selector26~2_combout ),
	.cin(gnd),
	.combout(\Selector26~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~3 .lut_mask = 16'hFF48;
defparam \Selector26~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N16
cycloneive_lcell_comb \Selector26~4 (
// Equation(s):
// \Selector26~4_combout  = (\Selector5~1_combout  & (\Selector5~0_combout )) # (!\Selector5~1_combout  & ((\Selector5~0_combout  & (\ShiftRight0~130_combout )) # (!\Selector5~0_combout  & ((\ShiftRight0~128_combout )))))

	.dataa(\Selector5~1_combout ),
	.datab(\Selector5~0_combout ),
	.datac(\ShiftRight0~130_combout ),
	.datad(\ShiftRight0~128_combout ),
	.cin(gnd),
	.combout(\Selector26~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~4 .lut_mask = 16'hD9C8;
defparam \Selector26~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N14
cycloneive_lcell_comb \ShiftRight0~126 (
// Equation(s):
// \ShiftRight0~126_combout  = (\Mux34~3_combout  & ((\ShiftRight0~133_combout ))) # (!\Mux34~3_combout  & (\ShiftRight0~129_combout ))

	.dataa(Mux34),
	.datab(gnd),
	.datac(\ShiftRight0~129_combout ),
	.datad(\ShiftRight0~133_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~126_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~126 .lut_mask = 16'hFA50;
defparam \ShiftRight0~126 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N26
cycloneive_lcell_comb \ShiftRight0~115 (
// Equation(s):
// \ShiftRight0~115_combout  = (!\Mux33~3_combout  & ((\Mux34~3_combout  & (\ShiftRight0~131_combout )) # (!\Mux34~3_combout  & ((\ShiftRight0~132_combout )))))

	.dataa(Mux33),
	.datab(Mux34),
	.datac(\ShiftRight0~131_combout ),
	.datad(\ShiftRight0~132_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~115_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~115 .lut_mask = 16'h5140;
defparam \ShiftRight0~115 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N0
cycloneive_lcell_comb \ShiftRight0~116 (
// Equation(s):
// \ShiftRight0~116_combout  = (\ShiftRight0~115_combout ) # ((\Mux33~3_combout  & (!\Mux34~3_combout  & \ShiftRight0~75_combout )))

	.dataa(Mux33),
	.datab(Mux34),
	.datac(\ShiftRight0~115_combout ),
	.datad(\ShiftRight0~75_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~116_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~116 .lut_mask = 16'hF2F0;
defparam \ShiftRight0~116 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N22
cycloneive_lcell_comb \Selector26~5 (
// Equation(s):
// \Selector26~5_combout  = (\Selector5~1_combout  & ((\Selector26~4_combout  & ((\ShiftRight0~116_combout ))) # (!\Selector26~4_combout  & (\ShiftRight0~126_combout )))) # (!\Selector5~1_combout  & (\Selector26~4_combout ))

	.dataa(\Selector5~1_combout ),
	.datab(\Selector26~4_combout ),
	.datac(\ShiftRight0~126_combout ),
	.datad(\ShiftRight0~116_combout ),
	.cin(gnd),
	.combout(\Selector26~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector26~5 .lut_mask = 16'hEC64;
defparam \Selector26~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N10
cycloneive_lcell_comb \Selector27~0 (
// Equation(s):
// \Selector27~0_combout  = (\Selector0~8_combout ) # ((\Selector0~9_combout  & Mux27))

	.dataa(gnd),
	.datab(\Selector0~9_combout ),
	.datac(\Selector0~8_combout ),
	.datad(Mux271),
	.cin(gnd),
	.combout(\Selector27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~0 .lut_mask = 16'hFCF0;
defparam \Selector27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N26
cycloneive_lcell_comb \Selector27~1 (
// Equation(s):
// \Selector27~1_combout  = (\Mux32~4_combout  & ((\Selector27~0_combout ) # ((\Selector0~10_combout  & !Mux27)))) # (!\Mux32~4_combout  & (\Selector0~10_combout  & ((Mux27))))

	.dataa(Mux32),
	.datab(\Selector0~10_combout ),
	.datac(\Selector27~0_combout ),
	.datad(Mux271),
	.cin(gnd),
	.combout(\Selector27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~1 .lut_mask = 16'hE4A8;
defparam \Selector27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N8
cycloneive_lcell_comb \Selector27~2 (
// Equation(s):
// \Selector27~2_combout  = (!\Mux32~4_combout  & (\Selector0~11_combout  & !Mux27))

	.dataa(gnd),
	.datab(Mux32),
	.datac(\Selector0~11_combout ),
	.datad(Mux271),
	.cin(gnd),
	.combout(\Selector27~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~2 .lut_mask = 16'h0030;
defparam \Selector27~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N2
cycloneive_lcell_comb \Selector27~3 (
// Equation(s):
// \Selector27~3_combout  = (\Selector0~13_combout  & ((\Add0~8_combout ) # ((\Selector0~12_combout  & \Add1~8_combout )))) # (!\Selector0~13_combout  & (\Selector0~12_combout  & ((\Add1~8_combout ))))

	.dataa(\Selector0~13_combout ),
	.datab(\Selector0~12_combout ),
	.datac(\Add0~8_combout ),
	.datad(\Add1~8_combout ),
	.cin(gnd),
	.combout(\Selector27~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~3 .lut_mask = 16'hECA0;
defparam \Selector27~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N16
cycloneive_lcell_comb \Selector27~4 (
// Equation(s):
// \Selector27~4_combout  = (\Selector27~2_combout ) # ((\Selector27~3_combout ) # ((Mux27 & \Selector0~8_combout )))

	.dataa(Mux271),
	.datab(\Selector27~2_combout ),
	.datac(\Selector0~8_combout ),
	.datad(\Selector27~3_combout ),
	.cin(gnd),
	.combout(\Selector27~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~4 .lut_mask = 16'hFFEC;
defparam \Selector27~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N18
cycloneive_lcell_comb \ShiftRight0~127 (
// Equation(s):
// \ShiftRight0~127_combout  = (\Mux34~3_combout  & (\ShiftRight0~140_combout )) # (!\Mux34~3_combout  & ((\ShiftRight0~135_combout )))

	.dataa(gnd),
	.datab(Mux34),
	.datac(\ShiftRight0~140_combout ),
	.datad(\ShiftRight0~135_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~127_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~127 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~127 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N28
cycloneive_lcell_comb \Selector27~5 (
// Equation(s):
// \Selector27~5_combout  = (\Selector5~1_combout  & ((\Selector5~0_combout ) # ((\ShiftRight0~127_combout )))) # (!\Selector5~1_combout  & (!\Selector5~0_combout  & (\ShiftRight0~134_combout )))

	.dataa(\Selector5~1_combout ),
	.datab(\Selector5~0_combout ),
	.datac(\ShiftRight0~134_combout ),
	.datad(\ShiftRight0~127_combout ),
	.cin(gnd),
	.combout(\Selector27~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~5 .lut_mask = 16'hBA98;
defparam \Selector27~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y39_N22
cycloneive_lcell_comb \Selector27~6 (
// Equation(s):
// \Selector27~6_combout  = (\Selector5~0_combout  & ((\Selector27~5_combout  & (\ShiftRight0~118_combout )) # (!\Selector27~5_combout  & ((\ShiftRight0~136_combout ))))) # (!\Selector5~0_combout  & (\Selector27~5_combout ))

	.dataa(\Selector5~0_combout ),
	.datab(\Selector27~5_combout ),
	.datac(\ShiftRight0~118_combout ),
	.datad(\ShiftRight0~136_combout ),
	.cin(gnd),
	.combout(\Selector27~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector27~6 .lut_mask = 16'hE6C4;
defparam \Selector27~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y38_N28
cycloneive_lcell_comb \Equal10~5 (
// Equation(s):
// \Equal10~5_combout  = (!Selector271 & (!Selector261 & (!Selector13 & !Selector12)))

	.dataa(Selector271),
	.datab(Selector261),
	.datac(Selector13),
	.datad(Selector12),
	.cin(gnd),
	.combout(\Equal10~5_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~5 .lut_mask = 16'h0001;
defparam \Equal10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N0
cycloneive_lcell_comb \Equal10~3 (
// Equation(s):
// \Equal10~3_combout  = (!Selector6 & (!Selector71 & !Selector10))

	.dataa(gnd),
	.datab(Selector6),
	.datac(Selector71),
	.datad(Selector10),
	.cin(gnd),
	.combout(\Equal10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~3 .lut_mask = 16'h0003;
defparam \Equal10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y38_N20
cycloneive_lcell_comb \Equal10~4 (
// Equation(s):
// \Equal10~4_combout  = (!Selector242 & (!Selector251 & (!Selector11 & \Equal10~3_combout )))

	.dataa(Selector242),
	.datab(Selector251),
	.datac(Selector11),
	.datad(\Equal10~3_combout ),
	.cin(gnd),
	.combout(\Equal10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~4 .lut_mask = 16'h0100;
defparam \Equal10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y36_N16
cycloneive_lcell_comb \Equal10~0 (
// Equation(s):
// \Equal10~0_combout  = (!Selector29 & (!Selector28 & (!Selector30 & !Selector5)))

	.dataa(Selector29),
	.datab(Selector28),
	.datac(Selector30),
	.datad(Selector5),
	.cin(gnd),
	.combout(\Equal10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~0 .lut_mask = 16'h0001;
defparam \Equal10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N28
cycloneive_lcell_comb \Equal10~1 (
// Equation(s):
// \Equal10~1_combout  = (!Selector3 & (!Selector41 & !Selector1))

	.dataa(gnd),
	.datab(Selector3),
	.datac(Selector41),
	.datad(Selector1),
	.cin(gnd),
	.combout(\Equal10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~1 .lut_mask = 16'h0003;
defparam \Equal10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N2
cycloneive_lcell_comb \Equal10~2 (
// Equation(s):
// \Equal10~2_combout  = (\Equal10~0_combout  & (!Selector0 & (!Selector2 & \Equal10~1_combout )))

	.dataa(\Equal10~0_combout ),
	.datab(Selector0),
	.datac(Selector2),
	.datad(\Equal10~1_combout ),
	.cin(gnd),
	.combout(\Equal10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~2 .lut_mask = 16'h0200;
defparam \Equal10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N0
cycloneive_lcell_comb \Selector14~4 (
// Equation(s):
// \Selector14~4_combout  = (\Mux19~1_combout  & (((\Selector0~15_combout )))) # (!\Mux19~1_combout  & (!Mux14 & ((\Selector0~18_combout ))))

	.dataa(Mux141),
	.datab(\Selector0~15_combout ),
	.datac(\Selector0~18_combout ),
	.datad(Mux192),
	.cin(gnd),
	.combout(\Selector14~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~4 .lut_mask = 16'hCC50;
defparam \Selector14~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N4
cycloneive_lcell_comb \Selector14~5 (
// Equation(s):
// \Selector14~5_combout  = (\Selector14~4_combout ) # ((\Selector0~17_combout  & (Mux14 $ (\Mux19~1_combout ))))

	.dataa(Mux141),
	.datab(\Selector0~17_combout ),
	.datac(\Selector14~4_combout ),
	.datad(Mux192),
	.cin(gnd),
	.combout(\Selector14~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~5 .lut_mask = 16'hF4F8;
defparam \Selector14~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N8
cycloneive_lcell_comb \Selector14~1 (
// Equation(s):
// \Selector14~1_combout  = (!cuifaluOp_0 & (\ShiftLeft0~99_combout  & \Selector16~1_combout ))

	.dataa(gnd),
	.datab(cuifaluOp_0),
	.datac(\ShiftLeft0~99_combout ),
	.datad(\Selector16~1_combout ),
	.cin(gnd),
	.combout(\Selector14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~1 .lut_mask = 16'h3000;
defparam \Selector14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N2
cycloneive_lcell_comb \Selector14~2 (
// Equation(s):
// \Selector14~2_combout  = (\Add1~34_combout  & ((\Selector0~19_combout ) # ((\Selector0~20_combout  & \Add0~34_combout )))) # (!\Add1~34_combout  & (\Selector0~20_combout  & ((\Add0~34_combout ))))

	.dataa(\Add1~34_combout ),
	.datab(\Selector0~20_combout ),
	.datac(\Selector0~19_combout ),
	.datad(\Add0~34_combout ),
	.cin(gnd),
	.combout(\Selector14~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~2 .lut_mask = 16'hECA0;
defparam \Selector14~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N12
cycloneive_lcell_comb \Selector14~6 (
// Equation(s):
// \Selector14~6_combout  = (\Selector14~3_combout ) # ((\Selector14~5_combout ) # ((\Selector14~1_combout ) # (\Selector14~2_combout )))

	.dataa(\Selector14~3_combout ),
	.datab(\Selector14~5_combout ),
	.datac(\Selector14~1_combout ),
	.datad(\Selector14~2_combout ),
	.cin(gnd),
	.combout(\Selector14~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~6 .lut_mask = 16'hFFFE;
defparam \Selector14~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N8
cycloneive_lcell_comb \Selector14~0 (
// Equation(s):
// \Selector14~0_combout  = (\Selector0~27_combout  & ((\Mux34~3_combout  & ((\ShiftLeft0~113_combout ))) # (!\Mux34~3_combout  & (\ShiftLeft0~114_combout ))))

	.dataa(\ShiftLeft0~114_combout ),
	.datab(Mux34),
	.datac(\ShiftLeft0~113_combout ),
	.datad(\Selector0~27_combout ),
	.cin(gnd),
	.combout(\Selector14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~0 .lut_mask = 16'hE200;
defparam \Selector14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N16
cycloneive_lcell_comb \Selector14~7 (
// Equation(s):
// \Selector14~7_combout  = (\Selector14~6_combout ) # ((\Selector14~0_combout ) # ((\Selector8~0_combout  & \ShiftRight0~83_combout )))

	.dataa(\Selector14~6_combout ),
	.datab(\Selector8~0_combout ),
	.datac(\ShiftRight0~83_combout ),
	.datad(\Selector14~0_combout ),
	.cin(gnd),
	.combout(\Selector14~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector14~7 .lut_mask = 16'hFFEA;
defparam \Selector14~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N30
cycloneive_lcell_comb \Selector15~0 (
// Equation(s):
// \Selector15~0_combout  = (\Selector0~27_combout  & ((\Mux34~3_combout  & ((\ShiftLeft0~126_combout ))) # (!\Mux34~3_combout  & (\ShiftLeft0~127_combout ))))

	.dataa(\Selector0~27_combout ),
	.datab(\ShiftLeft0~127_combout ),
	.datac(\ShiftLeft0~126_combout ),
	.datad(Mux34),
	.cin(gnd),
	.combout(\Selector15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~0 .lut_mask = 16'hA088;
defparam \Selector15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N0
cycloneive_lcell_comb \Selector15~4 (
// Equation(s):
// \Selector15~4_combout  = (\Mux20~1_combout  & (\Selector0~15_combout )) # (!\Mux20~1_combout  & (((\Selector0~18_combout  & !Mux15))))

	.dataa(Mux20),
	.datab(\Selector0~15_combout ),
	.datac(\Selector0~18_combout ),
	.datad(Mux152),
	.cin(gnd),
	.combout(\Selector15~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~4 .lut_mask = 16'h88D8;
defparam \Selector15~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N4
cycloneive_lcell_comb \Selector15~2 (
// Equation(s):
// \Selector15~2_combout  = (Mux15 & ((\Selector0~15_combout ) # ((\Selector0~16_combout  & \Mux20~1_combout ))))

	.dataa(\Selector0~16_combout ),
	.datab(Mux20),
	.datac(Mux152),
	.datad(\Selector0~15_combout ),
	.cin(gnd),
	.combout(\Selector15~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~2 .lut_mask = 16'hF080;
defparam \Selector15~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N28
cycloneive_lcell_comb \Selector15~1 (
// Equation(s):
// \Selector15~1_combout  = (\Add0~32_combout  & ((\Selector0~20_combout ) # ((\Selector0~19_combout  & \Add1~32_combout )))) # (!\Add0~32_combout  & (((\Selector0~19_combout  & \Add1~32_combout ))))

	.dataa(\Add0~32_combout ),
	.datab(\Selector0~20_combout ),
	.datac(\Selector0~19_combout ),
	.datad(\Add1~32_combout ),
	.cin(gnd),
	.combout(\Selector15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~1 .lut_mask = 16'hF888;
defparam \Selector15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N22
cycloneive_lcell_comb \Selector15~5 (
// Equation(s):
// \Selector15~5_combout  = (\Selector15~3_combout ) # ((\Selector15~4_combout ) # ((\Selector15~2_combout ) # (\Selector15~1_combout )))

	.dataa(\Selector15~3_combout ),
	.datab(\Selector15~4_combout ),
	.datac(\Selector15~2_combout ),
	.datad(\Selector15~1_combout ),
	.cin(gnd),
	.combout(\Selector15~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~5 .lut_mask = 16'hFFFE;
defparam \Selector15~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N28
cycloneive_lcell_comb \Selector15~6 (
// Equation(s):
// \Selector15~6_combout  = (\Selector15~5_combout ) # ((!\ShiftRight0~106_combout  & (Mux31 & \Selector0~29_combout )))

	.dataa(\ShiftRight0~106_combout ),
	.datab(Mux311),
	.datac(\Selector15~5_combout ),
	.datad(\Selector0~29_combout ),
	.cin(gnd),
	.combout(\Selector15~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~6 .lut_mask = 16'hF4F0;
defparam \Selector15~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N6
cycloneive_lcell_comb \Selector15~7 (
// Equation(s):
// \Selector15~7_combout  = (\Selector15~6_combout ) # ((!cuifaluOp_0 & (\Selector16~1_combout  & \ShiftLeft0~103_combout )))

	.dataa(cuifaluOp_0),
	.datab(\Selector16~1_combout ),
	.datac(\ShiftLeft0~103_combout ),
	.datad(\Selector15~6_combout ),
	.cin(gnd),
	.combout(\Selector15~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector15~7 .lut_mask = 16'hFF40;
defparam \Selector15~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N16
cycloneive_lcell_comb \Selector16~10 (
// Equation(s):
// \Selector16~10_combout  = (cuifaluOp_0 & \Selector16~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(cuifaluOp_0),
	.datad(\Selector16~1_combout ),
	.cin(gnd),
	.combout(\Selector16~10_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~10 .lut_mask = 16'hF000;
defparam \Selector16~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N12
cycloneive_lcell_comb \Selector0~39 (
// Equation(s):
// \Selector0~39_combout  = (cuifaluOp_0 & (\Mux33~3_combout  & (!\Mux32~4_combout  & \Selector0~21_combout )))

	.dataa(cuifaluOp_0),
	.datab(Mux33),
	.datac(Mux32),
	.datad(\Selector0~21_combout ),
	.cin(gnd),
	.combout(\Selector0~39_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~39 .lut_mask = 16'h0800;
defparam \Selector0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N8
cycloneive_lcell_comb \Selector16~2 (
// Equation(s):
// \Selector16~2_combout  = (\Mux34~3_combout  & (\ShiftRight0~145_combout )) # (!\Mux34~3_combout  & ((\ShiftRight0~146_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~145_combout ),
	.datac(Mux34),
	.datad(\ShiftRight0~146_combout ),
	.cin(gnd),
	.combout(\Selector16~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~2 .lut_mask = 16'hCFC0;
defparam \Selector16~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N14
cycloneive_lcell_comb \Selector16~3 (
// Equation(s):
// \Selector16~3_combout  = (\Selector0~39_combout  & ((\Selector16~2_combout ) # ((\Selector16~0_combout  & \ShiftLeft0~65_combout )))) # (!\Selector0~39_combout  & (((\Selector16~0_combout  & \ShiftLeft0~65_combout ))))

	.dataa(\Selector0~39_combout ),
	.datab(\Selector16~2_combout ),
	.datac(\Selector16~0_combout ),
	.datad(\ShiftLeft0~65_combout ),
	.cin(gnd),
	.combout(\Selector16~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~3 .lut_mask = 16'hF888;
defparam \Selector16~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y41_N24
cycloneive_lcell_comb \Selector16~4 (
// Equation(s):
// \Selector16~4_combout  = (Mux16 & ((\Selector0~15_combout ) # ((\Selector0~16_combout  & \Mux21~1_combout )))) # (!Mux16 & (((\Selector0~15_combout  & \Mux21~1_combout ))))

	.dataa(Mux161),
	.datab(\Selector0~16_combout ),
	.datac(\Selector0~15_combout ),
	.datad(Mux21),
	.cin(gnd),
	.combout(\Selector16~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~4 .lut_mask = 16'hF8A0;
defparam \Selector16~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N6
cycloneive_lcell_comb \Selector16~5 (
// Equation(s):
// \Selector16~5_combout  = (\Selector0~20_combout  & ((\Add0~30_combout ) # ((\Selector0~19_combout  & \Add1~30_combout )))) # (!\Selector0~20_combout  & (\Selector0~19_combout  & (\Add1~30_combout )))

	.dataa(\Selector0~20_combout ),
	.datab(\Selector0~19_combout ),
	.datac(\Add1~30_combout ),
	.datad(\Add0~30_combout ),
	.cin(gnd),
	.combout(\Selector16~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~5 .lut_mask = 16'hEAC0;
defparam \Selector16~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N20
cycloneive_lcell_comb \Selector16~6 (
// Equation(s):
// \Selector16~6_combout  = (\Selector16~5_combout ) # ((!\Mux21~1_combout  & (!Mux16 & \Selector0~18_combout )))

	.dataa(Mux21),
	.datab(Mux161),
	.datac(\Selector0~18_combout ),
	.datad(\Selector16~5_combout ),
	.cin(gnd),
	.combout(\Selector16~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~6 .lut_mask = 16'hFF10;
defparam \Selector16~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y38_N30
cycloneive_lcell_comb \Selector16~7 (
// Equation(s):
// \Selector16~7_combout  = (\Selector16~6_combout ) # ((\Selector0~17_combout  & (\Mux21~1_combout  $ (Mux16))))

	.dataa(\Selector0~17_combout ),
	.datab(Mux21),
	.datac(Mux161),
	.datad(\Selector16~6_combout ),
	.cin(gnd),
	.combout(\Selector16~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~7 .lut_mask = 16'hFF28;
defparam \Selector16~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N4
cycloneive_lcell_comb \Selector16~8 (
// Equation(s):
// \Selector16~8_combout  = (Mux0 & (!\Mux36~4_combout  & (\ShiftRight0~107_combout  & !\Mux35~4_combout )))

	.dataa(Mux0),
	.datab(Mux36),
	.datac(\ShiftRight0~107_combout ),
	.datad(Mux352),
	.cin(gnd),
	.combout(\Selector16~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~8 .lut_mask = 16'h0020;
defparam \Selector16~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y37_N20
cycloneive_lcell_comb \Selector16~9 (
// Equation(s):
// \Selector16~9_combout  = (\Selector16~4_combout ) # ((\Selector16~7_combout ) # ((\Selector20~0_combout  & \Selector16~8_combout )))

	.dataa(\Selector20~0_combout ),
	.datab(\Selector16~4_combout ),
	.datac(\Selector16~7_combout ),
	.datad(\Selector16~8_combout ),
	.cin(gnd),
	.combout(\Selector16~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector16~9 .lut_mask = 16'hFEFC;
defparam \Selector16~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N10
cycloneive_lcell_comb \ShiftRight0~123 (
// Equation(s):
// \ShiftRight0~123_combout  = (!\Selector0~30_combout  & ((\Mux36~4_combout  & ((Mux0))) # (!\Mux36~4_combout  & (Mux1))))

	.dataa(\Selector0~30_combout ),
	.datab(Mux1),
	.datac(Mux36),
	.datad(Mux0),
	.cin(gnd),
	.combout(\ShiftRight0~123_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~123 .lut_mask = 16'h5404;
defparam \ShiftRight0~123 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N24
cycloneive_lcell_comb \Selector9~0 (
// Equation(s):
// \Selector9~0_combout  = (\Mux34~3_combout  & (\ShiftLeft0~124_combout )) # (!\Mux34~3_combout  & ((\ShiftLeft0~120_combout )))

	.dataa(\ShiftLeft0~124_combout ),
	.datab(gnd),
	.datac(Mux34),
	.datad(\ShiftLeft0~120_combout ),
	.cin(gnd),
	.combout(\Selector9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~0 .lut_mask = 16'hAFA0;
defparam \Selector9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N30
cycloneive_lcell_comb \ShiftLeft0~95 (
// Equation(s):
// \ShiftLeft0~95_combout  = (\Mux33~3_combout  & (ShiftLeft03)) # (!\Mux33~3_combout  & ((\Selector9~0_combout )))

	.dataa(gnd),
	.datab(Mux33),
	.datac(ShiftLeft03),
	.datad(\Selector9~0_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~95_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~95 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y42_N4
cycloneive_lcell_comb \Selector17~0 (
// Equation(s):
// \Selector17~0_combout  = (\Selector0~39_combout  & ((\Mux34~3_combout  & ((\ShiftRight0~151_combout ))) # (!\Mux34~3_combout  & (\ShiftRight0~152_combout ))))

	.dataa(Mux34),
	.datab(\ShiftRight0~152_combout ),
	.datac(\ShiftRight0~151_combout ),
	.datad(\Selector0~39_combout ),
	.cin(gnd),
	.combout(\Selector17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~0 .lut_mask = 16'hE400;
defparam \Selector17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N8
cycloneive_lcell_comb \Selector17~1 (
// Equation(s):
// \Selector17~1_combout  = (\Selector0~15_combout  & (((Mux17) # (\Mux22~1_combout )))) # (!\Selector0~15_combout  & (\Selector0~16_combout  & (Mux17 & \Mux22~1_combout )))

	.dataa(\Selector0~15_combout ),
	.datab(\Selector0~16_combout ),
	.datac(Mux171),
	.datad(Mux22),
	.cin(gnd),
	.combout(\Selector17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~1 .lut_mask = 16'hEAA0;
defparam \Selector17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N18
cycloneive_lcell_comb \Selector17~2 (
// Equation(s):
// \Selector17~2_combout  = (\Selector0~20_combout  & ((\Add0~28_combout ) # ((\Selector0~19_combout  & \Add1~28_combout )))) # (!\Selector0~20_combout  & (((\Selector0~19_combout  & \Add1~28_combout ))))

	.dataa(\Selector0~20_combout ),
	.datab(\Add0~28_combout ),
	.datac(\Selector0~19_combout ),
	.datad(\Add1~28_combout ),
	.cin(gnd),
	.combout(\Selector17~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~2 .lut_mask = 16'hF888;
defparam \Selector17~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N18
cycloneive_lcell_comb \Selector17~3 (
// Equation(s):
// \Selector17~3_combout  = (\Selector17~2_combout ) # ((\Selector0~18_combout  & (!\Mux22~1_combout  & !Mux17)))

	.dataa(\Selector0~18_combout ),
	.datab(Mux22),
	.datac(Mux171),
	.datad(\Selector17~2_combout ),
	.cin(gnd),
	.combout(\Selector17~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~3 .lut_mask = 16'hFF02;
defparam \Selector17~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N28
cycloneive_lcell_comb \Selector17~4 (
// Equation(s):
// \Selector17~4_combout  = (\Selector17~3_combout ) # ((\Selector0~17_combout  & (\Mux22~1_combout  $ (Mux17))))

	.dataa(\Selector0~17_combout ),
	.datab(Mux22),
	.datac(Mux171),
	.datad(\Selector17~3_combout ),
	.cin(gnd),
	.combout(\Selector17~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~4 .lut_mask = 16'hFF28;
defparam \Selector17~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N14
cycloneive_lcell_comb \Selector17~5 (
// Equation(s):
// \Selector17~5_combout  = (\Selector17~1_combout ) # ((\Selector17~4_combout ) # ((\Selector16~10_combout  & \ShiftRight0~122_combout )))

	.dataa(\Selector16~10_combout ),
	.datab(\Selector17~1_combout ),
	.datac(\ShiftRight0~122_combout ),
	.datad(\Selector17~4_combout ),
	.cin(gnd),
	.combout(\Selector17~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~5 .lut_mask = 16'hFFEC;
defparam \Selector17~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y37_N10
cycloneive_lcell_comb \Selector17~6 (
// Equation(s):
// \Selector17~6_combout  = (\Selector17~0_combout ) # ((\Selector17~5_combout ) # ((\ShiftLeft0~95_combout  & \Selector16~0_combout )))

	.dataa(\ShiftLeft0~95_combout ),
	.datab(\Selector16~0_combout ),
	.datac(\Selector17~0_combout ),
	.datad(\Selector17~5_combout ),
	.cin(gnd),
	.combout(\Selector17~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector17~6 .lut_mask = 16'hFFF8;
defparam \Selector17~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N8
cycloneive_lcell_comb \Selector20~2 (
// Equation(s):
// \Selector20~2_combout  = (!\Mux33~3_combout  & (\ShiftRight0~110_combout  & \Selector20~0_combout ))

	.dataa(Mux33),
	.datab(gnd),
	.datac(\ShiftRight0~110_combout ),
	.datad(\Selector20~0_combout ),
	.cin(gnd),
	.combout(\Selector20~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~2 .lut_mask = 16'h5000;
defparam \Selector20~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N20
cycloneive_lcell_comb \Selector20~4 (
// Equation(s):
// \Selector20~4_combout  = (\Selector0~19_combout  & ((\Add1~22_combout ) # ((\Selector0~20_combout  & \Add0~22_combout )))) # (!\Selector0~19_combout  & (((\Selector0~20_combout  & \Add0~22_combout ))))

	.dataa(\Selector0~19_combout ),
	.datab(\Add1~22_combout ),
	.datac(\Selector0~20_combout ),
	.datad(\Add0~22_combout ),
	.cin(gnd),
	.combout(\Selector20~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~4 .lut_mask = 16'hF888;
defparam \Selector20~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N2
cycloneive_lcell_comb \Selector20~5 (
// Equation(s):
// \Selector20~5_combout  = (\Selector20~4_combout ) # ((!\Mux25~1_combout  & (\Selector0~18_combout  & !Mux20)))

	.dataa(Mux25),
	.datab(\Selector0~18_combout ),
	.datac(Mux201),
	.datad(\Selector20~4_combout ),
	.cin(gnd),
	.combout(\Selector20~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~5 .lut_mask = 16'hFF04;
defparam \Selector20~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N8
cycloneive_lcell_comb \Selector20~6 (
// Equation(s):
// \Selector20~6_combout  = (\Selector20~5_combout ) # ((\Selector0~17_combout  & (\Mux25~1_combout  $ (Mux20))))

	.dataa(Mux25),
	.datab(\Selector0~17_combout ),
	.datac(Mux201),
	.datad(\Selector20~5_combout ),
	.cin(gnd),
	.combout(\Selector20~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~6 .lut_mask = 16'hFF48;
defparam \Selector20~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N26
cycloneive_lcell_comb \Selector20~7 (
// Equation(s):
// \Selector20~7_combout  = (\Selector20~3_combout ) # ((\Selector20~6_combout ) # ((\Selector16~0_combout  & \ShiftLeft0~98_combout )))

	.dataa(\Selector20~3_combout ),
	.datab(\Selector16~0_combout ),
	.datac(\Selector20~6_combout ),
	.datad(\ShiftLeft0~98_combout ),
	.cin(gnd),
	.combout(\Selector20~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~7 .lut_mask = 16'hFEFA;
defparam \Selector20~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y36_N24
cycloneive_lcell_comb \Selector20~8 (
// Equation(s):
// \Selector20~8_combout  = (\Selector20~7_combout ) # ((\Selector20~1_combout  & \Selector0~39_combout ))

	.dataa(\Selector20~1_combout ),
	.datab(\Selector0~39_combout ),
	.datac(\Selector20~7_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector20~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector20~8 .lut_mask = 16'hF8F8;
defparam \Selector20~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N14
cycloneive_lcell_comb \Selector21~3 (
// Equation(s):
// \Selector21~3_combout  = (\Add1~20_combout  & ((\Selector0~19_combout ) # ((\Selector0~20_combout  & \Add0~20_combout )))) # (!\Add1~20_combout  & (((\Selector0~20_combout  & \Add0~20_combout ))))

	.dataa(\Add1~20_combout ),
	.datab(\Selector0~19_combout ),
	.datac(\Selector0~20_combout ),
	.datad(\Add0~20_combout ),
	.cin(gnd),
	.combout(\Selector21~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~3 .lut_mask = 16'hF888;
defparam \Selector21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N28
cycloneive_lcell_comb \Selector21~4 (
// Equation(s):
// \Selector21~4_combout  = (\Selector21~3_combout ) # ((\Selector0~18_combout  & (!Mux21 & !\Mux26~1_combout )))

	.dataa(\Selector0~18_combout ),
	.datab(Mux211),
	.datac(Mux26),
	.datad(\Selector21~3_combout ),
	.cin(gnd),
	.combout(\Selector21~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~4 .lut_mask = 16'hFF02;
defparam \Selector21~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N22
cycloneive_lcell_comb \Selector21~5 (
// Equation(s):
// \Selector21~5_combout  = (\Selector21~4_combout ) # ((\Selector0~17_combout  & (Mux21 $ (\Mux26~1_combout ))))

	.dataa(\Selector0~17_combout ),
	.datab(Mux211),
	.datac(Mux26),
	.datad(\Selector21~4_combout ),
	.cin(gnd),
	.combout(\Selector21~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~5 .lut_mask = 16'hFF28;
defparam \Selector21~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N8
cycloneive_lcell_comb \Selector21~6 (
// Equation(s):
// \Selector21~6_combout  = (\Selector21~2_combout ) # ((\Selector21~5_combout ) # ((\ShiftLeft0~88_combout  & \Selector16~0_combout )))

	.dataa(\Selector21~2_combout ),
	.datab(\ShiftLeft0~88_combout ),
	.datac(\Selector21~5_combout ),
	.datad(\Selector16~0_combout ),
	.cin(gnd),
	.combout(\Selector21~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~6 .lut_mask = 16'hFEFA;
defparam \Selector21~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N18
cycloneive_lcell_comb \Selector21~7 (
// Equation(s):
// \Selector21~7_combout  = (\Selector21~6_combout ) # ((\Selector0~39_combout  & \Selector21~0_combout ))

	.dataa(\Selector0~39_combout ),
	.datab(gnd),
	.datac(\Selector21~6_combout ),
	.datad(\Selector21~0_combout ),
	.cin(gnd),
	.combout(\Selector21~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~7 .lut_mask = 16'hFAF0;
defparam \Selector21~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N14
cycloneive_lcell_comb \Selector21~1 (
// Equation(s):
// \Selector21~1_combout  = (!\Mux33~3_combout  & (\ShiftRight0~113_combout  & \Selector20~0_combout ))

	.dataa(gnd),
	.datab(Mux33),
	.datac(\ShiftRight0~113_combout ),
	.datad(\Selector20~0_combout ),
	.cin(gnd),
	.combout(\Selector21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector21~1 .lut_mask = 16'h3000;
defparam \Selector21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N2
cycloneive_lcell_comb \Selector18~0 (
// Equation(s):
// \Selector18~0_combout  = (\Selector0~39_combout  & ((\Mux34~3_combout  & ((\ShiftRight0~131_combout ))) # (!\Mux34~3_combout  & (\ShiftRight0~132_combout ))))

	.dataa(Mux34),
	.datab(\ShiftRight0~132_combout ),
	.datac(\Selector0~39_combout ),
	.datad(\ShiftRight0~131_combout ),
	.cin(gnd),
	.combout(\Selector18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~0 .lut_mask = 16'hE040;
defparam \Selector18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N20
cycloneive_lcell_comb \Selector18~2 (
// Equation(s):
// \Selector18~2_combout  = (\Selector0~19_combout  & ((\Add1~26_combout ) # ((\Selector0~20_combout  & \Add0~26_combout )))) # (!\Selector0~19_combout  & (\Selector0~20_combout  & (\Add0~26_combout )))

	.dataa(\Selector0~19_combout ),
	.datab(\Selector0~20_combout ),
	.datac(\Add0~26_combout ),
	.datad(\Add1~26_combout ),
	.cin(gnd),
	.combout(\Selector18~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~2 .lut_mask = 16'hEAC0;
defparam \Selector18~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N18
cycloneive_lcell_comb \Selector18~3 (
// Equation(s):
// \Selector18~3_combout  = (\Selector18~2_combout ) # ((\Selector0~18_combout  & (!Mux18 & !\Mux23~1_combout )))

	.dataa(\Selector0~18_combout ),
	.datab(Mux181),
	.datac(Mux23),
	.datad(\Selector18~2_combout ),
	.cin(gnd),
	.combout(\Selector18~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~3 .lut_mask = 16'hFF02;
defparam \Selector18~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N4
cycloneive_lcell_comb \Selector18~4 (
// Equation(s):
// \Selector18~4_combout  = (\Selector18~3_combout ) # ((\Selector0~17_combout  & (Mux18 $ (\Mux23~1_combout ))))

	.dataa(\Selector0~17_combout ),
	.datab(Mux181),
	.datac(Mux23),
	.datad(\Selector18~3_combout ),
	.cin(gnd),
	.combout(\Selector18~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~4 .lut_mask = 16'hFF28;
defparam \Selector18~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N26
cycloneive_lcell_comb \Selector18~5 (
// Equation(s):
// \Selector18~5_combout  = (\Selector18~1_combout ) # ((\Selector18~4_combout ) # ((\ShiftLeft0~70_combout  & \Selector16~0_combout )))

	.dataa(\Selector18~1_combout ),
	.datab(\ShiftLeft0~70_combout ),
	.datac(\Selector18~4_combout ),
	.datad(\Selector16~0_combout ),
	.cin(gnd),
	.combout(\Selector18~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~5 .lut_mask = 16'hFEFA;
defparam \Selector18~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N16
cycloneive_lcell_comb \Selector18~6 (
// Equation(s):
// \Selector18~6_combout  = (\Selector18~0_combout ) # ((\Selector18~5_combout ) # ((\ShiftRight0~126_combout  & \Selector16~10_combout )))

	.dataa(\ShiftRight0~126_combout ),
	.datab(\Selector18~0_combout ),
	.datac(\Selector18~5_combout ),
	.datad(\Selector16~10_combout ),
	.cin(gnd),
	.combout(\Selector18~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector18~6 .lut_mask = 16'hFEFC;
defparam \Selector18~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N20
cycloneive_lcell_comb \Selector19~1 (
// Equation(s):
// \Selector19~1_combout  = (\Selector0~15_combout  & (((Mux19) # (\Mux24~1_combout )))) # (!\Selector0~15_combout  & (\Selector0~16_combout  & (Mux19 & \Mux24~1_combout )))

	.dataa(\Selector0~16_combout ),
	.datab(\Selector0~15_combout ),
	.datac(Mux191),
	.datad(Mux24),
	.cin(gnd),
	.combout(\Selector19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~1 .lut_mask = 16'hECC0;
defparam \Selector19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N6
cycloneive_lcell_comb \Selector19~2 (
// Equation(s):
// \Selector19~2_combout  = (\Add0~24_combout  & ((\Selector0~20_combout ) # ((\Selector0~19_combout  & \Add1~24_combout )))) # (!\Add0~24_combout  & (((\Selector0~19_combout  & \Add1~24_combout ))))

	.dataa(\Add0~24_combout ),
	.datab(\Selector0~20_combout ),
	.datac(\Selector0~19_combout ),
	.datad(\Add1~24_combout ),
	.cin(gnd),
	.combout(\Selector19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~2 .lut_mask = 16'hF888;
defparam \Selector19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N24
cycloneive_lcell_comb \Selector19~3 (
// Equation(s):
// \Selector19~3_combout  = (\Selector19~2_combout ) # ((!\Mux24~1_combout  & (\Selector0~18_combout  & !Mux19)))

	.dataa(Mux24),
	.datab(\Selector0~18_combout ),
	.datac(Mux191),
	.datad(\Selector19~2_combout ),
	.cin(gnd),
	.combout(\Selector19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~3 .lut_mask = 16'hFF04;
defparam \Selector19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N22
cycloneive_lcell_comb \Selector19~4 (
// Equation(s):
// \Selector19~4_combout  = (\Selector19~3_combout ) # ((\Selector0~17_combout  & (Mux19 $ (\Mux24~1_combout ))))

	.dataa(Mux191),
	.datab(\Selector19~3_combout ),
	.datac(\Selector0~17_combout ),
	.datad(Mux24),
	.cin(gnd),
	.combout(\Selector19~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~4 .lut_mask = 16'hDCEC;
defparam \Selector19~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N20
cycloneive_lcell_comb \Selector19~5 (
// Equation(s):
// \Selector19~5_combout  = (\Selector19~1_combout ) # ((\Selector19~4_combout ) # ((\ShiftLeft0~91_combout  & \Selector16~0_combout )))

	.dataa(\ShiftLeft0~91_combout ),
	.datab(\Selector19~1_combout ),
	.datac(\Selector19~4_combout ),
	.datad(\Selector16~0_combout ),
	.cin(gnd),
	.combout(\Selector19~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~5 .lut_mask = 16'hFEFC;
defparam \Selector19~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y39_N14
cycloneive_lcell_comb \Selector19~0 (
// Equation(s):
// \Selector19~0_combout  = (\Selector0~39_combout  & ((\Mux34~3_combout  & ((\ShiftRight0~138_combout ))) # (!\Mux34~3_combout  & (\ShiftRight0~139_combout ))))

	.dataa(\ShiftRight0~139_combout ),
	.datab(Mux34),
	.datac(\ShiftRight0~138_combout ),
	.datad(\Selector0~39_combout ),
	.cin(gnd),
	.combout(\Selector19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~0 .lut_mask = 16'hE200;
defparam \Selector19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N10
cycloneive_lcell_comb \Selector19~6 (
// Equation(s):
// \Selector19~6_combout  = (\Selector19~5_combout ) # ((\Selector19~0_combout ) # ((\Selector16~10_combout  & \ShiftRight0~127_combout )))

	.dataa(\Selector16~10_combout ),
	.datab(\ShiftRight0~127_combout ),
	.datac(\Selector19~5_combout ),
	.datad(\Selector19~0_combout ),
	.cin(gnd),
	.combout(\Selector19~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector19~6 .lut_mask = 16'hFFF8;
defparam \Selector19~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N14
cycloneive_lcell_comb \Selector8~5 (
// Equation(s):
// \Selector8~5_combout  = (Mux8 & ((\Selector0~15_combout ) # ((\Selector0~16_combout  & \Mux13~1_combout ))))

	.dataa(Mux81),
	.datab(\Selector0~15_combout ),
	.datac(\Selector0~16_combout ),
	.datad(Mux132),
	.cin(gnd),
	.combout(\Selector8~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~5 .lut_mask = 16'hA888;
defparam \Selector8~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N28
cycloneive_lcell_comb \Selector8~6 (
// Equation(s):
// \Selector8~6_combout  = (\Selector0~17_combout  & (Mux8 $ (((\Mux5~1_combout ) # (\Mux13~0_combout )))))

	.dataa(Mux81),
	.datab(Mux5),
	.datac(Mux13),
	.datad(\Selector0~17_combout ),
	.cin(gnd),
	.combout(\Selector8~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~6 .lut_mask = 16'h5600;
defparam \Selector8~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y42_N20
cycloneive_lcell_comb \Selector8~8 (
// Equation(s):
// \Selector8~8_combout  = (\Selector8~7_combout ) # ((\Selector8~5_combout ) # (\Selector8~6_combout ))

	.dataa(\Selector8~7_combout ),
	.datab(gnd),
	.datac(\Selector8~5_combout ),
	.datad(\Selector8~6_combout ),
	.cin(gnd),
	.combout(\Selector8~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~8 .lut_mask = 16'hFFFA;
defparam \Selector8~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N10
cycloneive_lcell_comb \Selector8~4 (
// Equation(s):
// \Selector8~4_combout  = (\Selector0~19_combout  & ((\Add1~46_combout ) # ((\Selector0~20_combout  & \Add0~46_combout )))) # (!\Selector0~19_combout  & (\Selector0~20_combout  & (\Add0~46_combout )))

	.dataa(\Selector0~19_combout ),
	.datab(\Selector0~20_combout ),
	.datac(\Add0~46_combout ),
	.datad(\Add1~46_combout ),
	.cin(gnd),
	.combout(\Selector8~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~4 .lut_mask = 16'hEAC0;
defparam \Selector8~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N20
cycloneive_lcell_comb \Selector8~9 (
// Equation(s):
// \Selector8~9_combout  = (\Selector8~8_combout ) # ((\Selector8~4_combout ) # ((\ShiftRight0~121_combout  & \Selector8~0_combout )))

	.dataa(\ShiftRight0~121_combout ),
	.datab(\Selector8~8_combout ),
	.datac(\Selector8~0_combout ),
	.datad(\Selector8~4_combout ),
	.cin(gnd),
	.combout(\Selector8~9_combout ),
	.cout());
// synopsys translate_off
defparam \Selector8~9 .lut_mask = 16'hFFEC;
defparam \Selector8~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N14
cycloneive_lcell_comb \Selector9~1 (
// Equation(s):
// \Selector9~1_combout  = (!cuifaluOp_0 & (\Selector1~6_combout  & \Selector16~1_combout ))

	.dataa(gnd),
	.datab(cuifaluOp_0),
	.datac(\Selector1~6_combout ),
	.datad(\Selector16~1_combout ),
	.cin(gnd),
	.combout(\Selector9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~1 .lut_mask = 16'h3000;
defparam \Selector9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N18
cycloneive_lcell_comb \Selector9~4 (
// Equation(s):
// \Selector9~4_combout  = (Mux9 & ((\Selector0~15_combout ) # ((\Selector0~16_combout  & \Mux14~1_combout ))))

	.dataa(Mux91),
	.datab(\Selector0~16_combout ),
	.datac(\Selector0~15_combout ),
	.datad(Mux14),
	.cin(gnd),
	.combout(\Selector9~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~4 .lut_mask = 16'hA8A0;
defparam \Selector9~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N4
cycloneive_lcell_comb \Selector9~3 (
// Equation(s):
// \Selector9~3_combout  = (\Add0~44_combout  & ((\Selector0~20_combout ) # ((\Selector0~19_combout  & \Add1~44_combout )))) # (!\Add0~44_combout  & (\Selector0~19_combout  & (\Add1~44_combout )))

	.dataa(\Add0~44_combout ),
	.datab(\Selector0~19_combout ),
	.datac(\Add1~44_combout ),
	.datad(\Selector0~20_combout ),
	.cin(gnd),
	.combout(\Selector9~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~3 .lut_mask = 16'hEAC0;
defparam \Selector9~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y38_N16
cycloneive_lcell_comb \Selector9~2 (
// Equation(s):
// \Selector9~2_combout  = (!\Mux32~4_combout  & (\ShiftRight0~125_combout  & (\Selector0~25_combout  & !\ShiftRight0~61_combout )))

	.dataa(Mux32),
	.datab(\ShiftRight0~125_combout ),
	.datac(\Selector0~25_combout ),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\Selector9~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~2 .lut_mask = 16'h0040;
defparam \Selector9~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N28
cycloneive_lcell_comb \Selector9~7 (
// Equation(s):
// \Selector9~7_combout  = (\Selector9~6_combout ) # ((\Selector9~4_combout ) # ((\Selector9~3_combout ) # (\Selector9~2_combout )))

	.dataa(\Selector9~6_combout ),
	.datab(\Selector9~4_combout ),
	.datac(\Selector9~3_combout ),
	.datad(\Selector9~2_combout ),
	.cin(gnd),
	.combout(\Selector9~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~7 .lut_mask = 16'hFFFE;
defparam \Selector9~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y39_N10
cycloneive_lcell_comb \Selector9~8 (
// Equation(s):
// \Selector9~8_combout  = (\Selector9~1_combout ) # ((\Selector9~7_combout ) # ((\Selector0~27_combout  & \Selector9~0_combout )))

	.dataa(\Selector0~27_combout ),
	.datab(\Selector9~0_combout ),
	.datac(\Selector9~1_combout ),
	.datad(\Selector9~7_combout ),
	.cin(gnd),
	.combout(\Selector9~8_combout ),
	.cout());
// synopsys translate_off
defparam \Selector9~8 .lut_mask = 16'hFFF8;
defparam \Selector9~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N28
cycloneive_lcell_comb \Selector22~2 (
// Equation(s):
// \Selector22~2_combout  = (\Mux27~1_combout  & ((\Selector0~15_combout ) # ((\Selector0~16_combout  & Mux22)))) # (!\Mux27~1_combout  & (((\Selector0~15_combout  & Mux22))))

	.dataa(\Selector0~16_combout ),
	.datab(Mux27),
	.datac(\Selector0~15_combout ),
	.datad(Mux221),
	.cin(gnd),
	.combout(\Selector22~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~2 .lut_mask = 16'hF8C0;
defparam \Selector22~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N6
cycloneive_lcell_comb \Selector22~3 (
// Equation(s):
// \Selector22~3_combout  = (\Add0~18_combout  & ((\Selector0~20_combout ) # ((\Selector0~19_combout  & \Add1~18_combout )))) # (!\Add0~18_combout  & (((\Selector0~19_combout  & \Add1~18_combout ))))

	.dataa(\Add0~18_combout ),
	.datab(\Selector0~20_combout ),
	.datac(\Selector0~19_combout ),
	.datad(\Add1~18_combout ),
	.cin(gnd),
	.combout(\Selector22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~3 .lut_mask = 16'hF888;
defparam \Selector22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N16
cycloneive_lcell_comb \Selector22~4 (
// Equation(s):
// \Selector22~4_combout  = (\Selector22~3_combout ) # ((\Selector0~18_combout  & (!Mux22 & !\Mux27~1_combout )))

	.dataa(\Selector0~18_combout ),
	.datab(Mux221),
	.datac(Mux27),
	.datad(\Selector22~3_combout ),
	.cin(gnd),
	.combout(\Selector22~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~4 .lut_mask = 16'hFF02;
defparam \Selector22~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N22
cycloneive_lcell_comb \Selector22~5 (
// Equation(s):
// \Selector22~5_combout  = (\Selector22~4_combout ) # ((\Selector0~17_combout  & (\Mux27~1_combout  $ (Mux22))))

	.dataa(Mux27),
	.datab(Mux221),
	.datac(\Selector0~17_combout ),
	.datad(\Selector22~4_combout ),
	.cin(gnd),
	.combout(\Selector22~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~5 .lut_mask = 16'hFF60;
defparam \Selector22~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N0
cycloneive_lcell_comb \Selector22~6 (
// Equation(s):
// \Selector22~6_combout  = (\Selector22~2_combout ) # ((\Selector22~5_combout ) # ((\ShiftLeft0~102_combout  & \Selector16~0_combout )))

	.dataa(\ShiftLeft0~102_combout ),
	.datab(\Selector22~2_combout ),
	.datac(\Selector22~5_combout ),
	.datad(\Selector16~0_combout ),
	.cin(gnd),
	.combout(\Selector22~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~6 .lut_mask = 16'hFEFC;
defparam \Selector22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N26
cycloneive_lcell_comb \Selector22~7 (
// Equation(s):
// \Selector22~7_combout  = (\Selector22~6_combout ) # ((\Selector22~0_combout  & \Selector0~39_combout ))

	.dataa(\Selector22~0_combout ),
	.datab(gnd),
	.datac(\Selector0~39_combout ),
	.datad(\Selector22~6_combout ),
	.cin(gnd),
	.combout(\Selector22~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~7 .lut_mask = 16'hFFA0;
defparam \Selector22~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N18
cycloneive_lcell_comb \Selector22~1 (
// Equation(s):
// \Selector22~1_combout  = (!\Mux33~3_combout  & (\ShiftRight0~78_combout  & \Selector20~0_combout ))

	.dataa(gnd),
	.datab(Mux33),
	.datac(\ShiftRight0~78_combout ),
	.datad(\Selector20~0_combout ),
	.cin(gnd),
	.combout(\Selector22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector22~1 .lut_mask = 16'h3000;
defparam \Selector22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N0
cycloneive_lcell_comb \Selector23~1 (
// Equation(s):
// \Selector23~1_combout  = (\Selector20~0_combout  & (!\Mux33~3_combout  & ShiftRight0))

	.dataa(\Selector20~0_combout ),
	.datab(Mux33),
	.datac(gnd),
	.datad(ShiftRight0),
	.cin(gnd),
	.combout(\Selector23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~1 .lut_mask = 16'h2200;
defparam \Selector23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N12
cycloneive_lcell_comb \Selector23~3 (
// Equation(s):
// \Selector23~3_combout  = (\Selector0~19_combout  & ((\Add1~16_combout ) # ((\Selector0~20_combout  & \Add0~16_combout )))) # (!\Selector0~19_combout  & (\Selector0~20_combout  & ((\Add0~16_combout ))))

	.dataa(\Selector0~19_combout ),
	.datab(\Selector0~20_combout ),
	.datac(\Add1~16_combout ),
	.datad(\Add0~16_combout ),
	.cin(gnd),
	.combout(\Selector23~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~3 .lut_mask = 16'hECA0;
defparam \Selector23~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N10
cycloneive_lcell_comb \Selector23~4 (
// Equation(s):
// \Selector23~4_combout  = (\Selector23~3_combout ) # ((\Selector0~18_combout  & (!Mux23 & !\Mux28~1_combout )))

	.dataa(\Selector0~18_combout ),
	.datab(Mux231),
	.datac(Mux28),
	.datad(\Selector23~3_combout ),
	.cin(gnd),
	.combout(\Selector23~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~4 .lut_mask = 16'hFF02;
defparam \Selector23~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N8
cycloneive_lcell_comb \Selector23~5 (
// Equation(s):
// \Selector23~5_combout  = (\Selector23~4_combout ) # ((\Selector0~17_combout  & (Mux23 $ (\Mux28~1_combout ))))

	.dataa(\Selector0~17_combout ),
	.datab(Mux231),
	.datac(Mux28),
	.datad(\Selector23~4_combout ),
	.cin(gnd),
	.combout(\Selector23~5_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~5 .lut_mask = 16'hFF28;
defparam \Selector23~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N14
cycloneive_lcell_comb \Selector23~6 (
// Equation(s):
// \Selector23~6_combout  = (\Selector23~2_combout ) # ((\Selector23~5_combout ) # ((\ShiftLeft0~105_combout  & \Selector16~0_combout )))

	.dataa(\Selector23~2_combout ),
	.datab(\ShiftLeft0~105_combout ),
	.datac(\Selector23~5_combout ),
	.datad(\Selector16~0_combout ),
	.cin(gnd),
	.combout(\Selector23~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~6 .lut_mask = 16'hFEFA;
defparam \Selector23~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N10
cycloneive_lcell_comb \Selector23~7 (
// Equation(s):
// \Selector23~7_combout  = (\Selector23~6_combout ) # ((\Selector0~39_combout  & \Selector23~0_combout ))

	.dataa(gnd),
	.datab(\Selector0~39_combout ),
	.datac(\Selector23~0_combout ),
	.datad(\Selector23~6_combout ),
	.cin(gnd),
	.combout(\Selector23~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector23~7 .lut_mask = 16'hFFC0;
defparam \Selector23~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y39_N22
cycloneive_lcell_comb \Equal10~8 (
// Equation(s):
// \Equal10~8_combout  = (!Selector81 & (!Selector8 & (!Selector82 & !Selector9)))

	.dataa(Selector81),
	.datab(Selector8),
	.datac(Selector82),
	.datad(Selector9),
	.cin(gnd),
	.combout(\Equal10~8_combout ),
	.cout());
// synopsys translate_off
defparam \Equal10~8 .lut_mask = 16'h0001;
defparam \Equal10~8 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module control_unit (
	always1,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	iwait,
	instr_28,
	instr_27,
	instr_29,
	instr_26,
	Equal12,
	instr_30,
	dcifimemload_30,
	instr_31,
	dcifimemload_31,
	dcifimemload_19,
	dcifimemload_29,
	dcifimemload_28,
	dcifimemload_26,
	dcifimemload_27,
	Equal2,
	Equal21,
	cuifregT_0,
	cuifregT_3,
	dcifimemload_18,
	cuifregT_2,
	dcifimemload_16,
	cuifregT_01,
	dcifimemload_17,
	cuifregT_1,
	dcifimemload_20,
	cuifregT_4,
	dcifimemload_3,
	dcifimemload_4,
	cuifaluOp_3,
	dcifimemload_0,
	dcifimemload_1,
	dcifimemload_2,
	dcifimemload_5,
	cuifaluOp_31,
	cuifaluOp_2,
	cuifaluOp_1,
	cuifaluOp_0,
	cuifaluSrc_0,
	WideOr4,
	Equal22,
	Equal0,
	cuifaluSrc_1,
	dcifimemload_23,
	cuifregS_2,
	dcifimemload_24,
	cuifregS_3,
	dcifimemload_21,
	cuifregS_0,
	dcifimemload_22,
	cuifregS_1,
	dcifimemload_25,
	cuifregS_4,
	cuifJmpSel_1,
	cuifJmpSel_0,
	Equal01,
	cuifMemtoReg_1,
	cuifMemtoReg_0,
	cuifRegDst_0,
	Equal23,
	devpor,
	devclrn,
	devoe);
input 	always1;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
input 	iwait;
input 	instr_28;
input 	instr_27;
input 	instr_29;
input 	instr_26;
output 	Equal12;
input 	instr_30;
input 	dcifimemload_30;
input 	instr_31;
input 	dcifimemload_31;
input 	dcifimemload_19;
input 	dcifimemload_29;
input 	dcifimemload_28;
input 	dcifimemload_26;
input 	dcifimemload_27;
output 	Equal2;
output 	Equal21;
output 	cuifregT_0;
output 	cuifregT_3;
input 	dcifimemload_18;
output 	cuifregT_2;
input 	dcifimemload_16;
output 	cuifregT_01;
input 	dcifimemload_17;
output 	cuifregT_1;
input 	dcifimemload_20;
output 	cuifregT_4;
input 	dcifimemload_3;
input 	dcifimemload_4;
output 	cuifaluOp_3;
input 	dcifimemload_0;
input 	dcifimemload_1;
input 	dcifimemload_2;
input 	dcifimemload_5;
output 	cuifaluOp_31;
output 	cuifaluOp_2;
output 	cuifaluOp_1;
output 	cuifaluOp_0;
output 	cuifaluSrc_0;
output 	WideOr4;
output 	Equal22;
output 	Equal0;
output 	cuifaluSrc_1;
input 	dcifimemload_23;
output 	cuifregS_2;
input 	dcifimemload_24;
output 	cuifregS_3;
input 	dcifimemload_21;
output 	cuifregS_0;
input 	dcifimemload_22;
output 	cuifregS_1;
input 	dcifimemload_25;
output 	cuifregS_4;
output 	cuifJmpSel_1;
output 	cuifJmpSel_0;
input 	Equal01;
output 	cuifMemtoReg_1;
output 	cuifMemtoReg_0;
output 	cuifRegDst_0;
output 	Equal23;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \WideOr4~1_combout ;
wire \Equal12~0_combout ;
wire \Equal12~1_combout ;
wire \Equal2~3_combout ;
wire \Equal2~2_combout ;
wire \Equal2~5_combout ;
wire \Equal2~6_combout ;
wire \cuif.regT[0]~0_combout ;
wire \cuif.aluOp[3]~0_combout ;
wire \cuif.MemtoReg[1]~0_combout ;
wire \WideOr1~0_combout ;
wire \cuif.aluOp[3]~2_combout ;
wire \cuif.aluOp[2]~5_combout ;
wire \cuif.aluOp[2]~6_combout ;
wire \cuif.aluOp[2]~7_combout ;
wire \cuif.aluOp[2]~4_combout ;
wire \cuif.aluOp[1]~9_combout ;
wire \cuif.aluOp[1]~10_combout ;
wire \cuif.aluOp[1]~11_combout ;
wire \cuif.aluOp[1]~12_combout ;
wire \WideOr4~0_combout ;
wire \cuif.aluOp[0]~15_combout ;
wire \cuif.aluOp[0]~16_combout ;
wire \cuif.aluOp[0]~14_combout ;
wire \cuif.JmpSel[1]~0_combout ;
wire \cuif.MemtoReg[1]~1_combout ;
wire \cuif.MemtoReg[0]~3_combout ;


// Location: LCCOMB_X55_Y35_N6
cycloneive_lcell_comb \WideOr4~1 (
// Equation(s):
// \WideOr4~1_combout  = (!dcifimemload_2 & (!dcifimemload_3 & (!dcifimemload_1 & !dcifimemload_0)))

	.dataa(dcifimemload_2),
	.datab(dcifimemload_3),
	.datac(dcifimemload_1),
	.datad(dcifimemload_0),
	.cin(gnd),
	.combout(\WideOr4~1_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr4~1 .lut_mask = 16'h0001;
defparam \WideOr4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N24
cycloneive_lcell_comb \Equal12~2 (
// Equation(s):
// Equal12 = (iwait & (\Equal12~0_combout )) # (!iwait & ((always1 & ((\Equal12~1_combout ))) # (!always1 & (\Equal12~0_combout ))))

	.dataa(\Equal12~0_combout ),
	.datab(iwait),
	.datac(always1),
	.datad(\Equal12~1_combout ),
	.cin(gnd),
	.combout(Equal12),
	.cout());
// synopsys translate_off
defparam \Equal12~2 .lut_mask = 16'hBA8A;
defparam \Equal12~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N10
cycloneive_lcell_comb \Equal2~4 (
// Equation(s):
// Equal2 = (iwait & (((\Equal2~3_combout )))) # (!iwait & ((always1 & ((\Equal2~2_combout ))) # (!always1 & (\Equal2~3_combout ))))

	.dataa(iwait),
	.datab(always1),
	.datac(\Equal2~3_combout ),
	.datad(\Equal2~2_combout ),
	.cin(gnd),
	.combout(Equal2),
	.cout());
// synopsys translate_off
defparam \Equal2~4 .lut_mask = 16'hF4B0;
defparam \Equal2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N18
cycloneive_lcell_comb \Equal2~7 (
// Equation(s):
// Equal21 = (iwait & (\Equal2~5_combout )) # (!iwait & ((always1 & ((\Equal2~6_combout ))) # (!always1 & (\Equal2~5_combout ))))

	.dataa(\Equal2~5_combout ),
	.datab(iwait),
	.datac(always1),
	.datad(\Equal2~6_combout ),
	.cin(gnd),
	.combout(Equal21),
	.cout());
// synopsys translate_off
defparam \Equal2~7 .lut_mask = 16'hBA8A;
defparam \Equal2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N28
cycloneive_lcell_comb \cuif.regT[0]~1 (
// Equation(s):
// cuifregT_0 = ((dcifimemload_30 & ((!Equal12))) # (!dcifimemload_30 & (!Equal21))) # (!dcifimemload_31)

	.dataa(dcifimemload_30),
	.datab(dcifimemload_31),
	.datac(Equal21),
	.datad(Equal12),
	.cin(gnd),
	.combout(cuifregT_0),
	.cout());
// synopsys translate_off
defparam \cuif.regT[0]~1 .lut_mask = 16'h37BF;
defparam \cuif.regT[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N22
cycloneive_lcell_comb \cuif.regT[3]~2 (
// Equation(s):
// cuifregT_3 = (dcifimemload_19 & (((Equal2 & \cuif.regT[0]~0_combout )) # (!cuifregT_0)))

	.dataa(Equal2),
	.datab(dcifimemload_19),
	.datac(\cuif.regT[0]~0_combout ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(cuifregT_3),
	.cout());
// synopsys translate_off
defparam \cuif.regT[3]~2 .lut_mask = 16'h80CC;
defparam \cuif.regT[3]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N8
cycloneive_lcell_comb \cuif.regT[2]~3 (
// Equation(s):
// cuifregT_2 = (dcifimemload_18 & (((\cuif.regT[0]~0_combout  & Equal2)) # (!cuifregT_0)))

	.dataa(dcifimemload_18),
	.datab(\cuif.regT[0]~0_combout ),
	.datac(Equal2),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(cuifregT_2),
	.cout());
// synopsys translate_off
defparam \cuif.regT[2]~3 .lut_mask = 16'h80AA;
defparam \cuif.regT[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N18
cycloneive_lcell_comb \cuif.regT[0]~4 (
// Equation(s):
// cuifregT_01 = (dcifimemload_16 & (((Equal2 & \cuif.regT[0]~0_combout )) # (!cuifregT_0)))

	.dataa(dcifimemload_16),
	.datab(Equal2),
	.datac(\cuif.regT[0]~0_combout ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(cuifregT_01),
	.cout());
// synopsys translate_off
defparam \cuif.regT[0]~4 .lut_mask = 16'h80AA;
defparam \cuif.regT[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N12
cycloneive_lcell_comb \cuif.regT[1]~5 (
// Equation(s):
// cuifregT_1 = (dcifimemload_17 & (((Equal2 & \cuif.regT[0]~0_combout )) # (!cuifregT_0)))

	.dataa(Equal2),
	.datab(\cuif.regT[0]~0_combout ),
	.datac(dcifimemload_17),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(cuifregT_1),
	.cout());
// synopsys translate_off
defparam \cuif.regT[1]~5 .lut_mask = 16'h80F0;
defparam \cuif.regT[1]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N10
cycloneive_lcell_comb \cuif.regT[4]~6 (
// Equation(s):
// cuifregT_4 = (dcifimemload_20 & (((Equal2 & \cuif.regT[0]~0_combout )) # (!cuifregT_0)))

	.dataa(Equal2),
	.datab(cuifregT_0),
	.datac(\cuif.regT[0]~0_combout ),
	.datad(dcifimemload_20),
	.cin(gnd),
	.combout(cuifregT_4),
	.cout());
// synopsys translate_off
defparam \cuif.regT[4]~6 .lut_mask = 16'hB300;
defparam \cuif.regT[4]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N12
cycloneive_lcell_comb \cuif.aluOp[3]~1 (
// Equation(s):
// cuifaluOp_3 = (!dcifimemload_26 & (!dcifimemload_27 & (!dcifimemload_28 & !dcifimemload_4)))

	.dataa(dcifimemload_26),
	.datab(dcifimemload_27),
	.datac(dcifimemload_28),
	.datad(dcifimemload_4),
	.cin(gnd),
	.combout(cuifaluOp_3),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[3]~1 .lut_mask = 16'h0001;
defparam \cuif.aluOp[3]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N14
cycloneive_lcell_comb \cuif.aluOp[3]~3 (
// Equation(s):
// cuifaluOp_31 = (Equal2 & ((dcifimemload_29 & (\cuif.aluOp[3]~0_combout )) # (!dcifimemload_29 & ((\cuif.aluOp[3]~2_combout )))))

	.dataa(Equal2),
	.datab(dcifimemload_29),
	.datac(\cuif.aluOp[3]~0_combout ),
	.datad(\cuif.aluOp[3]~2_combout ),
	.cin(gnd),
	.combout(cuifaluOp_31),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[3]~3 .lut_mask = 16'hA280;
defparam \cuif.aluOp[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N14
cycloneive_lcell_comb \cuif.aluOp[2]~8 (
// Equation(s):
// cuifaluOp_2 = (\cuif.aluOp[2]~4_combout ) # ((!dcifimemload_29 & (\cuif.aluOp[2]~7_combout  & !dcifimemload_27)))

	.dataa(dcifimemload_29),
	.datab(\cuif.aluOp[2]~7_combout ),
	.datac(\cuif.aluOp[2]~4_combout ),
	.datad(dcifimemload_27),
	.cin(gnd),
	.combout(cuifaluOp_2),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[2]~8 .lut_mask = 16'hF0F4;
defparam \cuif.aluOp[2]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N28
cycloneive_lcell_comb \cuif.aluOp[1]~13 (
// Equation(s):
// cuifaluOp_1 = (\cuif.aluOp[1]~9_combout ) # ((!dcifimemload_29 & \cuif.aluOp[1]~12_combout ))

	.dataa(dcifimemload_29),
	.datab(\cuif.aluOp[1]~9_combout ),
	.datac(\cuif.aluOp[1]~12_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(cuifaluOp_1),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[1]~13 .lut_mask = 16'hDCDC;
defparam \cuif.aluOp[1]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N16
cycloneive_lcell_comb \cuif.aluOp[0]~17 (
// Equation(s):
// cuifaluOp_0 = (Equal2 & ((\cuif.aluOp[0]~14_combout ) # ((\cuif.aluOp[0]~16_combout  & !dcifimemload_29))))

	.dataa(\cuif.aluOp[0]~16_combout ),
	.datab(\cuif.aluOp[0]~14_combout ),
	.datac(Equal2),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(cuifaluOp_0),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[0]~17 .lut_mask = 16'hC0E0;
defparam \cuif.aluOp[0]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N16
cycloneive_lcell_comb \cuif.aluSrc[0]~0 (
// Equation(s):
// cuifaluSrc_0 = (Equal2 & (dcifimemload_29)) # (!Equal2 & ((!cuifregT_0)))

	.dataa(gnd),
	.datab(dcifimemload_29),
	.datac(cuifregT_0),
	.datad(Equal2),
	.cin(gnd),
	.combout(cuifaluSrc_0),
	.cout());
// synopsys translate_off
defparam \cuif.aluSrc[0]~0 .lut_mask = 16'hCC0F;
defparam \cuif.aluSrc[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N4
cycloneive_lcell_comb \WideOr4~2 (
// Equation(s):
// WideOr4 = (!dcifimemload_3 & (!dcifimemload_0 & !dcifimemload_2))

	.dataa(dcifimemload_3),
	.datab(gnd),
	.datac(dcifimemload_0),
	.datad(dcifimemload_2),
	.cin(gnd),
	.combout(WideOr4),
	.cout());
// synopsys translate_off
defparam \WideOr4~2 .lut_mask = 16'h0005;
defparam \WideOr4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N18
cycloneive_lcell_comb \Equal2~8 (
// Equation(s):
// Equal22 = (!dcifimemload_30 & (!dcifimemload_31 & !dcifimemload_29))

	.dataa(dcifimemload_30),
	.datab(gnd),
	.datac(dcifimemload_31),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(Equal22),
	.cout());
// synopsys translate_off
defparam \Equal2~8 .lut_mask = 16'h0005;
defparam \Equal2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N18
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// Equal0 = (dcifimemload_28) # ((dcifimemload_27) # ((dcifimemload_26) # (!Equal22)))

	.dataa(dcifimemload_28),
	.datab(dcifimemload_27),
	.datac(dcifimemload_26),
	.datad(Equal22),
	.cin(gnd),
	.combout(Equal0),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'hFEFF;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N0
cycloneive_lcell_comb \cuif.aluSrc[1]~1 (
// Equation(s):
// cuifaluSrc_1 = (!dcifimemload_4 & (!dcifimemload_5 & (WideOr4 & !Equal0)))

	.dataa(dcifimemload_4),
	.datab(dcifimemload_5),
	.datac(WideOr4),
	.datad(Equal0),
	.cin(gnd),
	.combout(cuifaluSrc_1),
	.cout());
// synopsys translate_off
defparam \cuif.aluSrc[1]~1 .lut_mask = 16'h0010;
defparam \cuif.aluSrc[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N6
cycloneive_lcell_comb \cuif.regS[2]~0 (
// Equation(s):
// cuifregS_2 = (dcifimemload_23 & (((Equal2 & \cuif.regT[0]~0_combout )) # (!cuifregT_0)))

	.dataa(Equal2),
	.datab(dcifimemload_23),
	.datac(\cuif.regT[0]~0_combout ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(cuifregS_2),
	.cout());
// synopsys translate_off
defparam \cuif.regS[2]~0 .lut_mask = 16'h80CC;
defparam \cuif.regS[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N10
cycloneive_lcell_comb \cuif.regS[3]~1 (
// Equation(s):
// cuifregS_3 = (dcifimemload_24 & (((\cuif.regT[0]~0_combout  & Equal2)) # (!cuifregT_0)))

	.dataa(dcifimemload_24),
	.datab(cuifregT_0),
	.datac(\cuif.regT[0]~0_combout ),
	.datad(Equal2),
	.cin(gnd),
	.combout(cuifregS_3),
	.cout());
// synopsys translate_off
defparam \cuif.regS[3]~1 .lut_mask = 16'hA222;
defparam \cuif.regS[3]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N2
cycloneive_lcell_comb \cuif.regS[0]~2 (
// Equation(s):
// cuifregS_0 = (dcifimemload_21 & (((Equal2 & \cuif.regT[0]~0_combout )) # (!cuifregT_0)))

	.dataa(Equal2),
	.datab(dcifimemload_21),
	.datac(\cuif.regT[0]~0_combout ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(cuifregS_0),
	.cout());
// synopsys translate_off
defparam \cuif.regS[0]~2 .lut_mask = 16'h80CC;
defparam \cuif.regS[0]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N14
cycloneive_lcell_comb \cuif.regS[1]~3 (
// Equation(s):
// cuifregS_1 = (dcifimemload_22 & (((Equal2 & \cuif.regT[0]~0_combout )) # (!cuifregT_0)))

	.dataa(Equal2),
	.datab(dcifimemload_22),
	.datac(\cuif.regT[0]~0_combout ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(cuifregS_1),
	.cout());
// synopsys translate_off
defparam \cuif.regS[1]~3 .lut_mask = 16'h80CC;
defparam \cuif.regS[1]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N10
cycloneive_lcell_comb \cuif.regS[4]~4 (
// Equation(s):
// cuifregS_4 = (dcifimemload_25 & (((\cuif.regT[0]~0_combout  & Equal2)) # (!cuifregT_0)))

	.dataa(\cuif.regT[0]~0_combout ),
	.datab(dcifimemload_25),
	.datac(Equal2),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(cuifregS_4),
	.cout());
// synopsys translate_off
defparam \cuif.regS[4]~4 .lut_mask = 16'h80CC;
defparam \cuif.regS[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N6
cycloneive_lcell_comb \cuif.JmpSel[1]~1 (
// Equation(s):
// cuifJmpSel_1 = (!dcifimemload_5 & (!dcifimemload_2 & (\cuif.JmpSel[1]~0_combout  & \cuif.aluOp[2]~6_combout )))

	.dataa(dcifimemload_5),
	.datab(dcifimemload_2),
	.datac(\cuif.JmpSel[1]~0_combout ),
	.datad(\cuif.aluOp[2]~6_combout ),
	.cin(gnd),
	.combout(cuifJmpSel_1),
	.cout());
// synopsys translate_off
defparam \cuif.JmpSel[1]~1 .lut_mask = 16'h1000;
defparam \cuif.JmpSel[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N16
cycloneive_lcell_comb \cuif.JmpSel[0]~2 (
// Equation(s):
// cuifJmpSel_0 = (dcifimemload_27 & (!dcifimemload_28 & Equal22))

	.dataa(dcifimemload_27),
	.datab(dcifimemload_28),
	.datac(gnd),
	.datad(Equal22),
	.cin(gnd),
	.combout(cuifJmpSel_0),
	.cout());
// synopsys translate_off
defparam \cuif.JmpSel[0]~2 .lut_mask = 16'h2200;
defparam \cuif.JmpSel[0]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N6
cycloneive_lcell_comb \cuif.MemtoReg[1]~2 (
// Equation(s):
// cuifMemtoReg_1 = (\cuif.MemtoReg[1]~1_combout  & (Equal2 & ((Equal12) # (!dcifimemload_29))))

	.dataa(dcifimemload_29),
	.datab(\cuif.MemtoReg[1]~1_combout ),
	.datac(Equal2),
	.datad(Equal12),
	.cin(gnd),
	.combout(cuifMemtoReg_1),
	.cout());
// synopsys translate_off
defparam \cuif.MemtoReg[1]~2 .lut_mask = 16'hC040;
defparam \cuif.MemtoReg[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N0
cycloneive_lcell_comb \cuif.MemtoReg[0]~4 (
// Equation(s):
// cuifMemtoReg_0 = (Equal2 & (!dcifimemload_29 & ((\cuif.MemtoReg[0]~3_combout ) # (Equal21)))) # (!Equal2 & (!\cuif.MemtoReg[0]~3_combout ))

	.dataa(\cuif.MemtoReg[0]~3_combout ),
	.datab(Equal21),
	.datac(Equal2),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(cuifMemtoReg_0),
	.cout());
// synopsys translate_off
defparam \cuif.MemtoReg[0]~4 .lut_mask = 16'h05E5;
defparam \cuif.MemtoReg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N20
cycloneive_lcell_comb \cuif.RegDst[0]~0 (
// Equation(s):
// cuifRegDst_0 = (Equal22 & ((dcifimemload_28 & ((!dcifimemload_27))) # (!dcifimemload_28 & (!dcifimemload_26))))

	.dataa(dcifimemload_28),
	.datab(dcifimemload_26),
	.datac(Equal22),
	.datad(dcifimemload_27),
	.cin(gnd),
	.combout(cuifRegDst_0),
	.cout());
// synopsys translate_off
defparam \cuif.RegDst[0]~0 .lut_mask = 16'h10B0;
defparam \cuif.RegDst[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N26
cycloneive_lcell_comb \Equal2~9 (
// Equation(s):
// Equal23 = (!dcifimemload_31 & (Equal21 & (!dcifimemload_29 & !dcifimemload_30)))

	.dataa(dcifimemload_31),
	.datab(Equal21),
	.datac(dcifimemload_29),
	.datad(dcifimemload_30),
	.cin(gnd),
	.combout(Equal23),
	.cout());
// synopsys translate_off
defparam \Equal2~9 .lut_mask = 16'h0004;
defparam \Equal2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N4
cycloneive_lcell_comb \Equal12~0 (
// Equation(s):
// \Equal12~0_combout  = (instr_27 & (instr_28 & (instr_26 & instr_29)))

	.dataa(instr_27),
	.datab(instr_28),
	.datac(instr_26),
	.datad(instr_29),
	.cin(gnd),
	.combout(\Equal12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal12~0 .lut_mask = 16'h8000;
defparam \Equal12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N14
cycloneive_lcell_comb \Equal12~1 (
// Equation(s):
// \Equal12~1_combout  = (ramiframload_29 & (ramiframload_26 & (ramiframload_28 & ramiframload_27)))

	.dataa(ramiframload_29),
	.datab(ramiframload_26),
	.datac(ramiframload_28),
	.datad(ramiframload_27),
	.cin(gnd),
	.combout(\Equal12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal12~1 .lut_mask = 16'h8000;
defparam \Equal12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N12
cycloneive_lcell_comb \Equal2~3 (
// Equation(s):
// \Equal2~3_combout  = (!instr_30 & !instr_31)

	.dataa(gnd),
	.datab(instr_30),
	.datac(instr_31),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~3 .lut_mask = 16'h0303;
defparam \Equal2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y35_N0
cycloneive_lcell_comb \Equal2~2 (
// Equation(s):
// \Equal2~2_combout  = (iwait & (((!instr_31)))) # (!iwait & (!ramiframload_30 & (!ramiframload_31)))

	.dataa(ramiframload_30),
	.datab(ramiframload_31),
	.datac(instr_31),
	.datad(iwait),
	.cin(gnd),
	.combout(\Equal2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~2 .lut_mask = 16'h0F11;
defparam \Equal2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N0
cycloneive_lcell_comb \Equal2~5 (
// Equation(s):
// \Equal2~5_combout  = (instr_27 & (instr_26 & !instr_28))

	.dataa(instr_27),
	.datab(instr_26),
	.datac(gnd),
	.datad(instr_28),
	.cin(gnd),
	.combout(\Equal2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~5 .lut_mask = 16'h0088;
defparam \Equal2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N16
cycloneive_lcell_comb \Equal2~6 (
// Equation(s):
// \Equal2~6_combout  = (!ramiframload_28 & (ramiframload_26 & ramiframload_27))

	.dataa(ramiframload_28),
	.datab(gnd),
	.datac(ramiframload_26),
	.datad(ramiframload_27),
	.cin(gnd),
	.combout(\Equal2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~6 .lut_mask = 16'h5000;
defparam \Equal2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y35_N2
cycloneive_lcell_comb \cuif.regT[0]~0 (
// Equation(s):
// \cuif.regT[0]~0_combout  = (dcifimemload_29) # ((!dcifimemload_27 & ((dcifimemload_28) # (!dcifimemload_26))))

	.dataa(dcifimemload_27),
	.datab(dcifimemload_26),
	.datac(dcifimemload_28),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(\cuif.regT[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.regT[0]~0 .lut_mask = 16'hFF51;
defparam \cuif.regT[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N8
cycloneive_lcell_comb \cuif.aluOp[3]~0 (
// Equation(s):
// \cuif.aluOp[3]~0_combout  = (dcifimemload_28 & (Equal12 & ((Equal2)))) # (!dcifimemload_28 & (((dcifimemload_27))))

	.dataa(Equal12),
	.datab(dcifimemload_28),
	.datac(dcifimemload_27),
	.datad(Equal2),
	.cin(gnd),
	.combout(\cuif.aluOp[3]~0_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[3]~0 .lut_mask = 16'hB830;
defparam \cuif.aluOp[3]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N2
cycloneive_lcell_comb \cuif.MemtoReg[1]~0 (
// Equation(s):
// \cuif.MemtoReg[1]~0_combout  = (dcifimemload_27 & (dcifimemload_28 $ (((!Equal2) # (!Equal12)))))

	.dataa(Equal12),
	.datab(dcifimemload_28),
	.datac(dcifimemload_27),
	.datad(Equal2),
	.cin(gnd),
	.combout(\cuif.MemtoReg[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.MemtoReg[1]~0 .lut_mask = 16'h9030;
defparam \cuif.MemtoReg[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N18
cycloneive_lcell_comb \WideOr1~0 (
// Equation(s):
// \WideOr1~0_combout  = (dcifimemload_2) # ((dcifimemload_5 & ((!dcifimemload_1))) # (!dcifimemload_5 & ((dcifimemload_0) # (dcifimemload_1))))

	.dataa(dcifimemload_5),
	.datab(dcifimemload_0),
	.datac(dcifimemload_2),
	.datad(dcifimemload_1),
	.cin(gnd),
	.combout(\WideOr1~0_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr1~0 .lut_mask = 16'hF5FE;
defparam \WideOr1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N24
cycloneive_lcell_comb \cuif.aluOp[3]~2 (
// Equation(s):
// \cuif.aluOp[3]~2_combout  = (\cuif.MemtoReg[1]~0_combout ) # ((dcifimemload_3 & (cuifaluOp_3 & !\WideOr1~0_combout )))

	.dataa(dcifimemload_3),
	.datab(\cuif.MemtoReg[1]~0_combout ),
	.datac(cuifaluOp_3),
	.datad(\WideOr1~0_combout ),
	.cin(gnd),
	.combout(\cuif.aluOp[3]~2_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[3]~2 .lut_mask = 16'hCCEC;
defparam \cuif.aluOp[3]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N24
cycloneive_lcell_comb \cuif.aluOp[2]~5 (
// Equation(s):
// \cuif.aluOp[2]~5_combout  = (dcifimemload_26) # ((dcifimemload_4) # ((dcifimemload_3 & dcifimemload_5)))

	.dataa(dcifimemload_3),
	.datab(dcifimemload_26),
	.datac(dcifimemload_5),
	.datad(dcifimemload_4),
	.cin(gnd),
	.combout(\cuif.aluOp[2]~5_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[2]~5 .lut_mask = 16'hFFEC;
defparam \cuif.aluOp[2]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N22
cycloneive_lcell_comb \cuif.aluOp[2]~6 (
// Equation(s):
// \cuif.aluOp[2]~6_combout  = (!dcifimemload_0 & (dcifimemload_3 & !dcifimemload_1))

	.dataa(dcifimemload_0),
	.datab(gnd),
	.datac(dcifimemload_3),
	.datad(dcifimemload_1),
	.cin(gnd),
	.combout(\cuif.aluOp[2]~6_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[2]~6 .lut_mask = 16'h0050;
defparam \cuif.aluOp[2]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N16
cycloneive_lcell_comb \cuif.aluOp[2]~7 (
// Equation(s):
// \cuif.aluOp[2]~7_combout  = (\cuif.aluOp[2]~5_combout ) # ((dcifimemload_2 & (!dcifimemload_5)) # (!dcifimemload_2 & ((!\cuif.aluOp[2]~6_combout ))))

	.dataa(dcifimemload_5),
	.datab(\cuif.aluOp[2]~5_combout ),
	.datac(\cuif.aluOp[2]~6_combout ),
	.datad(dcifimemload_2),
	.cin(gnd),
	.combout(\cuif.aluOp[2]~7_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[2]~7 .lut_mask = 16'hDDCF;
defparam \cuif.aluOp[2]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N4
cycloneive_lcell_comb \cuif.aluOp[2]~4 (
// Equation(s):
// \cuif.aluOp[2]~4_combout  = (dcifimemload_31) # ((dcifimemload_30) # (dcifimemload_29 $ (dcifimemload_28)))

	.dataa(dcifimemload_29),
	.datab(dcifimemload_31),
	.datac(dcifimemload_28),
	.datad(dcifimemload_30),
	.cin(gnd),
	.combout(\cuif.aluOp[2]~4_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[2]~4 .lut_mask = 16'hFFDE;
defparam \cuif.aluOp[2]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N8
cycloneive_lcell_comb \cuif.aluOp[1]~9 (
// Equation(s):
// \cuif.aluOp[1]~9_combout  = ((dcifimemload_27) # ((dcifimemload_29 & !dcifimemload_28))) # (!Equal2)

	.dataa(dcifimemload_29),
	.datab(dcifimemload_28),
	.datac(Equal2),
	.datad(dcifimemload_27),
	.cin(gnd),
	.combout(\cuif.aluOp[1]~9_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[1]~9 .lut_mask = 16'hFF2F;
defparam \cuif.aluOp[1]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N26
cycloneive_lcell_comb \cuif.aluOp[1]~10 (
// Equation(s):
// \cuif.aluOp[1]~10_combout  = (dcifimemload_5 & ((dcifimemload_2 & (dcifimemload_1 & !dcifimemload_3)) # (!dcifimemload_2 & ((dcifimemload_1) # (!dcifimemload_3)))))

	.dataa(dcifimemload_2),
	.datab(dcifimemload_5),
	.datac(dcifimemload_1),
	.datad(dcifimemload_3),
	.cin(gnd),
	.combout(\cuif.aluOp[1]~10_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[1]~10 .lut_mask = 16'h40C4;
defparam \cuif.aluOp[1]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N20
cycloneive_lcell_comb \cuif.aluOp[1]~11 (
// Equation(s):
// \cuif.aluOp[1]~11_combout  = (\cuif.aluOp[1]~10_combout ) # ((!dcifimemload_2 & (!dcifimemload_5 & \cuif.aluOp[2]~6_combout )))

	.dataa(dcifimemload_2),
	.datab(dcifimemload_5),
	.datac(\cuif.aluOp[1]~10_combout ),
	.datad(\cuif.aluOp[2]~6_combout ),
	.cin(gnd),
	.combout(\cuif.aluOp[1]~11_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[1]~11 .lut_mask = 16'hF1F0;
defparam \cuif.aluOp[1]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N30
cycloneive_lcell_comb \cuif.aluOp[1]~12 (
// Equation(s):
// \cuif.aluOp[1]~12_combout  = (dcifimemload_26) # ((dcifimemload_28) # ((!dcifimemload_4 & \cuif.aluOp[1]~11_combout )))

	.dataa(dcifimemload_26),
	.datab(dcifimemload_4),
	.datac(dcifimemload_28),
	.datad(\cuif.aluOp[1]~11_combout ),
	.cin(gnd),
	.combout(\cuif.aluOp[1]~12_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[1]~12 .lut_mask = 16'hFBFA;
defparam \cuif.aluOp[1]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N26
cycloneive_lcell_comb \WideOr4~0 (
// Equation(s):
// \WideOr4~0_combout  = (dcifimemload_1 & ((dcifimemload_0) # (dcifimemload_3 $ (!dcifimemload_2)))) # (!dcifimemload_1 & ((dcifimemload_3) # ((dcifimemload_0 & dcifimemload_2))))

	.dataa(dcifimemload_1),
	.datab(dcifimemload_0),
	.datac(dcifimemload_3),
	.datad(dcifimemload_2),
	.cin(gnd),
	.combout(\WideOr4~0_combout ),
	.cout());
// synopsys translate_off
defparam \WideOr4~0 .lut_mask = 16'hFCDA;
defparam \WideOr4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N24
cycloneive_lcell_comb \cuif.aluOp[0]~15 (
// Equation(s):
// \cuif.aluOp[0]~15_combout  = (dcifimemload_4) # ((dcifimemload_5 & ((\WideOr4~0_combout ))) # (!dcifimemload_5 & (!\WideOr4~1_combout )))

	.dataa(\WideOr4~1_combout ),
	.datab(dcifimemload_5),
	.datac(dcifimemload_4),
	.datad(\WideOr4~0_combout ),
	.cin(gnd),
	.combout(\cuif.aluOp[0]~15_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[0]~15 .lut_mask = 16'hFDF1;
defparam \cuif.aluOp[0]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y35_N14
cycloneive_lcell_comb \cuif.aluOp[0]~16 (
// Equation(s):
// \cuif.aluOp[0]~16_combout  = (dcifimemload_27 & (((!dcifimemload_28)))) # (!dcifimemload_27 & ((dcifimemload_28) # ((!dcifimemload_26 & \cuif.aluOp[0]~15_combout ))))

	.dataa(dcifimemload_27),
	.datab(dcifimemload_26),
	.datac(dcifimemload_28),
	.datad(\cuif.aluOp[0]~15_combout ),
	.cin(gnd),
	.combout(\cuif.aluOp[0]~16_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[0]~16 .lut_mask = 16'h5B5A;
defparam \cuif.aluOp[0]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N0
cycloneive_lcell_comb \cuif.aluOp[0]~14 (
// Equation(s):
// \cuif.aluOp[0]~14_combout  = (dcifimemload_26 & (dcifimemload_29 & ((dcifimemload_28) # (dcifimemload_27))))

	.dataa(dcifimemload_26),
	.datab(dcifimemload_28),
	.datac(dcifimemload_27),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(\cuif.aluOp[0]~14_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.aluOp[0]~14 .lut_mask = 16'hA800;
defparam \cuif.aluOp[0]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N4
cycloneive_lcell_comb \cuif.JmpSel[1]~0 (
// Equation(s):
// \cuif.JmpSel[1]~0_combout  = (!Equal0 & !dcifimemload_4)

	.dataa(gnd),
	.datab(Equal0),
	.datac(gnd),
	.datad(dcifimemload_4),
	.cin(gnd),
	.combout(\cuif.JmpSel[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.JmpSel[1]~0 .lut_mask = 16'h0033;
defparam \cuif.JmpSel[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N24
cycloneive_lcell_comb \cuif.MemtoReg[1]~1 (
// Equation(s):
// \cuif.MemtoReg[1]~1_combout  = (dcifimemload_29 & (((dcifimemload_26)))) # (!dcifimemload_29 & ((Equal0) # ((\cuif.MemtoReg[1]~0_combout  & dcifimemload_26))))

	.dataa(\cuif.MemtoReg[1]~0_combout ),
	.datab(Equal01),
	.datac(dcifimemload_26),
	.datad(dcifimemload_29),
	.cin(gnd),
	.combout(\cuif.MemtoReg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.MemtoReg[1]~1 .lut_mask = 16'hF0EC;
defparam \cuif.MemtoReg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N26
cycloneive_lcell_comb \cuif.MemtoReg[0]~3 (
// Equation(s):
// \cuif.MemtoReg[0]~3_combout  = (Equal2 & (dcifimemload_28 & ((!cuifregT_0) # (!dcifimemload_27)))) # (!Equal2 & (((cuifregT_0))))

	.dataa(dcifimemload_27),
	.datab(Equal2),
	.datac(cuifregT_0),
	.datad(dcifimemload_28),
	.cin(gnd),
	.combout(\cuif.MemtoReg[0]~3_combout ),
	.cout());
// synopsys translate_off
defparam \cuif.MemtoReg[0]~3 .lut_mask = 16'h7C30;
defparam \cuif.MemtoReg[0]~3 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module pc_logic (
	pcifimemaddr_29,
	pcifimemaddr_28,
	pcifimemaddr_31,
	pcifimemaddr_30,
	dpifhalt,
	pcifimemaddr_1,
	ruifdmemREN,
	ruifdmemWEN,
	pcifimemaddr_0,
	pcifimemaddr_3,
	pcifimemaddr_2,
	pcifimemaddr_5,
	pcifimemaddr_4,
	pcifimemaddr_7,
	pcifimemaddr_6,
	pcifimemaddr_9,
	pcifimemaddr_8,
	pcifimemaddr_11,
	pcifimemaddr_10,
	pcifimemaddr_13,
	pcifimemaddr_12,
	pcifimemaddr_15,
	pcifimemaddr_14,
	pcifimemaddr_17,
	pcifimemaddr_16,
	pcifimemaddr_19,
	pcifimemaddr_18,
	pcifimemaddr_21,
	pcifimemaddr_20,
	pcifimemaddr_23,
	pcifimemaddr_22,
	pcifimemaddr_25,
	pcifimemaddr_24,
	pcifimemaddr_27,
	pcifimemaddr_26,
	always1,
	dcifimemload_19,
	dcifimemload_28,
	dcifimemload_27,
	dcifimemload_18,
	dcifimemload_16,
	dcifimemload_17,
	dcifimemload_20,
	dcifimemload_3,
	dcifimemload_4,
	dcifimemload_0,
	dcifimemload_1,
	dcifimemload_2,
	dcifimemload_5,
	dcifimemload_15,
	Equal2,
	dcifimemload_14,
	dcifimemload_13,
	dcifimemload_12,
	dcifimemload_11,
	dcifimemload_10,
	dcifimemload_9,
	dcifimemload_8,
	dcifimemload_7,
	dcifimemload_6,
	dcifimemload_23,
	dcifimemload_24,
	dcifimemload_21,
	dcifimemload_22,
	dcifimemload_25,
	Mux29,
	Mux30,
	Mux27,
	Mux28,
	Mux23,
	Mux24,
	Mux25,
	Mux26,
	Mux15,
	Mux16,
	Mux17,
	Mux18,
	Mux19,
	Mux20,
	Mux21,
	Mux22,
	Mux0,
	Mux2,
	Mux1,
	Mux3,
	Mux4,
	Mux5,
	Mux6,
	Mux7,
	Mux8,
	Mux9,
	Mux10,
	Mux11,
	Mux12,
	Mux13,
	Mux14,
	Mux31,
	cuifJmpSel_1,
	cuifJmpSel_0,
	Equal0,
	dcifimemload_26,
	Equal10,
	Equal101,
	Selector20,
	Selector21,
	Selector18,
	Selector19,
	Equal102,
	dcifimemload_261,
	CPUCLK,
	nRST,
	devpor,
	devclrn,
	devoe);
output 	pcifimemaddr_29;
output 	pcifimemaddr_28;
output 	pcifimemaddr_31;
output 	pcifimemaddr_30;
input 	dpifhalt;
output 	pcifimemaddr_1;
input 	ruifdmemREN;
input 	ruifdmemWEN;
output 	pcifimemaddr_0;
output 	pcifimemaddr_3;
output 	pcifimemaddr_2;
output 	pcifimemaddr_5;
output 	pcifimemaddr_4;
output 	pcifimemaddr_7;
output 	pcifimemaddr_6;
output 	pcifimemaddr_9;
output 	pcifimemaddr_8;
output 	pcifimemaddr_11;
output 	pcifimemaddr_10;
output 	pcifimemaddr_13;
output 	pcifimemaddr_12;
output 	pcifimemaddr_15;
output 	pcifimemaddr_14;
output 	pcifimemaddr_17;
output 	pcifimemaddr_16;
output 	pcifimemaddr_19;
output 	pcifimemaddr_18;
output 	pcifimemaddr_21;
output 	pcifimemaddr_20;
output 	pcifimemaddr_23;
output 	pcifimemaddr_22;
output 	pcifimemaddr_25;
output 	pcifimemaddr_24;
output 	pcifimemaddr_27;
output 	pcifimemaddr_26;
input 	always1;
input 	dcifimemload_19;
input 	dcifimemload_28;
input 	dcifimemload_27;
input 	dcifimemload_18;
input 	dcifimemload_16;
input 	dcifimemload_17;
input 	dcifimemload_20;
input 	dcifimemload_3;
input 	dcifimemload_4;
input 	dcifimemload_0;
input 	dcifimemload_1;
input 	dcifimemload_2;
input 	dcifimemload_5;
input 	dcifimemload_15;
input 	Equal2;
input 	dcifimemload_14;
input 	dcifimemload_13;
input 	dcifimemload_12;
input 	dcifimemload_11;
input 	dcifimemload_10;
input 	dcifimemload_9;
input 	dcifimemload_8;
input 	dcifimemload_7;
input 	dcifimemload_6;
input 	dcifimemload_23;
input 	dcifimemload_24;
input 	dcifimemload_21;
input 	dcifimemload_22;
input 	dcifimemload_25;
input 	Mux29;
input 	Mux30;
input 	Mux27;
input 	Mux28;
input 	Mux23;
input 	Mux24;
input 	Mux25;
input 	Mux26;
input 	Mux15;
input 	Mux16;
input 	Mux17;
input 	Mux18;
input 	Mux19;
input 	Mux20;
input 	Mux21;
input 	Mux22;
input 	Mux0;
input 	Mux2;
input 	Mux1;
input 	Mux3;
input 	Mux4;
input 	Mux5;
input 	Mux6;
input 	Mux7;
input 	Mux8;
input 	Mux9;
input 	Mux10;
input 	Mux11;
input 	Mux12;
input 	Mux13;
input 	Mux14;
input 	Mux31;
input 	cuifJmpSel_1;
input 	cuifJmpSel_0;
output 	Equal0;
input 	dcifimemload_26;
input 	Equal10;
input 	Equal101;
input 	Selector20;
input 	Selector21;
input 	Selector18;
input 	Selector19;
input 	Equal102;
input 	dcifimemload_261;
input 	CPUCLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~0_combout ;
wire \Add1~2_combout ;
wire \tempReg[5]~6_combout ;
wire \tempReg[7]~10_combout ;
wire \Add1~8_combout ;
wire \Add1~34_combout ;
wire \Add1~38_combout ;
wire \Add1~42_combout ;
wire \Add1~48_combout ;
wire \pcif.imemaddr[31]~9_combout ;
wire \tempReg[2]~1 ;
wire \tempReg[3]~3 ;
wire \tempReg[4]~5 ;
wire \tempReg[5]~7 ;
wire \tempReg[6]~9 ;
wire \tempReg[7]~11 ;
wire \tempReg[8]~13 ;
wire \tempReg[9]~15 ;
wire \tempReg[10]~17 ;
wire \tempReg[11]~19 ;
wire \tempReg[12]~21 ;
wire \tempReg[13]~23 ;
wire \tempReg[14]~25 ;
wire \tempReg[15]~27 ;
wire \tempReg[16]~29 ;
wire \tempReg[17]~31 ;
wire \tempReg[18]~33 ;
wire \tempReg[19]~35 ;
wire \tempReg[20]~37 ;
wire \tempReg[21]~39 ;
wire \tempReg[22]~41 ;
wire \tempReg[23]~43 ;
wire \tempReg[24]~45 ;
wire \tempReg[25]~47 ;
wire \tempReg[26]~49 ;
wire \tempReg[27]~51 ;
wire \tempReg[28]~52_combout ;
wire \tempReg[27]~50_combout ;
wire \tempReg[26]~48_combout ;
wire \tempReg[20]~36_combout ;
wire \tempReg[19]~34_combout ;
wire \tempReg[17]~30_combout ;
wire \tempReg[15]~26_combout ;
wire \tempReg[14]~24_combout ;
wire \tempReg[13]~22_combout ;
wire \tempReg[12]~20_combout ;
wire \tempReg[11]~18_combout ;
wire \tempReg[10]~16_combout ;
wire \tempReg[6]~8_combout ;
wire \tempReg[4]~4_combout ;
wire \tempReg[3]~2_combout ;
wire \Add1~1 ;
wire \Add1~3 ;
wire \Add1~5 ;
wire \Add1~7 ;
wire \Add1~9 ;
wire \Add1~11 ;
wire \Add1~13 ;
wire \Add1~15 ;
wire \Add1~17 ;
wire \Add1~19 ;
wire \Add1~21 ;
wire \Add1~23 ;
wire \Add1~25 ;
wire \Add1~27 ;
wire \Add1~29 ;
wire \Add1~31 ;
wire \Add1~33 ;
wire \Add1~35 ;
wire \Add1~37 ;
wire \Add1~39 ;
wire \Add1~41 ;
wire \Add1~43 ;
wire \Add1~45 ;
wire \Add1~47 ;
wire \Add1~49 ;
wire \Add1~51 ;
wire \Add1~53 ;
wire \Add1~54_combout ;
wire \pcif.imemaddr[31]~14_combout ;
wire \pcif.imemaddr[29]~1_combout ;
wire \tempReg[28]~53 ;
wire \tempReg[29]~54_combout ;
wire \pcif.imemaddr[31]~10_combout ;
wire \pcif.imemaddr[31]~15_combout ;
wire \pcif.imemaddr[31]~16_combout ;
wire \pcif.imemaddr[31]~11_combout ;
wire \pcif.imemaddr[31]~12_combout ;
wire \pcif.imemaddr[31]~13_combout ;
wire \Add1~52_combout ;
wire \pcif.imemaddr[28]~0_combout ;
wire \tempReg[29]~55 ;
wire \tempReg[30]~56_combout ;
wire \Add1~55 ;
wire \Add1~57 ;
wire \Add1~58_combout ;
wire \pcif.imemaddr[31]~3_combout ;
wire \tempReg[30]~57 ;
wire \tempReg[31]~58_combout ;
wire \Add1~56_combout ;
wire \pcif.imemaddr[30]~2_combout ;
wire \haltReg~0_combout ;
wire \pcif.imemaddr[1]~8_combout ;
wire \haltReg~1_combout ;
wire \haltReg[3]~2_combout ;
wire \haltReg[3]~3_combout ;
wire \tempReg[2]~0_combout ;
wire \haltReg[2]~4_combout ;
wire \haltReg[2]~5_combout ;
wire \Add1~6_combout ;
wire \haltReg[5]~6_combout ;
wire \haltReg[5]~7_combout ;
wire \Add1~4_combout ;
wire \haltReg[4]~8_combout ;
wire \haltReg[4]~9_combout ;
wire \Add1~10_combout ;
wire \haltReg[7]~10_combout ;
wire \haltReg[7]~11_combout ;
wire \haltReg[6]~12_combout ;
wire \haltReg[6]~13_combout ;
wire \Add1~14_combout ;
wire \tempReg[9]~14_combout ;
wire \haltReg[9]~14_combout ;
wire \haltReg[9]~15_combout ;
wire \tempReg[8]~12_combout ;
wire \Add1~12_combout ;
wire \haltReg[8]~16_combout ;
wire \haltReg[8]~17_combout ;
wire \Add1~18_combout ;
wire \haltReg[11]~18_combout ;
wire \haltReg[11]~19_combout ;
wire \Add1~16_combout ;
wire \haltReg[10]~20_combout ;
wire \haltReg[10]~21_combout ;
wire \Add1~22_combout ;
wire \haltReg[13]~22_combout ;
wire \haltReg[13]~23_combout ;
wire \Add1~20_combout ;
wire \haltReg[12]~24_combout ;
wire \haltReg[12]~25_combout ;
wire \Add1~26_combout ;
wire \haltReg[15]~26_combout ;
wire \haltReg[15]~27_combout ;
wire \Add1~24_combout ;
wire \haltReg[14]~28_combout ;
wire \haltReg[14]~29_combout ;
wire \Add1~30_combout ;
wire \haltReg[17]~30_combout ;
wire \haltReg[17]~31_combout ;
wire \tempReg[16]~28_combout ;
wire \Add1~28_combout ;
wire \haltReg[16]~32_combout ;
wire \haltReg[16]~33_combout ;
wire \haltReg[19]~34_combout ;
wire \haltReg[19]~35_combout ;
wire \tempReg[18]~32_combout ;
wire \Add1~32_combout ;
wire \haltReg[18]~36_combout ;
wire \haltReg[18]~37_combout ;
wire \tempReg[21]~38_combout ;
wire \haltReg[21]~38_combout ;
wire \haltReg[21]~39_combout ;
wire \Add1~36_combout ;
wire \haltReg[20]~40_combout ;
wire \haltReg[20]~41_combout ;
wire \tempReg[23]~42_combout ;
wire \haltReg[23]~42_combout ;
wire \haltReg[23]~43_combout ;
wire \tempReg[22]~40_combout ;
wire \Add1~40_combout ;
wire \haltReg[22]~44_combout ;
wire \haltReg[22]~45_combout ;
wire \tempReg[25]~46_combout ;
wire \Add1~46_combout ;
wire \haltReg[25]~46_combout ;
wire \haltReg[25]~47_combout ;
wire \tempReg[24]~44_combout ;
wire \Add1~44_combout ;
wire \haltReg[24]~48_combout ;
wire \haltReg[24]~49_combout ;
wire \Add1~50_combout ;
wire \haltReg[27]~50_combout ;
wire \haltReg[27]~51_combout ;
wire \haltReg[26]~52_combout ;
wire \haltReg[26]~53_combout ;


// Location: LCCOMB_X50_Y37_N2
cycloneive_lcell_comb \Add1~0 (
// Equation(s):
// \Add1~0_combout  = (\tempReg[2]~0_combout  & (dcifimemload_0 $ (VCC))) # (!\tempReg[2]~0_combout  & (dcifimemload_0 & VCC))
// \Add1~1  = CARRY((\tempReg[2]~0_combout  & dcifimemload_0))

	.dataa(\tempReg[2]~0_combout ),
	.datab(dcifimemload_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h6688;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N4
cycloneive_lcell_comb \Add1~2 (
// Equation(s):
// \Add1~2_combout  = (dcifimemload_1 & ((\tempReg[3]~2_combout  & (\Add1~1  & VCC)) # (!\tempReg[3]~2_combout  & (!\Add1~1 )))) # (!dcifimemload_1 & ((\tempReg[3]~2_combout  & (!\Add1~1 )) # (!\tempReg[3]~2_combout  & ((\Add1~1 ) # (GND)))))
// \Add1~3  = CARRY((dcifimemload_1 & (!\tempReg[3]~2_combout  & !\Add1~1 )) # (!dcifimemload_1 & ((!\Add1~1 ) # (!\tempReg[3]~2_combout ))))

	.dataa(dcifimemload_1),
	.datab(\tempReg[3]~2_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h9617;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N8
cycloneive_lcell_comb \tempReg[5]~6 (
// Equation(s):
// \tempReg[5]~6_combout  = (pcifimemaddr_5 & (!\tempReg[4]~5 )) # (!pcifimemaddr_5 & ((\tempReg[4]~5 ) # (GND)))
// \tempReg[5]~7  = CARRY((!\tempReg[4]~5 ) # (!pcifimemaddr_5))

	.dataa(gnd),
	.datab(pcifimemaddr_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[4]~5 ),
	.combout(\tempReg[5]~6_combout ),
	.cout(\tempReg[5]~7 ));
// synopsys translate_off
defparam \tempReg[5]~6 .lut_mask = 16'h3C3F;
defparam \tempReg[5]~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N12
cycloneive_lcell_comb \tempReg[7]~10 (
// Equation(s):
// \tempReg[7]~10_combout  = (pcifimemaddr_7 & (!\tempReg[6]~9 )) # (!pcifimemaddr_7 & ((\tempReg[6]~9 ) # (GND)))
// \tempReg[7]~11  = CARRY((!\tempReg[6]~9 ) # (!pcifimemaddr_7))

	.dataa(gnd),
	.datab(pcifimemaddr_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[6]~9 ),
	.combout(\tempReg[7]~10_combout ),
	.cout(\tempReg[7]~11 ));
// synopsys translate_off
defparam \tempReg[7]~10 .lut_mask = 16'h3C3F;
defparam \tempReg[7]~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N10
cycloneive_lcell_comb \Add1~8 (
// Equation(s):
// \Add1~8_combout  = ((dcifimemload_4 $ (\tempReg[6]~8_combout  $ (!\Add1~7 )))) # (GND)
// \Add1~9  = CARRY((dcifimemload_4 & ((\tempReg[6]~8_combout ) # (!\Add1~7 ))) # (!dcifimemload_4 & (\tempReg[6]~8_combout  & !\Add1~7 )))

	.dataa(dcifimemload_4),
	.datab(\tempReg[6]~8_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'h698E;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N4
cycloneive_lcell_comb \Add1~34 (
// Equation(s):
// \Add1~34_combout  = (dcifimemload_15 & ((\tempReg[19]~34_combout  & (\Add1~33  & VCC)) # (!\tempReg[19]~34_combout  & (!\Add1~33 )))) # (!dcifimemload_15 & ((\tempReg[19]~34_combout  & (!\Add1~33 )) # (!\tempReg[19]~34_combout  & ((\Add1~33 ) # (GND)))))
// \Add1~35  = CARRY((dcifimemload_15 & (!\tempReg[19]~34_combout  & !\Add1~33 )) # (!dcifimemload_15 & ((!\Add1~33 ) # (!\tempReg[19]~34_combout ))))

	.dataa(dcifimemload_15),
	.datab(\tempReg[19]~34_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~33 ),
	.combout(\Add1~34_combout ),
	.cout(\Add1~35 ));
// synopsys translate_off
defparam \Add1~34 .lut_mask = 16'h9617;
defparam \Add1~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N8
cycloneive_lcell_comb \Add1~38 (
// Equation(s):
// \Add1~38_combout  = (\tempReg[21]~38_combout  & ((dcifimemload_15 & (\Add1~37  & VCC)) # (!dcifimemload_15 & (!\Add1~37 )))) # (!\tempReg[21]~38_combout  & ((dcifimemload_15 & (!\Add1~37 )) # (!dcifimemload_15 & ((\Add1~37 ) # (GND)))))
// \Add1~39  = CARRY((\tempReg[21]~38_combout  & (!dcifimemload_15 & !\Add1~37 )) # (!\tempReg[21]~38_combout  & ((!\Add1~37 ) # (!dcifimemload_15))))

	.dataa(\tempReg[21]~38_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~37 ),
	.combout(\Add1~38_combout ),
	.cout(\Add1~39 ));
// synopsys translate_off
defparam \Add1~38 .lut_mask = 16'h9617;
defparam \Add1~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N12
cycloneive_lcell_comb \Add1~42 (
// Equation(s):
// \Add1~42_combout  = (\tempReg[23]~42_combout  & ((dcifimemload_15 & (\Add1~41  & VCC)) # (!dcifimemload_15 & (!\Add1~41 )))) # (!\tempReg[23]~42_combout  & ((dcifimemload_15 & (!\Add1~41 )) # (!dcifimemload_15 & ((\Add1~41 ) # (GND)))))
// \Add1~43  = CARRY((\tempReg[23]~42_combout  & (!dcifimemload_15 & !\Add1~41 )) # (!\tempReg[23]~42_combout  & ((!\Add1~41 ) # (!dcifimemload_15))))

	.dataa(\tempReg[23]~42_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~41 ),
	.combout(\Add1~42_combout ),
	.cout(\Add1~43 ));
// synopsys translate_off
defparam \Add1~42 .lut_mask = 16'h9617;
defparam \Add1~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N18
cycloneive_lcell_comb \Add1~48 (
// Equation(s):
// \Add1~48_combout  = ((dcifimemload_15 $ (\tempReg[26]~48_combout  $ (!\Add1~47 )))) # (GND)
// \Add1~49  = CARRY((dcifimemload_15 & ((\tempReg[26]~48_combout ) # (!\Add1~47 ))) # (!dcifimemload_15 & (\tempReg[26]~48_combout  & !\Add1~47 )))

	.dataa(dcifimemload_15),
	.datab(\tempReg[26]~48_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~47 ),
	.combout(\Add1~48_combout ),
	.cout(\Add1~49 ));
// synopsys translate_off
defparam \Add1~48 .lut_mask = 16'h698E;
defparam \Add1~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N12
cycloneive_lcell_comb \pcif.imemaddr[31]~9 (
// Equation(s):
// \pcif.imemaddr[31]~9_combout  = (!dcifimemload_27 & (dcifimemload_28 & Equal22))

	.dataa(dcifimemload_27),
	.datab(dcifimemload_28),
	.datac(gnd),
	.datad(Equal2),
	.cin(gnd),
	.combout(\pcif.imemaddr[31]~9_combout ),
	.cout());
// synopsys translate_off
defparam \pcif.imemaddr[31]~9 .lut_mask = 16'h4400;
defparam \pcif.imemaddr[31]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X50_Y36_N31
dffeas \pcif.imemaddr[29] (
	.clk(CPUCLK),
	.d(\pcif.imemaddr[29]~1_combout ),
	.asdata(\tempReg[29]~54_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(\pcif.imemaddr[31]~12_combout ),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_29),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[29] .is_wysiwyg = "true";
defparam \pcif.imemaddr[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N25
dffeas \pcif.imemaddr[28] (
	.clk(CPUCLK),
	.d(\pcif.imemaddr[28]~0_combout ),
	.asdata(\tempReg[28]~52_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(\pcif.imemaddr[31]~12_combout ),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_28),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[28] .is_wysiwyg = "true";
defparam \pcif.imemaddr[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N9
dffeas \pcif.imemaddr[31] (
	.clk(CPUCLK),
	.d(\pcif.imemaddr[31]~3_combout ),
	.asdata(\tempReg[31]~58_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(\pcif.imemaddr[31]~12_combout ),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_31),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[31] .is_wysiwyg = "true";
defparam \pcif.imemaddr[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N31
dffeas \pcif.imemaddr[30] (
	.clk(CPUCLK),
	.d(\pcif.imemaddr[30]~2_combout ),
	.asdata(\tempReg[30]~56_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(\pcif.imemaddr[31]~12_combout ),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_30),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[30] .is_wysiwyg = "true";
defparam \pcif.imemaddr[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N21
dffeas \pcif.imemaddr[1] (
	.clk(CPUCLK),
	.d(\haltReg~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_1),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[1] .is_wysiwyg = "true";
defparam \pcif.imemaddr[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y36_N1
dffeas \pcif.imemaddr[0] (
	.clk(CPUCLK),
	.d(\haltReg~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[1]~8_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_0),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[0] .is_wysiwyg = "true";
defparam \pcif.imemaddr[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N29
dffeas \pcif.imemaddr[3] (
	.clk(CPUCLK),
	.d(\haltReg[3]~3_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_3),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[3] .is_wysiwyg = "true";
defparam \pcif.imemaddr[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N7
dffeas \pcif.imemaddr[2] (
	.clk(CPUCLK),
	.d(\haltReg[2]~5_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_2),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[2] .is_wysiwyg = "true";
defparam \pcif.imemaddr[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N5
dffeas \pcif.imemaddr[5] (
	.clk(CPUCLK),
	.d(\haltReg[5]~7_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_5),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[5] .is_wysiwyg = "true";
defparam \pcif.imemaddr[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N21
dffeas \pcif.imemaddr[4] (
	.clk(CPUCLK),
	.d(\haltReg[4]~9_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_4),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[4] .is_wysiwyg = "true";
defparam \pcif.imemaddr[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y35_N31
dffeas \pcif.imemaddr[7] (
	.clk(CPUCLK),
	.d(\haltReg[7]~11_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_7),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[7] .is_wysiwyg = "true";
defparam \pcif.imemaddr[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y36_N19
dffeas \pcif.imemaddr[6] (
	.clk(CPUCLK),
	.d(\haltReg[6]~13_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_6),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[6] .is_wysiwyg = "true";
defparam \pcif.imemaddr[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N9
dffeas \pcif.imemaddr[9] (
	.clk(CPUCLK),
	.d(\haltReg[9]~15_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_9),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[9] .is_wysiwyg = "true";
defparam \pcif.imemaddr[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N27
dffeas \pcif.imemaddr[8] (
	.clk(CPUCLK),
	.d(\haltReg[8]~17_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_8),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[8] .is_wysiwyg = "true";
defparam \pcif.imemaddr[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N13
dffeas \pcif.imemaddr[11] (
	.clk(CPUCLK),
	.d(\haltReg[11]~19_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_11),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[11] .is_wysiwyg = "true";
defparam \pcif.imemaddr[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N31
dffeas \pcif.imemaddr[10] (
	.clk(CPUCLK),
	.d(\haltReg[10]~21_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_10),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[10] .is_wysiwyg = "true";
defparam \pcif.imemaddr[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N5
dffeas \pcif.imemaddr[13] (
	.clk(CPUCLK),
	.d(\haltReg[13]~23_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_13),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[13] .is_wysiwyg = "true";
defparam \pcif.imemaddr[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N23
dffeas \pcif.imemaddr[12] (
	.clk(CPUCLK),
	.d(\haltReg[12]~25_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_12),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[12] .is_wysiwyg = "true";
defparam \pcif.imemaddr[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N13
dffeas \pcif.imemaddr[15] (
	.clk(CPUCLK),
	.d(\haltReg[15]~27_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_15),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[15] .is_wysiwyg = "true";
defparam \pcif.imemaddr[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N3
dffeas \pcif.imemaddr[14] (
	.clk(CPUCLK),
	.d(\haltReg[14]~29_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_14),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[14] .is_wysiwyg = "true";
defparam \pcif.imemaddr[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N1
dffeas \pcif.imemaddr[17] (
	.clk(CPUCLK),
	.d(\haltReg[17]~31_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_17),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[17] .is_wysiwyg = "true";
defparam \pcif.imemaddr[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N7
dffeas \pcif.imemaddr[16] (
	.clk(CPUCLK),
	.d(\haltReg[16]~33_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_16),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[16] .is_wysiwyg = "true";
defparam \pcif.imemaddr[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y36_N13
dffeas \pcif.imemaddr[19] (
	.clk(CPUCLK),
	.d(\haltReg[19]~35_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_19),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[19] .is_wysiwyg = "true";
defparam \pcif.imemaddr[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N29
dffeas \pcif.imemaddr[18] (
	.clk(CPUCLK),
	.d(\haltReg[18]~37_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_18),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[18] .is_wysiwyg = "true";
defparam \pcif.imemaddr[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N5
dffeas \pcif.imemaddr[21] (
	.clk(CPUCLK),
	.d(\haltReg[21]~39_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_21),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[21] .is_wysiwyg = "true";
defparam \pcif.imemaddr[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N23
dffeas \pcif.imemaddr[20] (
	.clk(CPUCLK),
	.d(\haltReg[20]~41_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_20),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[20] .is_wysiwyg = "true";
defparam \pcif.imemaddr[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y35_N27
dffeas \pcif.imemaddr[23] (
	.clk(CPUCLK),
	.d(\haltReg[23]~43_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_23),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[23] .is_wysiwyg = "true";
defparam \pcif.imemaddr[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y36_N25
dffeas \pcif.imemaddr[22] (
	.clk(CPUCLK),
	.d(\haltReg[22]~45_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_22),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[22] .is_wysiwyg = "true";
defparam \pcif.imemaddr[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y36_N21
dffeas \pcif.imemaddr[25] (
	.clk(CPUCLK),
	.d(\haltReg[25]~47_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_25),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[25] .is_wysiwyg = "true";
defparam \pcif.imemaddr[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N5
dffeas \pcif.imemaddr[24] (
	.clk(CPUCLK),
	.d(\haltReg[24]~49_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_24),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[24] .is_wysiwyg = "true";
defparam \pcif.imemaddr[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y36_N19
dffeas \pcif.imemaddr[27] (
	.clk(CPUCLK),
	.d(\haltReg[27]~51_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_27),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[27] .is_wysiwyg = "true";
defparam \pcif.imemaddr[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N21
dffeas \pcif.imemaddr[26] (
	.clk(CPUCLK),
	.d(\haltReg[26]~53_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pcif.imemaddr[31]~13_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pcifimemaddr_26),
	.prn(vcc));
// synopsys translate_off
defparam \pcif.imemaddr[26] .is_wysiwyg = "true";
defparam \pcif.imemaddr[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N0
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// Equal0 = (dcifimemload_28 & !dcifimemload_27)

	.dataa(gnd),
	.datab(dcifimemload_28),
	.datac(gnd),
	.datad(dcifimemload_27),
	.cin(gnd),
	.combout(Equal0),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h00CC;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N2
cycloneive_lcell_comb \tempReg[2]~0 (
// Equation(s):
// \tempReg[2]~0_combout  = pcifimemaddr_2 $ (VCC)
// \tempReg[2]~1  = CARRY(pcifimemaddr_2)

	.dataa(pcifimemaddr_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\tempReg[2]~0_combout ),
	.cout(\tempReg[2]~1 ));
// synopsys translate_off
defparam \tempReg[2]~0 .lut_mask = 16'h55AA;
defparam \tempReg[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N4
cycloneive_lcell_comb \tempReg[3]~2 (
// Equation(s):
// \tempReg[3]~2_combout  = (pcifimemaddr_3 & (!\tempReg[2]~1 )) # (!pcifimemaddr_3 & ((\tempReg[2]~1 ) # (GND)))
// \tempReg[3]~3  = CARRY((!\tempReg[2]~1 ) # (!pcifimemaddr_3))

	.dataa(gnd),
	.datab(pcifimemaddr_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[2]~1 ),
	.combout(\tempReg[3]~2_combout ),
	.cout(\tempReg[3]~3 ));
// synopsys translate_off
defparam \tempReg[3]~2 .lut_mask = 16'h3C3F;
defparam \tempReg[3]~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N6
cycloneive_lcell_comb \tempReg[4]~4 (
// Equation(s):
// \tempReg[4]~4_combout  = (pcifimemaddr_4 & (\tempReg[3]~3  $ (GND))) # (!pcifimemaddr_4 & (!\tempReg[3]~3  & VCC))
// \tempReg[4]~5  = CARRY((pcifimemaddr_4 & !\tempReg[3]~3 ))

	.dataa(pcifimemaddr_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[3]~3 ),
	.combout(\tempReg[4]~4_combout ),
	.cout(\tempReg[4]~5 ));
// synopsys translate_off
defparam \tempReg[4]~4 .lut_mask = 16'hA50A;
defparam \tempReg[4]~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N10
cycloneive_lcell_comb \tempReg[6]~8 (
// Equation(s):
// \tempReg[6]~8_combout  = (pcifimemaddr_6 & (\tempReg[5]~7  $ (GND))) # (!pcifimemaddr_6 & (!\tempReg[5]~7  & VCC))
// \tempReg[6]~9  = CARRY((pcifimemaddr_6 & !\tempReg[5]~7 ))

	.dataa(gnd),
	.datab(pcifimemaddr_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[5]~7 ),
	.combout(\tempReg[6]~8_combout ),
	.cout(\tempReg[6]~9 ));
// synopsys translate_off
defparam \tempReg[6]~8 .lut_mask = 16'hC30C;
defparam \tempReg[6]~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N14
cycloneive_lcell_comb \tempReg[8]~12 (
// Equation(s):
// \tempReg[8]~12_combout  = (pcifimemaddr_8 & (\tempReg[7]~11  $ (GND))) # (!pcifimemaddr_8 & (!\tempReg[7]~11  & VCC))
// \tempReg[8]~13  = CARRY((pcifimemaddr_8 & !\tempReg[7]~11 ))

	.dataa(pcifimemaddr_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[7]~11 ),
	.combout(\tempReg[8]~12_combout ),
	.cout(\tempReg[8]~13 ));
// synopsys translate_off
defparam \tempReg[8]~12 .lut_mask = 16'hA50A;
defparam \tempReg[8]~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N16
cycloneive_lcell_comb \tempReg[9]~14 (
// Equation(s):
// \tempReg[9]~14_combout  = (pcifimemaddr_9 & (!\tempReg[8]~13 )) # (!pcifimemaddr_9 & ((\tempReg[8]~13 ) # (GND)))
// \tempReg[9]~15  = CARRY((!\tempReg[8]~13 ) # (!pcifimemaddr_9))

	.dataa(pcifimemaddr_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[8]~13 ),
	.combout(\tempReg[9]~14_combout ),
	.cout(\tempReg[9]~15 ));
// synopsys translate_off
defparam \tempReg[9]~14 .lut_mask = 16'h5A5F;
defparam \tempReg[9]~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N18
cycloneive_lcell_comb \tempReg[10]~16 (
// Equation(s):
// \tempReg[10]~16_combout  = (pcifimemaddr_10 & (\tempReg[9]~15  $ (GND))) # (!pcifimemaddr_10 & (!\tempReg[9]~15  & VCC))
// \tempReg[10]~17  = CARRY((pcifimemaddr_10 & !\tempReg[9]~15 ))

	.dataa(gnd),
	.datab(pcifimemaddr_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[9]~15 ),
	.combout(\tempReg[10]~16_combout ),
	.cout(\tempReg[10]~17 ));
// synopsys translate_off
defparam \tempReg[10]~16 .lut_mask = 16'hC30C;
defparam \tempReg[10]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N20
cycloneive_lcell_comb \tempReg[11]~18 (
// Equation(s):
// \tempReg[11]~18_combout  = (pcifimemaddr_11 & (!\tempReg[10]~17 )) # (!pcifimemaddr_11 & ((\tempReg[10]~17 ) # (GND)))
// \tempReg[11]~19  = CARRY((!\tempReg[10]~17 ) # (!pcifimemaddr_11))

	.dataa(gnd),
	.datab(pcifimemaddr_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[10]~17 ),
	.combout(\tempReg[11]~18_combout ),
	.cout(\tempReg[11]~19 ));
// synopsys translate_off
defparam \tempReg[11]~18 .lut_mask = 16'h3C3F;
defparam \tempReg[11]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N22
cycloneive_lcell_comb \tempReg[12]~20 (
// Equation(s):
// \tempReg[12]~20_combout  = (pcifimemaddr_12 & (\tempReg[11]~19  $ (GND))) # (!pcifimemaddr_12 & (!\tempReg[11]~19  & VCC))
// \tempReg[12]~21  = CARRY((pcifimemaddr_12 & !\tempReg[11]~19 ))

	.dataa(gnd),
	.datab(pcifimemaddr_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[11]~19 ),
	.combout(\tempReg[12]~20_combout ),
	.cout(\tempReg[12]~21 ));
// synopsys translate_off
defparam \tempReg[12]~20 .lut_mask = 16'hC30C;
defparam \tempReg[12]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N24
cycloneive_lcell_comb \tempReg[13]~22 (
// Equation(s):
// \tempReg[13]~22_combout  = (pcifimemaddr_13 & (!\tempReg[12]~21 )) # (!pcifimemaddr_13 & ((\tempReg[12]~21 ) # (GND)))
// \tempReg[13]~23  = CARRY((!\tempReg[12]~21 ) # (!pcifimemaddr_13))

	.dataa(pcifimemaddr_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[12]~21 ),
	.combout(\tempReg[13]~22_combout ),
	.cout(\tempReg[13]~23 ));
// synopsys translate_off
defparam \tempReg[13]~22 .lut_mask = 16'h5A5F;
defparam \tempReg[13]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N26
cycloneive_lcell_comb \tempReg[14]~24 (
// Equation(s):
// \tempReg[14]~24_combout  = (pcifimemaddr_14 & (\tempReg[13]~23  $ (GND))) # (!pcifimemaddr_14 & (!\tempReg[13]~23  & VCC))
// \tempReg[14]~25  = CARRY((pcifimemaddr_14 & !\tempReg[13]~23 ))

	.dataa(gnd),
	.datab(pcifimemaddr_14),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[13]~23 ),
	.combout(\tempReg[14]~24_combout ),
	.cout(\tempReg[14]~25 ));
// synopsys translate_off
defparam \tempReg[14]~24 .lut_mask = 16'hC30C;
defparam \tempReg[14]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N28
cycloneive_lcell_comb \tempReg[15]~26 (
// Equation(s):
// \tempReg[15]~26_combout  = (pcifimemaddr_15 & (!\tempReg[14]~25 )) # (!pcifimemaddr_15 & ((\tempReg[14]~25 ) # (GND)))
// \tempReg[15]~27  = CARRY((!\tempReg[14]~25 ) # (!pcifimemaddr_15))

	.dataa(pcifimemaddr_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[14]~25 ),
	.combout(\tempReg[15]~26_combout ),
	.cout(\tempReg[15]~27 ));
// synopsys translate_off
defparam \tempReg[15]~26 .lut_mask = 16'h5A5F;
defparam \tempReg[15]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y37_N30
cycloneive_lcell_comb \tempReg[16]~28 (
// Equation(s):
// \tempReg[16]~28_combout  = (pcifimemaddr_16 & (\tempReg[15]~27  $ (GND))) # (!pcifimemaddr_16 & (!\tempReg[15]~27  & VCC))
// \tempReg[16]~29  = CARRY((pcifimemaddr_16 & !\tempReg[15]~27 ))

	.dataa(gnd),
	.datab(pcifimemaddr_16),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[15]~27 ),
	.combout(\tempReg[16]~28_combout ),
	.cout(\tempReg[16]~29 ));
// synopsys translate_off
defparam \tempReg[16]~28 .lut_mask = 16'hC30C;
defparam \tempReg[16]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N0
cycloneive_lcell_comb \tempReg[17]~30 (
// Equation(s):
// \tempReg[17]~30_combout  = (pcifimemaddr_17 & (!\tempReg[16]~29 )) # (!pcifimemaddr_17 & ((\tempReg[16]~29 ) # (GND)))
// \tempReg[17]~31  = CARRY((!\tempReg[16]~29 ) # (!pcifimemaddr_17))

	.dataa(gnd),
	.datab(pcifimemaddr_17),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[16]~29 ),
	.combout(\tempReg[17]~30_combout ),
	.cout(\tempReg[17]~31 ));
// synopsys translate_off
defparam \tempReg[17]~30 .lut_mask = 16'h3C3F;
defparam \tempReg[17]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N2
cycloneive_lcell_comb \tempReg[18]~32 (
// Equation(s):
// \tempReg[18]~32_combout  = (pcifimemaddr_18 & (\tempReg[17]~31  $ (GND))) # (!pcifimemaddr_18 & (!\tempReg[17]~31  & VCC))
// \tempReg[18]~33  = CARRY((pcifimemaddr_18 & !\tempReg[17]~31 ))

	.dataa(pcifimemaddr_18),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[17]~31 ),
	.combout(\tempReg[18]~32_combout ),
	.cout(\tempReg[18]~33 ));
// synopsys translate_off
defparam \tempReg[18]~32 .lut_mask = 16'hA50A;
defparam \tempReg[18]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N4
cycloneive_lcell_comb \tempReg[19]~34 (
// Equation(s):
// \tempReg[19]~34_combout  = (pcifimemaddr_19 & (!\tempReg[18]~33 )) # (!pcifimemaddr_19 & ((\tempReg[18]~33 ) # (GND)))
// \tempReg[19]~35  = CARRY((!\tempReg[18]~33 ) # (!pcifimemaddr_19))

	.dataa(gnd),
	.datab(pcifimemaddr_19),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[18]~33 ),
	.combout(\tempReg[19]~34_combout ),
	.cout(\tempReg[19]~35 ));
// synopsys translate_off
defparam \tempReg[19]~34 .lut_mask = 16'h3C3F;
defparam \tempReg[19]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N6
cycloneive_lcell_comb \tempReg[20]~36 (
// Equation(s):
// \tempReg[20]~36_combout  = (pcifimemaddr_20 & (\tempReg[19]~35  $ (GND))) # (!pcifimemaddr_20 & (!\tempReg[19]~35  & VCC))
// \tempReg[20]~37  = CARRY((pcifimemaddr_20 & !\tempReg[19]~35 ))

	.dataa(gnd),
	.datab(pcifimemaddr_20),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[19]~35 ),
	.combout(\tempReg[20]~36_combout ),
	.cout(\tempReg[20]~37 ));
// synopsys translate_off
defparam \tempReg[20]~36 .lut_mask = 16'hC30C;
defparam \tempReg[20]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N8
cycloneive_lcell_comb \tempReg[21]~38 (
// Equation(s):
// \tempReg[21]~38_combout  = (pcifimemaddr_21 & (!\tempReg[20]~37 )) # (!pcifimemaddr_21 & ((\tempReg[20]~37 ) # (GND)))
// \tempReg[21]~39  = CARRY((!\tempReg[20]~37 ) # (!pcifimemaddr_21))

	.dataa(pcifimemaddr_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[20]~37 ),
	.combout(\tempReg[21]~38_combout ),
	.cout(\tempReg[21]~39 ));
// synopsys translate_off
defparam \tempReg[21]~38 .lut_mask = 16'h5A5F;
defparam \tempReg[21]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N10
cycloneive_lcell_comb \tempReg[22]~40 (
// Equation(s):
// \tempReg[22]~40_combout  = (pcifimemaddr_22 & (\tempReg[21]~39  $ (GND))) # (!pcifimemaddr_22 & (!\tempReg[21]~39  & VCC))
// \tempReg[22]~41  = CARRY((pcifimemaddr_22 & !\tempReg[21]~39 ))

	.dataa(gnd),
	.datab(pcifimemaddr_22),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[21]~39 ),
	.combout(\tempReg[22]~40_combout ),
	.cout(\tempReg[22]~41 ));
// synopsys translate_off
defparam \tempReg[22]~40 .lut_mask = 16'hC30C;
defparam \tempReg[22]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N12
cycloneive_lcell_comb \tempReg[23]~42 (
// Equation(s):
// \tempReg[23]~42_combout  = (pcifimemaddr_23 & (!\tempReg[22]~41 )) # (!pcifimemaddr_23 & ((\tempReg[22]~41 ) # (GND)))
// \tempReg[23]~43  = CARRY((!\tempReg[22]~41 ) # (!pcifimemaddr_23))

	.dataa(gnd),
	.datab(pcifimemaddr_23),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[22]~41 ),
	.combout(\tempReg[23]~42_combout ),
	.cout(\tempReg[23]~43 ));
// synopsys translate_off
defparam \tempReg[23]~42 .lut_mask = 16'h3C3F;
defparam \tempReg[23]~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N14
cycloneive_lcell_comb \tempReg[24]~44 (
// Equation(s):
// \tempReg[24]~44_combout  = (pcifimemaddr_24 & (\tempReg[23]~43  $ (GND))) # (!pcifimemaddr_24 & (!\tempReg[23]~43  & VCC))
// \tempReg[24]~45  = CARRY((pcifimemaddr_24 & !\tempReg[23]~43 ))

	.dataa(gnd),
	.datab(pcifimemaddr_24),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[23]~43 ),
	.combout(\tempReg[24]~44_combout ),
	.cout(\tempReg[24]~45 ));
// synopsys translate_off
defparam \tempReg[24]~44 .lut_mask = 16'hC30C;
defparam \tempReg[24]~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N16
cycloneive_lcell_comb \tempReg[25]~46 (
// Equation(s):
// \tempReg[25]~46_combout  = (pcifimemaddr_25 & (!\tempReg[24]~45 )) # (!pcifimemaddr_25 & ((\tempReg[24]~45 ) # (GND)))
// \tempReg[25]~47  = CARRY((!\tempReg[24]~45 ) # (!pcifimemaddr_25))

	.dataa(pcifimemaddr_25),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[24]~45 ),
	.combout(\tempReg[25]~46_combout ),
	.cout(\tempReg[25]~47 ));
// synopsys translate_off
defparam \tempReg[25]~46 .lut_mask = 16'h5A5F;
defparam \tempReg[25]~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N18
cycloneive_lcell_comb \tempReg[26]~48 (
// Equation(s):
// \tempReg[26]~48_combout  = (pcifimemaddr_26 & (\tempReg[25]~47  $ (GND))) # (!pcifimemaddr_26 & (!\tempReg[25]~47  & VCC))
// \tempReg[26]~49  = CARRY((pcifimemaddr_26 & !\tempReg[25]~47 ))

	.dataa(pcifimemaddr_26),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[25]~47 ),
	.combout(\tempReg[26]~48_combout ),
	.cout(\tempReg[26]~49 ));
// synopsys translate_off
defparam \tempReg[26]~48 .lut_mask = 16'hA50A;
defparam \tempReg[26]~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N20
cycloneive_lcell_comb \tempReg[27]~50 (
// Equation(s):
// \tempReg[27]~50_combout  = (pcifimemaddr_27 & (!\tempReg[26]~49 )) # (!pcifimemaddr_27 & ((\tempReg[26]~49 ) # (GND)))
// \tempReg[27]~51  = CARRY((!\tempReg[26]~49 ) # (!pcifimemaddr_27))

	.dataa(gnd),
	.datab(pcifimemaddr_27),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[26]~49 ),
	.combout(\tempReg[27]~50_combout ),
	.cout(\tempReg[27]~51 ));
// synopsys translate_off
defparam \tempReg[27]~50 .lut_mask = 16'h3C3F;
defparam \tempReg[27]~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N22
cycloneive_lcell_comb \tempReg[28]~52 (
// Equation(s):
// \tempReg[28]~52_combout  = (pcifimemaddr_28 & (\tempReg[27]~51  $ (GND))) # (!pcifimemaddr_28 & (!\tempReg[27]~51  & VCC))
// \tempReg[28]~53  = CARRY((pcifimemaddr_28 & !\tempReg[27]~51 ))

	.dataa(pcifimemaddr_28),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[27]~51 ),
	.combout(\tempReg[28]~52_combout ),
	.cout(\tempReg[28]~53 ));
// synopsys translate_off
defparam \tempReg[28]~52 .lut_mask = 16'hA50A;
defparam \tempReg[28]~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N6
cycloneive_lcell_comb \Add1~4 (
// Equation(s):
// \Add1~4_combout  = ((dcifimemload_2 $ (\tempReg[4]~4_combout  $ (!\Add1~3 )))) # (GND)
// \Add1~5  = CARRY((dcifimemload_2 & ((\tempReg[4]~4_combout ) # (!\Add1~3 ))) # (!dcifimemload_2 & (\tempReg[4]~4_combout  & !\Add1~3 )))

	.dataa(dcifimemload_2),
	.datab(\tempReg[4]~4_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'h698E;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N8
cycloneive_lcell_comb \Add1~6 (
// Equation(s):
// \Add1~6_combout  = (\tempReg[5]~6_combout  & ((dcifimemload_3 & (\Add1~5  & VCC)) # (!dcifimemload_3 & (!\Add1~5 )))) # (!\tempReg[5]~6_combout  & ((dcifimemload_3 & (!\Add1~5 )) # (!dcifimemload_3 & ((\Add1~5 ) # (GND)))))
// \Add1~7  = CARRY((\tempReg[5]~6_combout  & (!dcifimemload_3 & !\Add1~5 )) # (!\tempReg[5]~6_combout  & ((!\Add1~5 ) # (!dcifimemload_3))))

	.dataa(\tempReg[5]~6_combout ),
	.datab(dcifimemload_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h9617;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N12
cycloneive_lcell_comb \Add1~10 (
// Equation(s):
// \Add1~10_combout  = (\tempReg[7]~10_combout  & ((dcifimemload_5 & (\Add1~9  & VCC)) # (!dcifimemload_5 & (!\Add1~9 )))) # (!\tempReg[7]~10_combout  & ((dcifimemload_5 & (!\Add1~9 )) # (!dcifimemload_5 & ((\Add1~9 ) # (GND)))))
// \Add1~11  = CARRY((\tempReg[7]~10_combout  & (!dcifimemload_5 & !\Add1~9 )) # (!\tempReg[7]~10_combout  & ((!\Add1~9 ) # (!dcifimemload_5))))

	.dataa(\tempReg[7]~10_combout ),
	.datab(dcifimemload_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h9617;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N14
cycloneive_lcell_comb \Add1~12 (
// Equation(s):
// \Add1~12_combout  = ((\tempReg[8]~12_combout  $ (dcifimemload_6 $ (!\Add1~11 )))) # (GND)
// \Add1~13  = CARRY((\tempReg[8]~12_combout  & ((dcifimemload_6) # (!\Add1~11 ))) # (!\tempReg[8]~12_combout  & (dcifimemload_6 & !\Add1~11 )))

	.dataa(\tempReg[8]~12_combout ),
	.datab(dcifimemload_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout(\Add1~13 ));
// synopsys translate_off
defparam \Add1~12 .lut_mask = 16'h698E;
defparam \Add1~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N16
cycloneive_lcell_comb \Add1~14 (
// Equation(s):
// \Add1~14_combout  = (\tempReg[9]~14_combout  & ((dcifimemload_7 & (\Add1~13  & VCC)) # (!dcifimemload_7 & (!\Add1~13 )))) # (!\tempReg[9]~14_combout  & ((dcifimemload_7 & (!\Add1~13 )) # (!dcifimemload_7 & ((\Add1~13 ) # (GND)))))
// \Add1~15  = CARRY((\tempReg[9]~14_combout  & (!dcifimemload_7 & !\Add1~13 )) # (!\tempReg[9]~14_combout  & ((!\Add1~13 ) # (!dcifimemload_7))))

	.dataa(\tempReg[9]~14_combout ),
	.datab(dcifimemload_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~13 ),
	.combout(\Add1~14_combout ),
	.cout(\Add1~15 ));
// synopsys translate_off
defparam \Add1~14 .lut_mask = 16'h9617;
defparam \Add1~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N18
cycloneive_lcell_comb \Add1~16 (
// Equation(s):
// \Add1~16_combout  = ((dcifimemload_8 $ (\tempReg[10]~16_combout  $ (!\Add1~15 )))) # (GND)
// \Add1~17  = CARRY((dcifimemload_8 & ((\tempReg[10]~16_combout ) # (!\Add1~15 ))) # (!dcifimemload_8 & (\tempReg[10]~16_combout  & !\Add1~15 )))

	.dataa(dcifimemload_8),
	.datab(\tempReg[10]~16_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~15 ),
	.combout(\Add1~16_combout ),
	.cout(\Add1~17 ));
// synopsys translate_off
defparam \Add1~16 .lut_mask = 16'h698E;
defparam \Add1~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N20
cycloneive_lcell_comb \Add1~18 (
// Equation(s):
// \Add1~18_combout  = (dcifimemload_9 & ((\tempReg[11]~18_combout  & (\Add1~17  & VCC)) # (!\tempReg[11]~18_combout  & (!\Add1~17 )))) # (!dcifimemload_9 & ((\tempReg[11]~18_combout  & (!\Add1~17 )) # (!\tempReg[11]~18_combout  & ((\Add1~17 ) # (GND)))))
// \Add1~19  = CARRY((dcifimemload_9 & (!\tempReg[11]~18_combout  & !\Add1~17 )) # (!dcifimemload_9 & ((!\Add1~17 ) # (!\tempReg[11]~18_combout ))))

	.dataa(dcifimemload_9),
	.datab(\tempReg[11]~18_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~17 ),
	.combout(\Add1~18_combout ),
	.cout(\Add1~19 ));
// synopsys translate_off
defparam \Add1~18 .lut_mask = 16'h9617;
defparam \Add1~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N22
cycloneive_lcell_comb \Add1~20 (
// Equation(s):
// \Add1~20_combout  = ((dcifimemload_10 $ (\tempReg[12]~20_combout  $ (!\Add1~19 )))) # (GND)
// \Add1~21  = CARRY((dcifimemload_10 & ((\tempReg[12]~20_combout ) # (!\Add1~19 ))) # (!dcifimemload_10 & (\tempReg[12]~20_combout  & !\Add1~19 )))

	.dataa(dcifimemload_10),
	.datab(\tempReg[12]~20_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~19 ),
	.combout(\Add1~20_combout ),
	.cout(\Add1~21 ));
// synopsys translate_off
defparam \Add1~20 .lut_mask = 16'h698E;
defparam \Add1~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N24
cycloneive_lcell_comb \Add1~22 (
// Equation(s):
// \Add1~22_combout  = (dcifimemload_11 & ((\tempReg[13]~22_combout  & (\Add1~21  & VCC)) # (!\tempReg[13]~22_combout  & (!\Add1~21 )))) # (!dcifimemload_11 & ((\tempReg[13]~22_combout  & (!\Add1~21 )) # (!\tempReg[13]~22_combout  & ((\Add1~21 ) # (GND)))))
// \Add1~23  = CARRY((dcifimemload_11 & (!\tempReg[13]~22_combout  & !\Add1~21 )) # (!dcifimemload_11 & ((!\Add1~21 ) # (!\tempReg[13]~22_combout ))))

	.dataa(dcifimemload_11),
	.datab(\tempReg[13]~22_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~21 ),
	.combout(\Add1~22_combout ),
	.cout(\Add1~23 ));
// synopsys translate_off
defparam \Add1~22 .lut_mask = 16'h9617;
defparam \Add1~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N26
cycloneive_lcell_comb \Add1~24 (
// Equation(s):
// \Add1~24_combout  = ((dcifimemload_12 $ (\tempReg[14]~24_combout  $ (!\Add1~23 )))) # (GND)
// \Add1~25  = CARRY((dcifimemload_12 & ((\tempReg[14]~24_combout ) # (!\Add1~23 ))) # (!dcifimemload_12 & (\tempReg[14]~24_combout  & !\Add1~23 )))

	.dataa(dcifimemload_12),
	.datab(\tempReg[14]~24_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~23 ),
	.combout(\Add1~24_combout ),
	.cout(\Add1~25 ));
// synopsys translate_off
defparam \Add1~24 .lut_mask = 16'h698E;
defparam \Add1~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N28
cycloneive_lcell_comb \Add1~26 (
// Equation(s):
// \Add1~26_combout  = (dcifimemload_13 & ((\tempReg[15]~26_combout  & (\Add1~25  & VCC)) # (!\tempReg[15]~26_combout  & (!\Add1~25 )))) # (!dcifimemload_13 & ((\tempReg[15]~26_combout  & (!\Add1~25 )) # (!\tempReg[15]~26_combout  & ((\Add1~25 ) # (GND)))))
// \Add1~27  = CARRY((dcifimemload_13 & (!\tempReg[15]~26_combout  & !\Add1~25 )) # (!dcifimemload_13 & ((!\Add1~25 ) # (!\tempReg[15]~26_combout ))))

	.dataa(dcifimemload_13),
	.datab(\tempReg[15]~26_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~25 ),
	.combout(\Add1~26_combout ),
	.cout(\Add1~27 ));
// synopsys translate_off
defparam \Add1~26 .lut_mask = 16'h9617;
defparam \Add1~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y37_N30
cycloneive_lcell_comb \Add1~28 (
// Equation(s):
// \Add1~28_combout  = ((\tempReg[16]~28_combout  $ (dcifimemload_14 $ (!\Add1~27 )))) # (GND)
// \Add1~29  = CARRY((\tempReg[16]~28_combout  & ((dcifimemload_14) # (!\Add1~27 ))) # (!\tempReg[16]~28_combout  & (dcifimemload_14 & !\Add1~27 )))

	.dataa(\tempReg[16]~28_combout ),
	.datab(dcifimemload_14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~27 ),
	.combout(\Add1~28_combout ),
	.cout(\Add1~29 ));
// synopsys translate_off
defparam \Add1~28 .lut_mask = 16'h698E;
defparam \Add1~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N0
cycloneive_lcell_comb \Add1~30 (
// Equation(s):
// \Add1~30_combout  = (dcifimemload_15 & ((\tempReg[17]~30_combout  & (\Add1~29  & VCC)) # (!\tempReg[17]~30_combout  & (!\Add1~29 )))) # (!dcifimemload_15 & ((\tempReg[17]~30_combout  & (!\Add1~29 )) # (!\tempReg[17]~30_combout  & ((\Add1~29 ) # (GND)))))
// \Add1~31  = CARRY((dcifimemload_15 & (!\tempReg[17]~30_combout  & !\Add1~29 )) # (!dcifimemload_15 & ((!\Add1~29 ) # (!\tempReg[17]~30_combout ))))

	.dataa(dcifimemload_15),
	.datab(\tempReg[17]~30_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~29 ),
	.combout(\Add1~30_combout ),
	.cout(\Add1~31 ));
// synopsys translate_off
defparam \Add1~30 .lut_mask = 16'h9617;
defparam \Add1~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N2
cycloneive_lcell_comb \Add1~32 (
// Equation(s):
// \Add1~32_combout  = ((\tempReg[18]~32_combout  $ (dcifimemload_15 $ (!\Add1~31 )))) # (GND)
// \Add1~33  = CARRY((\tempReg[18]~32_combout  & ((dcifimemload_15) # (!\Add1~31 ))) # (!\tempReg[18]~32_combout  & (dcifimemload_15 & !\Add1~31 )))

	.dataa(\tempReg[18]~32_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~31 ),
	.combout(\Add1~32_combout ),
	.cout(\Add1~33 ));
// synopsys translate_off
defparam \Add1~32 .lut_mask = 16'h698E;
defparam \Add1~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N6
cycloneive_lcell_comb \Add1~36 (
// Equation(s):
// \Add1~36_combout  = ((dcifimemload_15 $ (\tempReg[20]~36_combout  $ (!\Add1~35 )))) # (GND)
// \Add1~37  = CARRY((dcifimemload_15 & ((\tempReg[20]~36_combout ) # (!\Add1~35 ))) # (!dcifimemload_15 & (\tempReg[20]~36_combout  & !\Add1~35 )))

	.dataa(dcifimemload_15),
	.datab(\tempReg[20]~36_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~35 ),
	.combout(\Add1~36_combout ),
	.cout(\Add1~37 ));
// synopsys translate_off
defparam \Add1~36 .lut_mask = 16'h698E;
defparam \Add1~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N10
cycloneive_lcell_comb \Add1~40 (
// Equation(s):
// \Add1~40_combout  = ((\tempReg[22]~40_combout  $ (dcifimemload_15 $ (!\Add1~39 )))) # (GND)
// \Add1~41  = CARRY((\tempReg[22]~40_combout  & ((dcifimemload_15) # (!\Add1~39 ))) # (!\tempReg[22]~40_combout  & (dcifimemload_15 & !\Add1~39 )))

	.dataa(\tempReg[22]~40_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~39 ),
	.combout(\Add1~40_combout ),
	.cout(\Add1~41 ));
// synopsys translate_off
defparam \Add1~40 .lut_mask = 16'h698E;
defparam \Add1~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N14
cycloneive_lcell_comb \Add1~44 (
// Equation(s):
// \Add1~44_combout  = ((\tempReg[24]~44_combout  $ (dcifimemload_15 $ (!\Add1~43 )))) # (GND)
// \Add1~45  = CARRY((\tempReg[24]~44_combout  & ((dcifimemload_15) # (!\Add1~43 ))) # (!\tempReg[24]~44_combout  & (dcifimemload_15 & !\Add1~43 )))

	.dataa(\tempReg[24]~44_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~43 ),
	.combout(\Add1~44_combout ),
	.cout(\Add1~45 ));
// synopsys translate_off
defparam \Add1~44 .lut_mask = 16'h698E;
defparam \Add1~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N16
cycloneive_lcell_comb \Add1~46 (
// Equation(s):
// \Add1~46_combout  = (\tempReg[25]~46_combout  & ((dcifimemload_15 & (\Add1~45  & VCC)) # (!dcifimemload_15 & (!\Add1~45 )))) # (!\tempReg[25]~46_combout  & ((dcifimemload_15 & (!\Add1~45 )) # (!dcifimemload_15 & ((\Add1~45 ) # (GND)))))
// \Add1~47  = CARRY((\tempReg[25]~46_combout  & (!dcifimemload_15 & !\Add1~45 )) # (!\tempReg[25]~46_combout  & ((!\Add1~45 ) # (!dcifimemload_15))))

	.dataa(\tempReg[25]~46_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~45 ),
	.combout(\Add1~46_combout ),
	.cout(\Add1~47 ));
// synopsys translate_off
defparam \Add1~46 .lut_mask = 16'h9617;
defparam \Add1~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N20
cycloneive_lcell_comb \Add1~50 (
// Equation(s):
// \Add1~50_combout  = (dcifimemload_15 & ((\tempReg[27]~50_combout  & (\Add1~49  & VCC)) # (!\tempReg[27]~50_combout  & (!\Add1~49 )))) # (!dcifimemload_15 & ((\tempReg[27]~50_combout  & (!\Add1~49 )) # (!\tempReg[27]~50_combout  & ((\Add1~49 ) # (GND)))))
// \Add1~51  = CARRY((dcifimemload_15 & (!\tempReg[27]~50_combout  & !\Add1~49 )) # (!dcifimemload_15 & ((!\Add1~49 ) # (!\tempReg[27]~50_combout ))))

	.dataa(dcifimemload_15),
	.datab(\tempReg[27]~50_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~49 ),
	.combout(\Add1~50_combout ),
	.cout(\Add1~51 ));
// synopsys translate_off
defparam \Add1~50 .lut_mask = 16'h9617;
defparam \Add1~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N22
cycloneive_lcell_comb \Add1~52 (
// Equation(s):
// \Add1~52_combout  = ((dcifimemload_15 $ (\tempReg[28]~52_combout  $ (!\Add1~51 )))) # (GND)
// \Add1~53  = CARRY((dcifimemload_15 & ((\tempReg[28]~52_combout ) # (!\Add1~51 ))) # (!dcifimemload_15 & (\tempReg[28]~52_combout  & !\Add1~51 )))

	.dataa(dcifimemload_15),
	.datab(\tempReg[28]~52_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~51 ),
	.combout(\Add1~52_combout ),
	.cout(\Add1~53 ));
// synopsys translate_off
defparam \Add1~52 .lut_mask = 16'h698E;
defparam \Add1~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N24
cycloneive_lcell_comb \Add1~54 (
// Equation(s):
// \Add1~54_combout  = (\tempReg[29]~54_combout  & ((dcifimemload_15 & (\Add1~53  & VCC)) # (!dcifimemload_15 & (!\Add1~53 )))) # (!\tempReg[29]~54_combout  & ((dcifimemload_15 & (!\Add1~53 )) # (!dcifimemload_15 & ((\Add1~53 ) # (GND)))))
// \Add1~55  = CARRY((\tempReg[29]~54_combout  & (!dcifimemload_15 & !\Add1~53 )) # (!\tempReg[29]~54_combout  & ((!\Add1~53 ) # (!dcifimemload_15))))

	.dataa(\tempReg[29]~54_combout ),
	.datab(dcifimemload_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~53 ),
	.combout(\Add1~54_combout ),
	.cout(\Add1~55 ));
// synopsys translate_off
defparam \Add1~54 .lut_mask = 16'h9617;
defparam \Add1~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N18
cycloneive_lcell_comb \pcif.imemaddr[31]~14 (
// Equation(s):
// \pcif.imemaddr[31]~14_combout  = cuifJmpSel_1 $ (((Equal22 & (!dcifimemload_28 & dcifimemload_27))))

	.dataa(Equal2),
	.datab(dcifimemload_28),
	.datac(dcifimemload_27),
	.datad(cuifJmpSel_1),
	.cin(gnd),
	.combout(\pcif.imemaddr[31]~14_combout ),
	.cout());
// synopsys translate_off
defparam \pcif.imemaddr[31]~14 .lut_mask = 16'hDF20;
defparam \pcif.imemaddr[31]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N30
cycloneive_lcell_comb \pcif.imemaddr[29]~1 (
// Equation(s):
// \pcif.imemaddr[29]~1_combout  = (\pcif.imemaddr[31]~14_combout  & ((Mux2))) # (!\pcif.imemaddr[31]~14_combout  & (\Add1~54_combout ))

	.dataa(\Add1~54_combout ),
	.datab(\pcif.imemaddr[31]~14_combout ),
	.datac(gnd),
	.datad(Mux2),
	.cin(gnd),
	.combout(\pcif.imemaddr[29]~1_combout ),
	.cout());
// synopsys translate_off
defparam \pcif.imemaddr[29]~1 .lut_mask = 16'hEE22;
defparam \pcif.imemaddr[29]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N24
cycloneive_lcell_comb \tempReg[29]~54 (
// Equation(s):
// \tempReg[29]~54_combout  = (pcifimemaddr_29 & (!\tempReg[28]~53 )) # (!pcifimemaddr_29 & ((\tempReg[28]~53 ) # (GND)))
// \tempReg[29]~55  = CARRY((!\tempReg[28]~53 ) # (!pcifimemaddr_29))

	.dataa(pcifimemaddr_29),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[28]~53 ),
	.combout(\tempReg[29]~54_combout ),
	.cout(\tempReg[29]~55 ));
// synopsys translate_off
defparam \tempReg[29]~54 .lut_mask = 16'h5A5F;
defparam \tempReg[29]~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N30
cycloneive_lcell_comb \pcif.imemaddr[31]~10 (
// Equation(s):
// \pcif.imemaddr[31]~10_combout  = (\pcif.imemaddr[31]~9_combout  & (cuifJmpSel_0 & !cuifJmpSel_1)) # (!\pcif.imemaddr[31]~9_combout  & ((cuifJmpSel_0) # (!cuifJmpSel_1)))

	.dataa(\pcif.imemaddr[31]~9_combout ),
	.datab(cuifJmpSel_0),
	.datac(gnd),
	.datad(cuifJmpSel_1),
	.cin(gnd),
	.combout(\pcif.imemaddr[31]~10_combout ),
	.cout());
// synopsys translate_off
defparam \pcif.imemaddr[31]~10 .lut_mask = 16'h44DD;
defparam \pcif.imemaddr[31]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N24
cycloneive_lcell_comb \pcif.imemaddr[31]~15 (
// Equation(s):
// \pcif.imemaddr[31]~15_combout  = (!Selector18 & (Equal102 & (Equal101 & Equal10)))

	.dataa(Selector18),
	.datab(Equal102),
	.datac(Equal101),
	.datad(Equal10),
	.cin(gnd),
	.combout(\pcif.imemaddr[31]~15_combout ),
	.cout());
// synopsys translate_off
defparam \pcif.imemaddr[31]~15 .lut_mask = 16'h4000;
defparam \pcif.imemaddr[31]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N10
cycloneive_lcell_comb \pcif.imemaddr[31]~16 (
// Equation(s):
// \pcif.imemaddr[31]~16_combout  = (!Selector20 & (!Selector21 & (!Selector19 & \pcif.imemaddr[31]~15_combout )))

	.dataa(Selector20),
	.datab(Selector21),
	.datac(Selector19),
	.datad(\pcif.imemaddr[31]~15_combout ),
	.cin(gnd),
	.combout(\pcif.imemaddr[31]~16_combout ),
	.cout());
// synopsys translate_off
defparam \pcif.imemaddr[31]~16 .lut_mask = 16'h0100;
defparam \pcif.imemaddr[31]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N18
cycloneive_lcell_comb \pcif.imemaddr[31]~11 (
// Equation(s):
// \pcif.imemaddr[31]~11_combout  = (Equal22 & (\pcif.imemaddr[31]~16_combout  $ (((dcifimemload_262) # (dcifimemload_261)))))

	.dataa(Equal2),
	.datab(dcifimemload_261),
	.datac(dcifimemload_26),
	.datad(\pcif.imemaddr[31]~16_combout ),
	.cin(gnd),
	.combout(\pcif.imemaddr[31]~11_combout ),
	.cout());
// synopsys translate_off
defparam \pcif.imemaddr[31]~11 .lut_mask = 16'h02A8;
defparam \pcif.imemaddr[31]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N28
cycloneive_lcell_comb \pcif.imemaddr[31]~12 (
// Equation(s):
// \pcif.imemaddr[31]~12_combout  = (\pcif.imemaddr[31]~10_combout ) # ((!\pcif.imemaddr[31]~14_combout  & ((!\pcif.imemaddr[31]~11_combout ) # (!Equal0))))

	.dataa(Equal0),
	.datab(\pcif.imemaddr[31]~14_combout ),
	.datac(\pcif.imemaddr[31]~10_combout ),
	.datad(\pcif.imemaddr[31]~11_combout ),
	.cin(gnd),
	.combout(\pcif.imemaddr[31]~12_combout ),
	.cout());
// synopsys translate_off
defparam \pcif.imemaddr[31]~12 .lut_mask = 16'hF1F3;
defparam \pcif.imemaddr[31]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N20
cycloneive_lcell_comb \pcif.imemaddr[31]~13 (
// Equation(s):
// \pcif.imemaddr[31]~13_combout  = (!ruifdmemWEN & (always1 & (!\dpif.halt~_Duplicate_1_q  & !ruifdmemREN)))

	.dataa(ruifdmemWEN),
	.datab(always1),
	.datac(dpifhalt),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(\pcif.imemaddr[31]~13_combout ),
	.cout());
// synopsys translate_off
defparam \pcif.imemaddr[31]~13 .lut_mask = 16'h0004;
defparam \pcif.imemaddr[31]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N24
cycloneive_lcell_comb \pcif.imemaddr[28]~0 (
// Equation(s):
// \pcif.imemaddr[28]~0_combout  = (\pcif.imemaddr[31]~14_combout  & (Mux3)) # (!\pcif.imemaddr[31]~14_combout  & ((\Add1~52_combout )))

	.dataa(Mux3),
	.datab(\pcif.imemaddr[31]~14_combout ),
	.datac(gnd),
	.datad(\Add1~52_combout ),
	.cin(gnd),
	.combout(\pcif.imemaddr[28]~0_combout ),
	.cout());
// synopsys translate_off
defparam \pcif.imemaddr[28]~0 .lut_mask = 16'hBB88;
defparam \pcif.imemaddr[28]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N26
cycloneive_lcell_comb \tempReg[30]~56 (
// Equation(s):
// \tempReg[30]~56_combout  = (pcifimemaddr_30 & (\tempReg[29]~55  $ (GND))) # (!pcifimemaddr_30 & (!\tempReg[29]~55  & VCC))
// \tempReg[30]~57  = CARRY((pcifimemaddr_30 & !\tempReg[29]~55 ))

	.dataa(gnd),
	.datab(pcifimemaddr_30),
	.datac(gnd),
	.datad(vcc),
	.cin(\tempReg[29]~55 ),
	.combout(\tempReg[30]~56_combout ),
	.cout(\tempReg[30]~57 ));
// synopsys translate_off
defparam \tempReg[30]~56 .lut_mask = 16'hC30C;
defparam \tempReg[30]~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N26
cycloneive_lcell_comb \Add1~56 (
// Equation(s):
// \Add1~56_combout  = ((dcifimemload_15 $ (\tempReg[30]~56_combout  $ (!\Add1~55 )))) # (GND)
// \Add1~57  = CARRY((dcifimemload_15 & ((\tempReg[30]~56_combout ) # (!\Add1~55 ))) # (!dcifimemload_15 & (\tempReg[30]~56_combout  & !\Add1~55 )))

	.dataa(dcifimemload_15),
	.datab(\tempReg[30]~56_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~55 ),
	.combout(\Add1~56_combout ),
	.cout(\Add1~57 ));
// synopsys translate_off
defparam \Add1~56 .lut_mask = 16'h698E;
defparam \Add1~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X50_Y36_N28
cycloneive_lcell_comb \Add1~58 (
// Equation(s):
// \Add1~58_combout  = \tempReg[31]~58_combout  $ (\Add1~57  $ (dcifimemload_15))

	.dataa(\tempReg[31]~58_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(dcifimemload_15),
	.cin(\Add1~57 ),
	.combout(\Add1~58_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~58 .lut_mask = 16'hA55A;
defparam \Add1~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N8
cycloneive_lcell_comb \pcif.imemaddr[31]~3 (
// Equation(s):
// \pcif.imemaddr[31]~3_combout  = (\pcif.imemaddr[31]~14_combout  & (Mux0)) # (!\pcif.imemaddr[31]~14_combout  & ((\Add1~58_combout )))

	.dataa(Mux0),
	.datab(\pcif.imemaddr[31]~14_combout ),
	.datac(gnd),
	.datad(\Add1~58_combout ),
	.cin(gnd),
	.combout(\pcif.imemaddr[31]~3_combout ),
	.cout());
// synopsys translate_off
defparam \pcif.imemaddr[31]~3 .lut_mask = 16'hBB88;
defparam \pcif.imemaddr[31]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y36_N28
cycloneive_lcell_comb \tempReg[31]~58 (
// Equation(s):
// \tempReg[31]~58_combout  = \tempReg[30]~57  $ (pcifimemaddr_31)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(pcifimemaddr_31),
	.cin(\tempReg[30]~57 ),
	.combout(\tempReg[31]~58_combout ),
	.cout());
// synopsys translate_off
defparam \tempReg[31]~58 .lut_mask = 16'h0FF0;
defparam \tempReg[31]~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N30
cycloneive_lcell_comb \pcif.imemaddr[30]~2 (
// Equation(s):
// \pcif.imemaddr[30]~2_combout  = (\pcif.imemaddr[31]~14_combout  & (Mux1)) # (!\pcif.imemaddr[31]~14_combout  & ((\Add1~56_combout )))

	.dataa(Mux1),
	.datab(\pcif.imemaddr[31]~14_combout ),
	.datac(gnd),
	.datad(\Add1~56_combout ),
	.cin(gnd),
	.combout(\pcif.imemaddr[30]~2_combout ),
	.cout());
// synopsys translate_off
defparam \pcif.imemaddr[30]~2 .lut_mask = 16'hBB88;
defparam \pcif.imemaddr[30]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N20
cycloneive_lcell_comb \haltReg~0 (
// Equation(s):
// \haltReg~0_combout  = (Mux30 & ((cuifJmpSel_1) # (!cuifJmpSel_0)))

	.dataa(cuifJmpSel_1),
	.datab(cuifJmpSel_0),
	.datac(Mux30),
	.datad(gnd),
	.cin(gnd),
	.combout(\haltReg~0_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg~0 .lut_mask = 16'hB0B0;
defparam \haltReg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N22
cycloneive_lcell_comb \pcif.imemaddr[1]~8 (
// Equation(s):
// \pcif.imemaddr[1]~8_combout  = (\pcif.imemaddr[31]~13_combout  & (cuifJmpSel_1 $ (cuifJmpSel_0)))

	.dataa(cuifJmpSel_1),
	.datab(cuifJmpSel_0),
	.datac(\pcif.imemaddr[31]~13_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\pcif.imemaddr[1]~8_combout ),
	.cout());
// synopsys translate_off
defparam \pcif.imemaddr[1]~8 .lut_mask = 16'h6060;
defparam \pcif.imemaddr[1]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y36_N0
cycloneive_lcell_comb \haltReg~1 (
// Equation(s):
// \haltReg~1_combout  = (Mux31 & ((cuifJmpSel_1) # (!cuifJmpSel_0)))

	.dataa(gnd),
	.datab(cuifJmpSel_0),
	.datac(cuifJmpSel_1),
	.datad(Mux31),
	.cin(gnd),
	.combout(\haltReg~1_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg~1 .lut_mask = 16'hF300;
defparam \haltReg~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N16
cycloneive_lcell_comb \haltReg[3]~2 (
// Equation(s):
// \haltReg[3]~2_combout  = (\pcif.imemaddr[31]~14_combout  & (((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & ((\pcif.imemaddr[31]~12_combout  & ((\tempReg[3]~2_combout ))) # (!\pcif.imemaddr[31]~12_combout  & (\Add1~2_combout ))))

	.dataa(\Add1~2_combout ),
	.datab(\tempReg[3]~2_combout ),
	.datac(\pcif.imemaddr[31]~14_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[3]~2_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[3]~2 .lut_mask = 16'hFC0A;
defparam \haltReg[3]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N28
cycloneive_lcell_comb \haltReg[3]~3 (
// Equation(s):
// \haltReg[3]~3_combout  = (\pcif.imemaddr[31]~14_combout  & ((\haltReg[3]~2_combout  & (dcifimemload_1)) # (!\haltReg[3]~2_combout  & ((Mux28))))) # (!\pcif.imemaddr[31]~14_combout  & (((\haltReg[3]~2_combout ))))

	.dataa(dcifimemload_1),
	.datab(Mux28),
	.datac(\pcif.imemaddr[31]~14_combout ),
	.datad(\haltReg[3]~2_combout ),
	.cin(gnd),
	.combout(\haltReg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[3]~3 .lut_mask = 16'hAFC0;
defparam \haltReg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N14
cycloneive_lcell_comb \haltReg[2]~4 (
// Equation(s):
// \haltReg[2]~4_combout  = (\pcif.imemaddr[31]~14_combout  & (((Mux29) # (\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & (\Add1~0_combout  & ((!\pcif.imemaddr[31]~12_combout ))))

	.dataa(\Add1~0_combout ),
	.datab(Mux29),
	.datac(\pcif.imemaddr[31]~14_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[2]~4_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[2]~4 .lut_mask = 16'hF0CA;
defparam \haltReg[2]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N6
cycloneive_lcell_comb \haltReg[2]~5 (
// Equation(s):
// \haltReg[2]~5_combout  = (\haltReg[2]~4_combout  & (((dcifimemload_0) # (!\pcif.imemaddr[31]~12_combout )))) # (!\haltReg[2]~4_combout  & (\tempReg[2]~0_combout  & ((\pcif.imemaddr[31]~12_combout ))))

	.dataa(\tempReg[2]~0_combout ),
	.datab(dcifimemload_0),
	.datac(\haltReg[2]~4_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[2]~5_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[2]~5 .lut_mask = 16'hCAF0;
defparam \haltReg[2]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N12
cycloneive_lcell_comb \haltReg[5]~6 (
// Equation(s):
// \haltReg[5]~6_combout  = (\pcif.imemaddr[31]~14_combout  & (((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & ((\pcif.imemaddr[31]~12_combout  & (\tempReg[5]~6_combout )) # (!\pcif.imemaddr[31]~12_combout  & ((\Add1~6_combout )))))

	.dataa(\tempReg[5]~6_combout ),
	.datab(\Add1~6_combout ),
	.datac(\pcif.imemaddr[31]~14_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[5]~6_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[5]~6 .lut_mask = 16'hFA0C;
defparam \haltReg[5]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N4
cycloneive_lcell_comb \haltReg[5]~7 (
// Equation(s):
// \haltReg[5]~7_combout  = (\pcif.imemaddr[31]~14_combout  & ((\haltReg[5]~6_combout  & ((dcifimemload_3))) # (!\haltReg[5]~6_combout  & (Mux26)))) # (!\pcif.imemaddr[31]~14_combout  & (((\haltReg[5]~6_combout ))))

	.dataa(Mux26),
	.datab(dcifimemload_3),
	.datac(\pcif.imemaddr[31]~14_combout ),
	.datad(\haltReg[5]~6_combout ),
	.cin(gnd),
	.combout(\haltReg[5]~7_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[5]~7 .lut_mask = 16'hCFA0;
defparam \haltReg[5]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N10
cycloneive_lcell_comb \haltReg[4]~8 (
// Equation(s):
// \haltReg[4]~8_combout  = (\pcif.imemaddr[31]~14_combout  & ((Mux27) # ((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & (((\Add1~4_combout  & !\pcif.imemaddr[31]~12_combout ))))

	.dataa(Mux27),
	.datab(\pcif.imemaddr[31]~14_combout ),
	.datac(\Add1~4_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[4]~8_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[4]~8 .lut_mask = 16'hCCB8;
defparam \haltReg[4]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N20
cycloneive_lcell_comb \haltReg[4]~9 (
// Equation(s):
// \haltReg[4]~9_combout  = (\pcif.imemaddr[31]~12_combout  & ((\haltReg[4]~8_combout  & (dcifimemload_2)) # (!\haltReg[4]~8_combout  & ((\tempReg[4]~4_combout ))))) # (!\pcif.imemaddr[31]~12_combout  & (((\haltReg[4]~8_combout ))))

	.dataa(dcifimemload_2),
	.datab(\pcif.imemaddr[31]~12_combout ),
	.datac(\tempReg[4]~4_combout ),
	.datad(\haltReg[4]~8_combout ),
	.cin(gnd),
	.combout(\haltReg[4]~9_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[4]~9 .lut_mask = 16'hBBC0;
defparam \haltReg[4]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N4
cycloneive_lcell_comb \haltReg[7]~10 (
// Equation(s):
// \haltReg[7]~10_combout  = (\pcif.imemaddr[31]~14_combout  & (((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & ((\pcif.imemaddr[31]~12_combout  & (\tempReg[7]~10_combout )) # (!\pcif.imemaddr[31]~12_combout  & ((\Add1~10_combout 
// )))))

	.dataa(\tempReg[7]~10_combout ),
	.datab(\pcif.imemaddr[31]~14_combout ),
	.datac(\Add1~10_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[7]~10_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[7]~10 .lut_mask = 16'hEE30;
defparam \haltReg[7]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y35_N30
cycloneive_lcell_comb \haltReg[7]~11 (
// Equation(s):
// \haltReg[7]~11_combout  = (\pcif.imemaddr[31]~14_combout  & ((\haltReg[7]~10_combout  & ((dcifimemload_5))) # (!\haltReg[7]~10_combout  & (Mux24)))) # (!\pcif.imemaddr[31]~14_combout  & (((\haltReg[7]~10_combout ))))

	.dataa(Mux24),
	.datab(\pcif.imemaddr[31]~14_combout ),
	.datac(\haltReg[7]~10_combout ),
	.datad(dcifimemload_5),
	.cin(gnd),
	.combout(\haltReg[7]~11_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[7]~11 .lut_mask = 16'hF838;
defparam \haltReg[7]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N22
cycloneive_lcell_comb \haltReg[6]~12 (
// Equation(s):
// \haltReg[6]~12_combout  = (\pcif.imemaddr[31]~14_combout  & (((Mux25) # (\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & (\Add1~8_combout  & ((!\pcif.imemaddr[31]~12_combout ))))

	.dataa(\Add1~8_combout ),
	.datab(Mux25),
	.datac(\pcif.imemaddr[31]~14_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[6]~12_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[6]~12 .lut_mask = 16'hF0CA;
defparam \haltReg[6]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y36_N18
cycloneive_lcell_comb \haltReg[6]~13 (
// Equation(s):
// \haltReg[6]~13_combout  = (\haltReg[6]~12_combout  & ((dcifimemload_4) # ((!\pcif.imemaddr[31]~12_combout )))) # (!\haltReg[6]~12_combout  & (((\tempReg[6]~8_combout  & \pcif.imemaddr[31]~12_combout ))))

	.dataa(dcifimemload_4),
	.datab(\tempReg[6]~8_combout ),
	.datac(\haltReg[6]~12_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[6]~13_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[6]~13 .lut_mask = 16'hACF0;
defparam \haltReg[6]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N6
cycloneive_lcell_comb \haltReg[9]~14 (
// Equation(s):
// \haltReg[9]~14_combout  = (\pcif.imemaddr[31]~14_combout  & (((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & ((\pcif.imemaddr[31]~12_combout  & ((\tempReg[9]~14_combout ))) # (!\pcif.imemaddr[31]~12_combout  & (\Add1~14_combout 
// ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(\Add1~14_combout ),
	.datac(\tempReg[9]~14_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[9]~14_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[9]~14 .lut_mask = 16'hFA44;
defparam \haltReg[9]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N8
cycloneive_lcell_comb \haltReg[9]~15 (
// Equation(s):
// \haltReg[9]~15_combout  = (\pcif.imemaddr[31]~14_combout  & ((\haltReg[9]~14_combout  & (dcifimemload_7)) # (!\haltReg[9]~14_combout  & ((Mux22))))) # (!\pcif.imemaddr[31]~14_combout  & (((\haltReg[9]~14_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(dcifimemload_7),
	.datac(Mux22),
	.datad(\haltReg[9]~14_combout ),
	.cin(gnd),
	.combout(\haltReg[9]~15_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[9]~15 .lut_mask = 16'hDDA0;
defparam \haltReg[9]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N24
cycloneive_lcell_comb \haltReg[8]~16 (
// Equation(s):
// \haltReg[8]~16_combout  = (\pcif.imemaddr[31]~14_combout  & (((Mux23) # (\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & (\Add1~12_combout  & ((!\pcif.imemaddr[31]~12_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(\Add1~12_combout ),
	.datac(Mux23),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[8]~16_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[8]~16 .lut_mask = 16'hAAE4;
defparam \haltReg[8]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N26
cycloneive_lcell_comb \haltReg[8]~17 (
// Equation(s):
// \haltReg[8]~17_combout  = (\pcif.imemaddr[31]~12_combout  & ((\haltReg[8]~16_combout  & (dcifimemload_6)) # (!\haltReg[8]~16_combout  & ((\tempReg[8]~12_combout ))))) # (!\pcif.imemaddr[31]~12_combout  & (((\haltReg[8]~16_combout ))))

	.dataa(dcifimemload_6),
	.datab(\pcif.imemaddr[31]~12_combout ),
	.datac(\tempReg[8]~12_combout ),
	.datad(\haltReg[8]~16_combout ),
	.cin(gnd),
	.combout(\haltReg[8]~17_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[8]~17 .lut_mask = 16'hBBC0;
defparam \haltReg[8]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N2
cycloneive_lcell_comb \haltReg[11]~18 (
// Equation(s):
// \haltReg[11]~18_combout  = (\pcif.imemaddr[31]~14_combout  & (((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & ((\pcif.imemaddr[31]~12_combout  & ((\tempReg[11]~18_combout ))) # (!\pcif.imemaddr[31]~12_combout  & (\Add1~18_combout 
// ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(\Add1~18_combout ),
	.datac(\tempReg[11]~18_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[11]~18_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[11]~18 .lut_mask = 16'hFA44;
defparam \haltReg[11]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N12
cycloneive_lcell_comb \haltReg[11]~19 (
// Equation(s):
// \haltReg[11]~19_combout  = (\pcif.imemaddr[31]~14_combout  & ((\haltReg[11]~18_combout  & (dcifimemload_9)) # (!\haltReg[11]~18_combout  & ((Mux20))))) # (!\pcif.imemaddr[31]~14_combout  & (((\haltReg[11]~18_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(dcifimemload_9),
	.datac(Mux20),
	.datad(\haltReg[11]~18_combout ),
	.cin(gnd),
	.combout(\haltReg[11]~19_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[11]~19 .lut_mask = 16'hDDA0;
defparam \haltReg[11]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N28
cycloneive_lcell_comb \haltReg[10]~20 (
// Equation(s):
// \haltReg[10]~20_combout  = (\pcif.imemaddr[31]~14_combout  & (((Mux21) # (\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & (\Add1~16_combout  & ((!\pcif.imemaddr[31]~12_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(\Add1~16_combout ),
	.datac(Mux21),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[10]~20_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[10]~20 .lut_mask = 16'hAAE4;
defparam \haltReg[10]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N30
cycloneive_lcell_comb \haltReg[10]~21 (
// Equation(s):
// \haltReg[10]~21_combout  = (\pcif.imemaddr[31]~12_combout  & ((\haltReg[10]~20_combout  & (dcifimemload_8)) # (!\haltReg[10]~20_combout  & ((\tempReg[10]~16_combout ))))) # (!\pcif.imemaddr[31]~12_combout  & (((\haltReg[10]~20_combout ))))

	.dataa(dcifimemload_8),
	.datab(\pcif.imemaddr[31]~12_combout ),
	.datac(\tempReg[10]~16_combout ),
	.datad(\haltReg[10]~20_combout ),
	.cin(gnd),
	.combout(\haltReg[10]~21_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[10]~21 .lut_mask = 16'hBBC0;
defparam \haltReg[10]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N10
cycloneive_lcell_comb \haltReg[13]~22 (
// Equation(s):
// \haltReg[13]~22_combout  = (\pcif.imemaddr[31]~14_combout  & (((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & ((\pcif.imemaddr[31]~12_combout  & ((\tempReg[13]~22_combout ))) # (!\pcif.imemaddr[31]~12_combout  & (\Add1~22_combout 
// ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(\Add1~22_combout ),
	.datac(\tempReg[13]~22_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[13]~22_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[13]~22 .lut_mask = 16'hFA44;
defparam \haltReg[13]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N4
cycloneive_lcell_comb \haltReg[13]~23 (
// Equation(s):
// \haltReg[13]~23_combout  = (\pcif.imemaddr[31]~14_combout  & ((\haltReg[13]~22_combout  & (dcifimemload_11)) # (!\haltReg[13]~22_combout  & ((Mux18))))) # (!\pcif.imemaddr[31]~14_combout  & (((\haltReg[13]~22_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(dcifimemload_11),
	.datac(Mux18),
	.datad(\haltReg[13]~22_combout ),
	.cin(gnd),
	.combout(\haltReg[13]~23_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[13]~23 .lut_mask = 16'hDDA0;
defparam \haltReg[13]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N16
cycloneive_lcell_comb \haltReg[12]~24 (
// Equation(s):
// \haltReg[12]~24_combout  = (\pcif.imemaddr[31]~14_combout  & ((Mux19) # ((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & (((\Add1~20_combout  & !\pcif.imemaddr[31]~12_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(Mux19),
	.datac(\Add1~20_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[12]~24_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[12]~24 .lut_mask = 16'hAAD8;
defparam \haltReg[12]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N22
cycloneive_lcell_comb \haltReg[12]~25 (
// Equation(s):
// \haltReg[12]~25_combout  = (\pcif.imemaddr[31]~12_combout  & ((\haltReg[12]~24_combout  & ((dcifimemload_10))) # (!\haltReg[12]~24_combout  & (\tempReg[12]~20_combout )))) # (!\pcif.imemaddr[31]~12_combout  & (((\haltReg[12]~24_combout ))))

	.dataa(\tempReg[12]~20_combout ),
	.datab(\pcif.imemaddr[31]~12_combout ),
	.datac(dcifimemload_10),
	.datad(\haltReg[12]~24_combout ),
	.cin(gnd),
	.combout(\haltReg[12]~25_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[12]~25 .lut_mask = 16'hF388;
defparam \haltReg[12]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N10
cycloneive_lcell_comb \haltReg[15]~26 (
// Equation(s):
// \haltReg[15]~26_combout  = (\pcif.imemaddr[31]~14_combout  & (((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & ((\pcif.imemaddr[31]~12_combout  & (\tempReg[15]~26_combout )) # (!\pcif.imemaddr[31]~12_combout  & ((\Add1~26_combout 
// )))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(\tempReg[15]~26_combout ),
	.datac(\Add1~26_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[15]~26_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[15]~26 .lut_mask = 16'hEE50;
defparam \haltReg[15]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N12
cycloneive_lcell_comb \haltReg[15]~27 (
// Equation(s):
// \haltReg[15]~27_combout  = (\pcif.imemaddr[31]~14_combout  & ((\haltReg[15]~26_combout  & (dcifimemload_13)) # (!\haltReg[15]~26_combout  & ((Mux16))))) # (!\pcif.imemaddr[31]~14_combout  & (((\haltReg[15]~26_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(dcifimemload_13),
	.datac(Mux16),
	.datad(\haltReg[15]~26_combout ),
	.cin(gnd),
	.combout(\haltReg[15]~27_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[15]~27 .lut_mask = 16'hDDA0;
defparam \haltReg[15]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N8
cycloneive_lcell_comb \haltReg[14]~28 (
// Equation(s):
// \haltReg[14]~28_combout  = (\pcif.imemaddr[31]~14_combout  & ((Mux17) # ((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & (((\Add1~24_combout  & !\pcif.imemaddr[31]~12_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(Mux17),
	.datac(\Add1~24_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[14]~28_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[14]~28 .lut_mask = 16'hAAD8;
defparam \haltReg[14]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N2
cycloneive_lcell_comb \haltReg[14]~29 (
// Equation(s):
// \haltReg[14]~29_combout  = (\haltReg[14]~28_combout  & ((dcifimemload_12) # ((!\pcif.imemaddr[31]~12_combout )))) # (!\haltReg[14]~28_combout  & (((\tempReg[14]~24_combout  & \pcif.imemaddr[31]~12_combout ))))

	.dataa(dcifimemload_12),
	.datab(\tempReg[14]~24_combout ),
	.datac(\haltReg[14]~28_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[14]~29_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[14]~29 .lut_mask = 16'hACF0;
defparam \haltReg[14]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N18
cycloneive_lcell_comb \haltReg[17]~30 (
// Equation(s):
// \haltReg[17]~30_combout  = (\pcif.imemaddr[31]~14_combout  & (((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & ((\pcif.imemaddr[31]~12_combout  & (\tempReg[17]~30_combout )) # (!\pcif.imemaddr[31]~12_combout  & ((\Add1~30_combout 
// )))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(\tempReg[17]~30_combout ),
	.datac(\Add1~30_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[17]~30_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[17]~30 .lut_mask = 16'hEE50;
defparam \haltReg[17]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N0
cycloneive_lcell_comb \haltReg[17]~31 (
// Equation(s):
// \haltReg[17]~31_combout  = (\pcif.imemaddr[31]~14_combout  & ((\haltReg[17]~30_combout  & (dcifimemload_15)) # (!\haltReg[17]~30_combout  & ((Mux14))))) # (!\pcif.imemaddr[31]~14_combout  & (((\haltReg[17]~30_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(dcifimemload_15),
	.datac(Mux14),
	.datad(\haltReg[17]~30_combout ),
	.cin(gnd),
	.combout(\haltReg[17]~31_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[17]~31 .lut_mask = 16'hDDA0;
defparam \haltReg[17]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N20
cycloneive_lcell_comb \haltReg[16]~32 (
// Equation(s):
// \haltReg[16]~32_combout  = (\pcif.imemaddr[31]~14_combout  & ((Mux15) # ((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & (((\Add1~28_combout  & !\pcif.imemaddr[31]~12_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(Mux15),
	.datac(\Add1~28_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[16]~32_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[16]~32 .lut_mask = 16'hAAD8;
defparam \haltReg[16]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N6
cycloneive_lcell_comb \haltReg[16]~33 (
// Equation(s):
// \haltReg[16]~33_combout  = (\pcif.imemaddr[31]~12_combout  & ((\haltReg[16]~32_combout  & ((dcifimemload_14))) # (!\haltReg[16]~32_combout  & (\tempReg[16]~28_combout )))) # (!\pcif.imemaddr[31]~12_combout  & (((\haltReg[16]~32_combout ))))

	.dataa(\tempReg[16]~28_combout ),
	.datab(\pcif.imemaddr[31]~12_combout ),
	.datac(dcifimemload_14),
	.datad(\haltReg[16]~32_combout ),
	.cin(gnd),
	.combout(\haltReg[16]~33_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[16]~33 .lut_mask = 16'hF388;
defparam \haltReg[16]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N30
cycloneive_lcell_comb \haltReg[19]~34 (
// Equation(s):
// \haltReg[19]~34_combout  = (\pcif.imemaddr[31]~14_combout  & (((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & ((\pcif.imemaddr[31]~12_combout  & ((\tempReg[19]~34_combout ))) # (!\pcif.imemaddr[31]~12_combout  & (\Add1~34_combout 
// ))))

	.dataa(\Add1~34_combout ),
	.datab(\pcif.imemaddr[31]~14_combout ),
	.datac(\tempReg[19]~34_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[19]~34_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[19]~34 .lut_mask = 16'hFC22;
defparam \haltReg[19]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y36_N12
cycloneive_lcell_comb \haltReg[19]~35 (
// Equation(s):
// \haltReg[19]~35_combout  = (\pcif.imemaddr[31]~14_combout  & ((\haltReg[19]~34_combout  & (dcifimemload_17)) # (!\haltReg[19]~34_combout  & ((Mux12))))) # (!\pcif.imemaddr[31]~14_combout  & (((\haltReg[19]~34_combout ))))

	.dataa(dcifimemload_17),
	.datab(\pcif.imemaddr[31]~14_combout ),
	.datac(\haltReg[19]~34_combout ),
	.datad(Mux12),
	.cin(gnd),
	.combout(\haltReg[19]~35_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[19]~35 .lut_mask = 16'hBCB0;
defparam \haltReg[19]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N14
cycloneive_lcell_comb \haltReg[18]~36 (
// Equation(s):
// \haltReg[18]~36_combout  = (\pcif.imemaddr[31]~14_combout  & ((Mux13) # ((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & (((\Add1~32_combout  & !\pcif.imemaddr[31]~12_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(Mux13),
	.datac(\Add1~32_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[18]~36_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[18]~36 .lut_mask = 16'hAAD8;
defparam \haltReg[18]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N28
cycloneive_lcell_comb \haltReg[18]~37 (
// Equation(s):
// \haltReg[18]~37_combout  = (\haltReg[18]~36_combout  & ((dcifimemload_16) # ((!\pcif.imemaddr[31]~12_combout )))) # (!\haltReg[18]~36_combout  & (((\tempReg[18]~32_combout  & \pcif.imemaddr[31]~12_combout ))))

	.dataa(dcifimemload_16),
	.datab(\tempReg[18]~32_combout ),
	.datac(\haltReg[18]~36_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[18]~37_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[18]~37 .lut_mask = 16'hACF0;
defparam \haltReg[18]~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N28
cycloneive_lcell_comb \haltReg[21]~38 (
// Equation(s):
// \haltReg[21]~38_combout  = (\pcif.imemaddr[31]~14_combout  & (((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & ((\pcif.imemaddr[31]~12_combout  & ((\tempReg[21]~38_combout ))) # (!\pcif.imemaddr[31]~12_combout  & (\Add1~38_combout 
// ))))

	.dataa(\Add1~38_combout ),
	.datab(\pcif.imemaddr[31]~14_combout ),
	.datac(\tempReg[21]~38_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[21]~38_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[21]~38 .lut_mask = 16'hFC22;
defparam \haltReg[21]~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N4
cycloneive_lcell_comb \haltReg[21]~39 (
// Equation(s):
// \haltReg[21]~39_combout  = (\pcif.imemaddr[31]~14_combout  & ((\haltReg[21]~38_combout  & ((dcifimemload_19))) # (!\haltReg[21]~38_combout  & (Mux10)))) # (!\pcif.imemaddr[31]~14_combout  & (((\haltReg[21]~38_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(Mux10),
	.datac(dcifimemload_19),
	.datad(\haltReg[21]~38_combout ),
	.cin(gnd),
	.combout(\haltReg[21]~39_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[21]~39 .lut_mask = 16'hF588;
defparam \haltReg[21]~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N4
cycloneive_lcell_comb \haltReg[20]~40 (
// Equation(s):
// \haltReg[20]~40_combout  = (\pcif.imemaddr[31]~14_combout  & ((Mux11) # ((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & (((\Add1~36_combout  & !\pcif.imemaddr[31]~12_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(Mux11),
	.datac(\Add1~36_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[20]~40_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[20]~40 .lut_mask = 16'hAAD8;
defparam \haltReg[20]~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N22
cycloneive_lcell_comb \haltReg[20]~41 (
// Equation(s):
// \haltReg[20]~41_combout  = (\haltReg[20]~40_combout  & (((dcifimemload_18) # (!\pcif.imemaddr[31]~12_combout )))) # (!\haltReg[20]~40_combout  & (\tempReg[20]~36_combout  & ((\pcif.imemaddr[31]~12_combout ))))

	.dataa(\tempReg[20]~36_combout ),
	.datab(dcifimemload_18),
	.datac(\haltReg[20]~40_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[20]~41_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[20]~41 .lut_mask = 16'hCAF0;
defparam \haltReg[20]~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N18
cycloneive_lcell_comb \haltReg[23]~42 (
// Equation(s):
// \haltReg[23]~42_combout  = (\pcif.imemaddr[31]~14_combout  & (((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & ((\pcif.imemaddr[31]~12_combout  & ((\tempReg[23]~42_combout ))) # (!\pcif.imemaddr[31]~12_combout  & (\Add1~42_combout 
// ))))

	.dataa(\Add1~42_combout ),
	.datab(\pcif.imemaddr[31]~14_combout ),
	.datac(\tempReg[23]~42_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[23]~42_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[23]~42 .lut_mask = 16'hFC22;
defparam \haltReg[23]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y35_N26
cycloneive_lcell_comb \haltReg[23]~43 (
// Equation(s):
// \haltReg[23]~43_combout  = (\pcif.imemaddr[31]~14_combout  & ((\haltReg[23]~42_combout  & (dcifimemload_21)) # (!\haltReg[23]~42_combout  & ((Mux8))))) # (!\pcif.imemaddr[31]~14_combout  & (((\haltReg[23]~42_combout ))))

	.dataa(dcifimemload_21),
	.datab(\pcif.imemaddr[31]~14_combout ),
	.datac(Mux8),
	.datad(\haltReg[23]~42_combout ),
	.cin(gnd),
	.combout(\haltReg[23]~43_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[23]~43 .lut_mask = 16'hBBC0;
defparam \haltReg[23]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N26
cycloneive_lcell_comb \haltReg[22]~44 (
// Equation(s):
// \haltReg[22]~44_combout  = (\pcif.imemaddr[31]~14_combout  & ((Mux9) # ((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & (((\Add1~40_combout  & !\pcif.imemaddr[31]~12_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(Mux9),
	.datac(\Add1~40_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[22]~44_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[22]~44 .lut_mask = 16'hAAD8;
defparam \haltReg[22]~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y36_N24
cycloneive_lcell_comb \haltReg[22]~45 (
// Equation(s):
// \haltReg[22]~45_combout  = (\haltReg[22]~44_combout  & (((dcifimemload_20) # (!\pcif.imemaddr[31]~12_combout )))) # (!\haltReg[22]~44_combout  & (\tempReg[22]~40_combout  & ((\pcif.imemaddr[31]~12_combout ))))

	.dataa(\tempReg[22]~40_combout ),
	.datab(dcifimemload_20),
	.datac(\haltReg[22]~44_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[22]~45_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[22]~45 .lut_mask = 16'hCAF0;
defparam \haltReg[22]~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N18
cycloneive_lcell_comb \haltReg[25]~46 (
// Equation(s):
// \haltReg[25]~46_combout  = (\pcif.imemaddr[31]~14_combout  & (((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & ((\pcif.imemaddr[31]~12_combout  & (\tempReg[25]~46_combout )) # (!\pcif.imemaddr[31]~12_combout  & ((\Add1~46_combout 
// )))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(\tempReg[25]~46_combout ),
	.datac(\Add1~46_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[25]~46_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[25]~46 .lut_mask = 16'hEE50;
defparam \haltReg[25]~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y36_N20
cycloneive_lcell_comb \haltReg[25]~47 (
// Equation(s):
// \haltReg[25]~47_combout  = (\pcif.imemaddr[31]~14_combout  & ((\haltReg[25]~46_combout  & ((dcifimemload_23))) # (!\haltReg[25]~46_combout  & (Mux6)))) # (!\pcif.imemaddr[31]~14_combout  & (((\haltReg[25]~46_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(Mux6),
	.datac(dcifimemload_23),
	.datad(\haltReg[25]~46_combout ),
	.cin(gnd),
	.combout(\haltReg[25]~47_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[25]~47 .lut_mask = 16'hF588;
defparam \haltReg[25]~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N6
cycloneive_lcell_comb \haltReg[24]~48 (
// Equation(s):
// \haltReg[24]~48_combout  = (\pcif.imemaddr[31]~14_combout  & ((Mux7) # ((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & (((\Add1~44_combout  & !\pcif.imemaddr[31]~12_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(Mux7),
	.datac(\Add1~44_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[24]~48_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[24]~48 .lut_mask = 16'hAAD8;
defparam \haltReg[24]~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N4
cycloneive_lcell_comb \haltReg[24]~49 (
// Equation(s):
// \haltReg[24]~49_combout  = (\pcif.imemaddr[31]~12_combout  & ((\haltReg[24]~48_combout  & (dcifimemload_22)) # (!\haltReg[24]~48_combout  & ((\tempReg[24]~44_combout ))))) # (!\pcif.imemaddr[31]~12_combout  & (((\haltReg[24]~48_combout ))))

	.dataa(dcifimemload_22),
	.datab(\tempReg[24]~44_combout ),
	.datac(\pcif.imemaddr[31]~12_combout ),
	.datad(\haltReg[24]~48_combout ),
	.cin(gnd),
	.combout(\haltReg[24]~49_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[24]~49 .lut_mask = 16'hAFC0;
defparam \haltReg[24]~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N20
cycloneive_lcell_comb \haltReg[27]~50 (
// Equation(s):
// \haltReg[27]~50_combout  = (\pcif.imemaddr[31]~14_combout  & ((Mux4) # ((\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & (((\Add1~50_combout  & !\pcif.imemaddr[31]~12_combout ))))

	.dataa(\pcif.imemaddr[31]~14_combout ),
	.datab(Mux4),
	.datac(\Add1~50_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[27]~50_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[27]~50 .lut_mask = 16'hAAD8;
defparam \haltReg[27]~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y36_N18
cycloneive_lcell_comb \haltReg[27]~51 (
// Equation(s):
// \haltReg[27]~51_combout  = (\pcif.imemaddr[31]~12_combout  & ((\haltReg[27]~50_combout  & ((dcifimemload_25))) # (!\haltReg[27]~50_combout  & (\tempReg[27]~50_combout )))) # (!\pcif.imemaddr[31]~12_combout  & (((\haltReg[27]~50_combout ))))

	.dataa(\tempReg[27]~50_combout ),
	.datab(dcifimemload_25),
	.datac(\pcif.imemaddr[31]~12_combout ),
	.datad(\haltReg[27]~50_combout ),
	.cin(gnd),
	.combout(\haltReg[27]~51_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[27]~51 .lut_mask = 16'hCFA0;
defparam \haltReg[27]~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N30
cycloneive_lcell_comb \haltReg[26]~52 (
// Equation(s):
// \haltReg[26]~52_combout  = (\pcif.imemaddr[31]~14_combout  & (((Mux5) # (\pcif.imemaddr[31]~12_combout )))) # (!\pcif.imemaddr[31]~14_combout  & (\Add1~48_combout  & ((!\pcif.imemaddr[31]~12_combout ))))

	.dataa(\Add1~48_combout ),
	.datab(\pcif.imemaddr[31]~14_combout ),
	.datac(Mux5),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[26]~52_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[26]~52 .lut_mask = 16'hCCE2;
defparam \haltReg[26]~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N20
cycloneive_lcell_comb \haltReg[26]~53 (
// Equation(s):
// \haltReg[26]~53_combout  = (\haltReg[26]~52_combout  & ((dcifimemload_24) # ((!\pcif.imemaddr[31]~12_combout )))) # (!\haltReg[26]~52_combout  & (((\tempReg[26]~48_combout  & \pcif.imemaddr[31]~12_combout ))))

	.dataa(dcifimemload_24),
	.datab(\tempReg[26]~48_combout ),
	.datac(\haltReg[26]~52_combout ),
	.datad(\pcif.imemaddr[31]~12_combout ),
	.cin(gnd),
	.combout(\haltReg[26]~53_combout ),
	.cout());
// synopsys translate_off
defparam \haltReg[26]~53 .lut_mask = 16'hACF0;
defparam \haltReg[26]~53 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module register_file (
	always1,
	cuifregT_3,
	cuifregT_2,
	cuifregT_0,
	cuifregT_1,
	Mux63,
	Mux631,
	Mux32,
	Mux321,
	Mux33,
	Mux331,
	Mux34,
	Mux341,
	Mux35,
	Mux351,
	Mux36,
	Mux361,
	Mux37,
	Mux371,
	Mux38,
	Mux381,
	Mux39,
	Mux391,
	Mux40,
	Mux401,
	Mux41,
	Mux411,
	Mux42,
	Mux421,
	Mux43,
	Mux431,
	Mux58,
	Mux581,
	Mux44,
	Mux441,
	Mux45,
	Mux451,
	Mux46,
	Mux461,
	Mux47,
	Mux471,
	Mux48,
	Mux481,
	Mux49,
	Mux491,
	Mux50,
	Mux501,
	Mux51,
	Mux511,
	Mux52,
	Mux521,
	Mux53,
	Mux531,
	Mux54,
	Mux541,
	Mux55,
	Mux551,
	Mux56,
	Mux561,
	Mux57,
	Mux571,
	cuifregS_2,
	cuifregS_3,
	cuifregS_0,
	cuifregS_1,
	cuifregS_4,
	Mux29,
	Mux30,
	Mux62,
	Mux621,
	Mux27,
	Mux28,
	Mux61,
	Mux611,
	Mux23,
	Mux24,
	Mux25,
	Mux26,
	Mux60,
	Mux601,
	Mux15,
	Mux16,
	Mux17,
	Mux18,
	Mux19,
	Mux20,
	Mux21,
	Mux22,
	Mux59,
	Mux591,
	Mux0,
	Mux2,
	Mux1,
	Mux3,
	Mux4,
	Mux5,
	Mux6,
	Mux7,
	Mux8,
	Mux9,
	Mux10,
	Mux11,
	Mux12,
	Mux13,
	Mux14,
	Mux31,
	Mux68,
	Mux410,
	Mux210,
	Mux01,
	Mux110,
	WEN,
	Mux310,
	Mux372,
	Mux382,
	Mux392,
	Mux402,
	Mux412,
	Mux422,
	Mux432,
	Mux442,
	Mux452,
	Mux462,
	Mux472,
	Mux482,
	Mux632,
	Mux492,
	Mux502,
	Mux512,
	Mux522,
	Mux532,
	Mux542,
	Mux552,
	Mux562,
	Mux572,
	Mux582,
	Mux592,
	Mux602,
	Mux612,
	Mux622,
	Mux66,
	Mux67,
	Mux64,
	Mux65,
	clk,
	n_rst,
	devpor,
	devclrn,
	devoe);
input 	always1;
input 	cuifregT_3;
input 	cuifregT_2;
input 	cuifregT_0;
input 	cuifregT_1;
output 	Mux63;
output 	Mux631;
output 	Mux32;
output 	Mux321;
output 	Mux33;
output 	Mux331;
output 	Mux34;
output 	Mux341;
output 	Mux35;
output 	Mux351;
output 	Mux36;
output 	Mux361;
output 	Mux37;
output 	Mux371;
output 	Mux38;
output 	Mux381;
output 	Mux39;
output 	Mux391;
output 	Mux40;
output 	Mux401;
output 	Mux41;
output 	Mux411;
output 	Mux42;
output 	Mux421;
output 	Mux43;
output 	Mux431;
output 	Mux58;
output 	Mux581;
output 	Mux44;
output 	Mux441;
output 	Mux45;
output 	Mux451;
output 	Mux46;
output 	Mux461;
output 	Mux47;
output 	Mux471;
output 	Mux48;
output 	Mux481;
output 	Mux49;
output 	Mux491;
output 	Mux50;
output 	Mux501;
output 	Mux51;
output 	Mux511;
output 	Mux52;
output 	Mux521;
output 	Mux53;
output 	Mux531;
output 	Mux54;
output 	Mux541;
output 	Mux55;
output 	Mux551;
output 	Mux56;
output 	Mux561;
output 	Mux57;
output 	Mux571;
input 	cuifregS_2;
input 	cuifregS_3;
input 	cuifregS_0;
input 	cuifregS_1;
input 	cuifregS_4;
output 	Mux29;
output 	Mux30;
output 	Mux62;
output 	Mux621;
output 	Mux27;
output 	Mux28;
output 	Mux61;
output 	Mux611;
output 	Mux23;
output 	Mux24;
output 	Mux25;
output 	Mux26;
output 	Mux60;
output 	Mux601;
output 	Mux15;
output 	Mux16;
output 	Mux17;
output 	Mux18;
output 	Mux19;
output 	Mux20;
output 	Mux21;
output 	Mux22;
output 	Mux59;
output 	Mux591;
output 	Mux0;
output 	Mux2;
output 	Mux1;
output 	Mux3;
output 	Mux4;
output 	Mux5;
output 	Mux6;
output 	Mux7;
output 	Mux8;
output 	Mux9;
output 	Mux10;
output 	Mux11;
output 	Mux12;
output 	Mux13;
output 	Mux14;
output 	Mux31;
input 	Mux68;
input 	Mux410;
input 	Mux210;
input 	Mux01;
input 	Mux110;
input 	WEN;
input 	Mux310;
input 	Mux372;
input 	Mux382;
input 	Mux392;
input 	Mux402;
input 	Mux412;
input 	Mux422;
input 	Mux432;
input 	Mux442;
input 	Mux452;
input 	Mux462;
input 	Mux472;
input 	Mux482;
input 	Mux632;
input 	Mux492;
input 	Mux502;
input 	Mux512;
input 	Mux522;
input 	Mux532;
input 	Mux542;
input 	Mux552;
input 	Mux562;
input 	Mux572;
input 	Mux582;
input 	Mux592;
input 	Mux602;
input 	Mux612;
input 	Mux622;
input 	Mux66;
input 	Mux67;
input 	Mux64;
input 	Mux65;
input 	clk;
input 	n_rst;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \registerArray[9][31]~q ;
wire \registerArray[1][31]~q ;
wire \registerArray[10][30]~q ;
wire \registerArray[6][30]~q ;
wire \registerArray[26][30]~q ;
wire \registerArray[24][29]~q ;
wire \registerArray[20][29]~q ;
wire \registerArray[9][29]~q ;
wire \registerArray[10][29]~q ;
wire \registerArray[5][28]~q ;
wire \Mux35~14_combout ;
wire \registerArray[16][27]~q ;
wire \Mux36~14_combout ;
wire \registerArray[3][26]~q ;
wire \registerArray[23][26]~q ;
wire \registerArray[26][25]~q ;
wire \registerArray[22][25]~q ;
wire \registerArray[20][24]~q ;
wire \registerArray[5][24]~q ;
wire \registerArray[12][24]~q ;
wire \registerArray[26][23]~q ;
wire \registerArray[20][23]~q ;
wire \registerArray[10][21]~q ;
wire \registerArray[26][21]~q ;
wire \registerArray[22][21]~q ;
wire \registerArray[27][21]~q ;
wire \registerArray[10][20]~q ;
wire \registerArray[3][20]~q ;
wire \registerArray[5][5]~q ;
wire \registerArray[11][5]~q ;
wire \registerArray[5][19]~q ;
wire \registerArray[13][19]~q ;
wire \registerArray[24][19]~q ;
wire \registerArray[20][19]~q ;
wire \registerArray[5][18]~q ;
wire \registerArray[3][18]~q ;
wire \registerArray[2][18]~q ;
wire \registerArray[13][18]~q ;
wire \registerArray[26][18]~q ;
wire \registerArray[10][17]~q ;
wire \registerArray[20][17]~q ;
wire \registerArray[21][16]~q ;
wire \registerArray[24][16]~q ;
wire \registerArray[16][16]~q ;
wire \Mux47~4_combout ;
wire \registerArray[23][16]~q ;
wire \registerArray[5][16]~q ;
wire \registerArray[3][16]~q ;
wire \registerArray[9][15]~q ;
wire \registerArray[10][15]~q ;
wire \registerArray[19][15]~q ;
wire \registerArray[10][14]~q ;
wire \registerArray[5][14]~q ;
wire \registerArray[5][13]~q ;
wire \registerArray[24][13]~q ;
wire \registerArray[20][13]~q ;
wire \registerArray[1][12]~q ;
wire \registerArray[21][12]~q ;
wire \registerArray[22][12]~q ;
wire \registerArray[10][10]~q ;
wire \registerArray[3][10]~q ;
wire \registerArray[21][10]~q ;
wire \registerArray[23][10]~q ;
wire \registerArray[16][9]~q ;
wire \Mux54~14_combout ;
wire \registerArray[5][8]~q ;
wire \registerArray[22][8]~q ;
wire \registerArray[26][8]~q ;
wire \registerArray[24][8]~q ;
wire \Mux55~14_combout ;
wire \registerArray[10][7]~q ;
wire \registerArray[3][7]~q ;
wire \registerArray[1][7]~q ;
wire \Mux56~4_combout ;
wire \registerArray[22][7]~q ;
wire \registerArray[6][6]~q ;
wire \registerArray[4][6]~q ;
wire \Mux30~7_combout ;
wire \registerArray[10][1]~q ;
wire \Mux30~10_combout ;
wire \registerArray[17][3]~q ;
wire \registerArray[26][3]~q ;
wire \Mux28~2_combout ;
wire \Mux23~2_combout ;
wire \Mux23~3_combout ;
wire \Mux24~10_combout ;
wire \Mux24~14_combout ;
wire \Mux24~15_combout ;
wire \Mux26~12_combout ;
wire \Mux26~13_combout ;
wire \Mux15~4_combout ;
wire \Mux15~5_combout ;
wire \Mux16~14_combout ;
wire \Mux16~15_combout ;
wire \Mux17~12_combout ;
wire \Mux19~14_combout ;
wire \Mux21~12_combout ;
wire \Mux21~14_combout ;
wire \Mux21~15_combout ;
wire \Mux2~4_combout ;
wire \Mux2~5_combout ;
wire \Mux1~2_combout ;
wire \Mux1~3_combout ;
wire \Mux1~12_combout ;
wire \Mux6~2_combout ;
wire \Mux6~3_combout ;
wire \Mux7~10_combout ;
wire \Mux8~2_combout ;
wire \Mux8~3_combout ;
wire \Mux10~2_combout ;
wire \Mux10~3_combout ;
wire \Mux10~10_combout ;
wire \Mux11~14_combout ;
wire \Mux11~15_combout ;
wire \Mux12~4_combout ;
wire \Mux12~5_combout ;
wire \Mux13~2_combout ;
wire \Mux13~3_combout ;
wire \Mux14~4_combout ;
wire \Mux14~5_combout ;
wire \Mux14~10_combout ;
wire \registerArray[9][31]~feeder_combout ;
wire \registerArray[1][31]~feeder_combout ;
wire \registerArray[6][30]~feeder_combout ;
wire \registerArray[10][29]~feeder_combout ;
wire \registerArray[9][29]~feeder_combout ;
wire \registerArray[20][29]~feeder_combout ;
wire \registerArray[5][28]~feeder_combout ;
wire \registerArray[23][26]~feeder_combout ;
wire \registerArray[3][26]~feeder_combout ;
wire \registerArray[12][24]~feeder_combout ;
wire \registerArray[20][24]~feeder_combout ;
wire \registerArray[20][23]~feeder_combout ;
wire \registerArray[27][21]~feeder_combout ;
wire \registerArray[10][20]~feeder_combout ;
wire \registerArray[5][5]~feeder_combout ;
wire \registerArray[11][5]~feeder_combout ;
wire \registerArray[5][19]~feeder_combout ;
wire \registerArray[20][19]~feeder_combout ;
wire \registerArray[13][19]~feeder_combout ;
wire \registerArray[2][18]~feeder_combout ;
wire \registerArray[13][18]~feeder_combout ;
wire \registerArray[5][18]~feeder_combout ;
wire \registerArray[20][17]~feeder_combout ;
wire \registerArray[23][16]~feeder_combout ;
wire \registerArray[21][16]~feeder_combout ;
wire \registerArray[5][16]~feeder_combout ;
wire \registerArray[3][16]~feeder_combout ;
wire \registerArray[19][15]~feeder_combout ;
wire \registerArray[9][15]~feeder_combout ;
wire \registerArray[10][15]~feeder_combout ;
wire \registerArray[5][14]~feeder_combout ;
wire \registerArray[24][13]~feeder_combout ;
wire \registerArray[20][13]~feeder_combout ;
wire \registerArray[5][13]~feeder_combout ;
wire \registerArray[1][12]~feeder_combout ;
wire \registerArray[22][12]~feeder_combout ;
wire \registerArray[21][12]~feeder_combout ;
wire \registerArray[23][10]~feeder_combout ;
wire \registerArray[3][10]~feeder_combout ;
wire \registerArray[5][8]~feeder_combout ;
wire \registerArray[24][8]~feeder_combout ;
wire \registerArray[3][7]~feeder_combout ;
wire \registerArray[22][7]~feeder_combout ;
wire \registerArray[6][6]~feeder_combout ;
wire \registerArray[17][3]~feeder_combout ;
wire \Decoder0~50_combout ;
wire \Decoder0~68_combout ;
wire \registerArray[27][0]~q ;
wire \Decoder0~71_combout ;
wire \registerArray[31][0]~q ;
wire \Decoder0~54_combout ;
wire \Decoder0~70_combout ;
wire \registerArray[19][0]~q ;
wire \Mux63~7_combout ;
wire \Mux63~8_combout ;
wire \registerArray[25][0]~feeder_combout ;
wire \Decoder0~60_combout ;
wire \registerArray[25][0]~q ;
wire \Decoder0~61_combout ;
wire \registerArray[29][0]~q ;
wire \Decoder0~51_combout ;
wire \Decoder0~53_combout ;
wire \registerArray[17][0]~q ;
wire \Mux63~0_combout ;
wire \Mux63~1_combout ;
wire \registerArray[22][0]~feeder_combout ;
wire \Decoder0~62_combout ;
wire \registerArray[22][0]~q ;
wire \Decoder0~65_combout ;
wire \registerArray[30][0]~q ;
wire \Decoder0~64_combout ;
wire \registerArray[18][0]~q ;
wire \Mux63~2_combout ;
wire \Mux63~3_combout ;
wire \Decoder0~67_combout ;
wire \registerArray[28][0]~q ;
wire \registerArray[24][0]~feeder_combout ;
wire \Decoder0~66_combout ;
wire \registerArray[24][0]~q ;
wire \Decoder0~56_combout ;
wire \registerArray[16][0]~q ;
wire \Mux63~4_combout ;
wire \Mux63~5_combout ;
wire \Mux63~6_combout ;
wire \Decoder0~57_combout ;
wire \Decoder0~75_combout ;
wire \registerArray[11][0]~q ;
wire \Decoder0~72_combout ;
wire \registerArray[9][0]~q ;
wire \registerArray[10][0]~feeder_combout ;
wire \Decoder0~73_combout ;
wire \registerArray[10][0]~q ;
wire \Mux63~10_combout ;
wire \Mux63~11_combout ;
wire \registerArray[3][0]~feeder_combout ;
wire \Decoder0~78_combout ;
wire \registerArray[3][0]~q ;
wire \Decoder0~79_combout ;
wire \registerArray[1][0]~q ;
wire \Mux63~14_combout ;
wire \Decoder0~80_combout ;
wire \registerArray[2][0]~q ;
wire \Mux63~15_combout ;
wire \Decoder0~77_combout ;
wire \registerArray[7][0]~q ;
wire \Decoder0~59_combout ;
wire \registerArray[4][0]~q ;
wire \Mux63~12_combout ;
wire \Mux63~13_combout ;
wire \Mux63~16_combout ;
wire \registerArray[14][0]~feeder_combout ;
wire \Decoder0~81_combout ;
wire \registerArray[14][0]~q ;
wire \Decoder0~84_combout ;
wire \registerArray[15][0]~q ;
wire \Decoder0~82_combout ;
wire \registerArray[13][0]~q ;
wire \Decoder0~83_combout ;
wire \registerArray[12][0]~q ;
wire \Mux63~17_combout ;
wire \Mux63~18_combout ;
wire \Decoder0~69_combout ;
wire \registerArray[23][31]~q ;
wire \registerArray[27][31]~q ;
wire \registerArray[19][31]~q ;
wire \Mux32~7_combout ;
wire \registerArray[31][31]~q ;
wire \Mux32~8_combout ;
wire \registerArray[16][31]~feeder_combout ;
wire \registerArray[16][31]~q ;
wire \Decoder0~55_combout ;
wire \registerArray[20][31]~q ;
wire \Mux32~4_combout ;
wire \registerArray[28][31]~q ;
wire \Mux32~5_combout ;
wire \registerArray[30][31]~q ;
wire \registerArray[18][31]~q ;
wire \Mux32~2_combout ;
wire \Mux32~3_combout ;
wire \Mux32~6_combout ;
wire \registerArray[21][31]~feeder_combout ;
wire \Decoder0~52_combout ;
wire \registerArray[21][31]~q ;
wire \registerArray[25][31]~feeder_combout ;
wire \registerArray[25][31]~q ;
wire \registerArray[17][31]~q ;
wire \Mux32~0_combout ;
wire \registerArray[29][31]~q ;
wire \Mux32~1_combout ;
wire \Decoder0~76_combout ;
wire \registerArray[6][31]~q ;
wire \Decoder0~58_combout ;
wire \registerArray[5][31]~q ;
wire \Mux32~10_combout ;
wire \registerArray[7][31]~q ;
wire \Mux32~11_combout ;
wire \registerArray[14][31]~q ;
wire \registerArray[15][31]~q ;
wire \registerArray[13][31]~q ;
wire \registerArray[12][31]~q ;
wire \Mux32~17_combout ;
wire \Mux32~18_combout ;
wire \Decoder0~74_combout ;
wire \registerArray[8][31]~q ;
wire \Mux32~12_combout ;
wire \registerArray[11][31]~q ;
wire \Mux32~13_combout ;
wire \registerArray[2][31]~q ;
wire \registerArray[3][31]~feeder_combout ;
wire \registerArray[3][31]~q ;
wire \Mux32~14_combout ;
wire \Mux32~15_combout ;
wire \Mux32~16_combout ;
wire \registerArray[7][30]~q ;
wire \registerArray[4][30]~q ;
wire \Mux33~2_combout ;
wire \Mux33~3_combout ;
wire \registerArray[2][30]~q ;
wire \registerArray[1][30]~q ;
wire \Mux33~4_combout ;
wire \Mux33~5_combout ;
wire \Mux33~6_combout ;
wire \registerArray[9][30]~q ;
wire \registerArray[11][30]~q ;
wire \registerArray[8][30]~q ;
wire \Mux33~0_combout ;
wire \Mux33~1_combout ;
wire \registerArray[14][30]~q ;
wire \registerArray[15][30]~q ;
wire \registerArray[12][30]~q ;
wire \Mux33~7_combout ;
wire \Mux33~8_combout ;
wire \registerArray[27][30]~q ;
wire \registerArray[31][30]~q ;
wire \registerArray[19][30]~q ;
wire \Mux33~17_combout ;
wire \Mux33~18_combout ;
wire \registerArray[25][30]~q ;
wire \registerArray[29][30]~q ;
wire \registerArray[21][30]~q ;
wire \registerArray[17][30]~q ;
wire \Mux33~10_combout ;
wire \Mux33~11_combout ;
wire \registerArray[22][30]~q ;
wire \registerArray[30][30]~q ;
wire \registerArray[18][30]~q ;
wire \Mux33~12_combout ;
wire \Mux33~13_combout ;
wire \registerArray[20][30]~feeder_combout ;
wire \registerArray[20][30]~q ;
wire \registerArray[16][30]~feeder_combout ;
wire \registerArray[16][30]~q ;
wire \Mux33~14_combout ;
wire \Mux33~15_combout ;
wire \Mux33~16_combout ;
wire \registerArray[23][29]~q ;
wire \registerArray[27][29]~q ;
wire \registerArray[19][29]~q ;
wire \Mux34~7_combout ;
wire \registerArray[31][29]~q ;
wire \Mux34~8_combout ;
wire \registerArray[21][29]~q ;
wire \registerArray[25][29]~feeder_combout ;
wire \registerArray[25][29]~q ;
wire \registerArray[17][29]~q ;
wire \Mux34~0_combout ;
wire \registerArray[29][29]~q ;
wire \Mux34~1_combout ;
wire \registerArray[28][29]~q ;
wire \registerArray[16][29]~q ;
wire \Mux34~4_combout ;
wire \Mux34~5_combout ;
wire \registerArray[30][29]~q ;
wire \registerArray[22][29]~feeder_combout ;
wire \registerArray[22][29]~q ;
wire \registerArray[18][29]~q ;
wire \Mux34~2_combout ;
wire \Mux34~3_combout ;
wire \Mux34~6_combout ;
wire \registerArray[6][29]~q ;
wire \registerArray[4][29]~q ;
wire \Mux34~10_combout ;
wire \registerArray[7][29]~q ;
wire \Mux34~11_combout ;
wire \registerArray[14][29]~q ;
wire \registerArray[15][29]~q ;
wire \registerArray[13][29]~q ;
wire \registerArray[12][29]~q ;
wire \Mux34~17_combout ;
wire \Mux34~18_combout ;
wire \registerArray[11][29]~q ;
wire \registerArray[8][29]~q ;
wire \Mux34~12_combout ;
wire \Mux34~13_combout ;
wire \registerArray[2][29]~q ;
wire \registerArray[3][29]~feeder_combout ;
wire \registerArray[3][29]~q ;
wire \registerArray[1][29]~q ;
wire \Mux34~14_combout ;
wire \Mux34~15_combout ;
wire \Mux34~16_combout ;
wire \registerArray[9][28]~q ;
wire \registerArray[10][28]~q ;
wire \registerArray[8][28]~q ;
wire \Mux35~0_combout ;
wire \registerArray[11][28]~q ;
wire \Mux35~1_combout ;
wire \registerArray[14][28]~q ;
wire \registerArray[15][28]~q ;
wire \registerArray[13][28]~q ;
wire \registerArray[12][28]~q ;
wire \Mux35~7_combout ;
wire \Mux35~8_combout ;
wire \registerArray[7][28]~q ;
wire \registerArray[4][28]~q ;
wire \Mux35~2_combout ;
wire \Mux35~3_combout ;
wire \registerArray[2][28]~q ;
wire \registerArray[3][28]~feeder_combout ;
wire \registerArray[3][28]~q ;
wire \registerArray[1][28]~q ;
wire \Mux35~4_combout ;
wire \Mux35~5_combout ;
wire \Mux35~6_combout ;
wire \registerArray[23][28]~feeder_combout ;
wire \registerArray[23][28]~q ;
wire \registerArray[19][28]~q ;
wire \Mux35~17_combout ;
wire \registerArray[31][28]~q ;
wire \registerArray[27][28]~feeder_combout ;
wire \registerArray[27][28]~q ;
wire \Mux35~18_combout ;
wire \registerArray[20][28]~q ;
wire \registerArray[28][28]~q ;
wire \Mux35~15_combout ;
wire \Decoder0~63_combout ;
wire \registerArray[26][28]~q ;
wire \registerArray[18][28]~q ;
wire \Mux35~12_combout ;
wire \registerArray[30][28]~q ;
wire \Mux35~13_combout ;
wire \Mux35~16_combout ;
wire \registerArray[29][28]~feeder_combout ;
wire \registerArray[29][28]~q ;
wire \registerArray[25][28]~feeder_combout ;
wire \registerArray[25][28]~q ;
wire \registerArray[21][28]~feeder_combout ;
wire \registerArray[21][28]~q ;
wire \Mux35~10_combout ;
wire \Mux35~11_combout ;
wire \registerArray[5][27]~q ;
wire \registerArray[4][27]~q ;
wire \Mux36~0_combout ;
wire \registerArray[7][27]~q ;
wire \registerArray[6][27]~q ;
wire \Mux36~1_combout ;
wire \registerArray[14][27]~q ;
wire \registerArray[13][27]~q ;
wire \registerArray[12][27]~q ;
wire \Mux36~7_combout ;
wire \registerArray[15][27]~q ;
wire \Mux36~8_combout ;
wire \registerArray[2][27]~q ;
wire \registerArray[3][27]~q ;
wire \registerArray[1][27]~q ;
wire \Mux36~4_combout ;
wire \Mux36~5_combout ;
wire \registerArray[9][27]~q ;
wire \registerArray[11][27]~q ;
wire \registerArray[8][27]~q ;
wire \Mux36~2_combout ;
wire \Mux36~3_combout ;
wire \Mux36~6_combout ;
wire \registerArray[21][27]~feeder_combout ;
wire \registerArray[21][27]~q ;
wire \registerArray[29][27]~q ;
wire \registerArray[25][27]~feeder_combout ;
wire \registerArray[25][27]~q ;
wire \registerArray[17][27]~feeder_combout ;
wire \registerArray[17][27]~q ;
wire \Mux36~10_combout ;
wire \Mux36~11_combout ;
wire \registerArray[18][27]~q ;
wire \Mux36~12_combout ;
wire \registerArray[30][27]~q ;
wire \Mux36~13_combout ;
wire \registerArray[24][27]~q ;
wire \registerArray[28][27]~q ;
wire \Mux36~15_combout ;
wire \Mux36~16_combout ;
wire \registerArray[27][27]~q ;
wire \registerArray[19][27]~q ;
wire \Mux36~17_combout ;
wire \registerArray[23][27]~feeder_combout ;
wire \registerArray[23][27]~q ;
wire \registerArray[31][27]~q ;
wire \Mux36~18_combout ;
wire \registerArray[14][26]~feeder_combout ;
wire \registerArray[14][26]~q ;
wire \registerArray[15][26]~q ;
wire \registerArray[13][26]~feeder_combout ;
wire \registerArray[13][26]~q ;
wire \registerArray[12][26]~q ;
wire \Mux37~7_combout ;
wire \Mux37~8_combout ;
wire \registerArray[6][26]~q ;
wire \registerArray[7][26]~q ;
wire \registerArray[5][26]~feeder_combout ;
wire \registerArray[5][26]~q ;
wire \registerArray[4][26]~q ;
wire \Mux37~2_combout ;
wire \Mux37~3_combout ;
wire \registerArray[2][26]~q ;
wire \registerArray[1][26]~q ;
wire \Mux37~4_combout ;
wire \Mux37~5_combout ;
wire \Mux37~6_combout ;
wire \registerArray[11][26]~q ;
wire \registerArray[9][26]~q ;
wire \registerArray[8][26]~q ;
wire \registerArray[10][26]~q ;
wire \Mux37~0_combout ;
wire \Mux37~1_combout ;
wire \registerArray[25][26]~q ;
wire \registerArray[29][26]~q ;
wire \registerArray[21][26]~q ;
wire \registerArray[17][26]~q ;
wire \Mux37~10_combout ;
wire \Mux37~11_combout ;
wire \registerArray[19][26]~q ;
wire \Mux37~17_combout ;
wire \registerArray[31][26]~q ;
wire \registerArray[27][26]~q ;
wire \Mux37~18_combout ;
wire \registerArray[28][26]~q ;
wire \registerArray[24][26]~feeder_combout ;
wire \registerArray[24][26]~q ;
wire \registerArray[16][26]~q ;
wire \Mux37~14_combout ;
wire \Mux37~15_combout ;
wire \registerArray[22][26]~q ;
wire \registerArray[30][26]~q ;
wire \registerArray[26][26]~q ;
wire \registerArray[18][26]~q ;
wire \Mux37~12_combout ;
wire \Mux37~13_combout ;
wire \Mux37~16_combout ;
wire \registerArray[14][25]~q ;
wire \registerArray[12][25]~q ;
wire \registerArray[13][25]~q ;
wire \Mux38~7_combout ;
wire \registerArray[15][25]~q ;
wire \Mux38~8_combout ;
wire \registerArray[6][25]~q ;
wire \registerArray[7][25]~q ;
wire \registerArray[5][25]~feeder_combout ;
wire \registerArray[5][25]~q ;
wire \registerArray[4][25]~q ;
wire \Mux38~0_combout ;
wire \Mux38~1_combout ;
wire \registerArray[11][25]~q ;
wire \registerArray[8][25]~q ;
wire \Mux38~2_combout ;
wire \Mux38~3_combout ;
wire \registerArray[2][25]~q ;
wire \registerArray[3][25]~q ;
wire \registerArray[1][25]~q ;
wire \Mux38~4_combout ;
wire \Mux38~5_combout ;
wire \Mux38~6_combout ;
wire \registerArray[30][25]~q ;
wire \registerArray[18][25]~q ;
wire \Mux38~12_combout ;
wire \Mux38~13_combout ;
wire \registerArray[28][25]~q ;
wire \registerArray[20][25]~q ;
wire \registerArray[16][25]~q ;
wire \Mux38~14_combout ;
wire \Mux38~15_combout ;
wire \Mux38~16_combout ;
wire \registerArray[23][25]~q ;
wire \registerArray[31][25]~q ;
wire \registerArray[19][25]~q ;
wire \Mux38~17_combout ;
wire \Mux38~18_combout ;
wire \registerArray[21][25]~q ;
wire \registerArray[29][25]~q ;
wire \registerArray[25][25]~q ;
wire \registerArray[17][25]~q ;
wire \Mux38~10_combout ;
wire \Mux38~11_combout ;
wire \registerArray[29][24]~feeder_combout ;
wire \registerArray[29][24]~q ;
wire \registerArray[25][24]~feeder_combout ;
wire \registerArray[25][24]~q ;
wire \registerArray[17][24]~feeder_combout ;
wire \registerArray[17][24]~q ;
wire \registerArray[21][24]~feeder_combout ;
wire \registerArray[21][24]~q ;
wire \Mux39~0_combout ;
wire \Mux39~1_combout ;
wire \registerArray[27][24]~q ;
wire \registerArray[31][24]~q ;
wire \registerArray[19][24]~q ;
wire \Mux39~7_combout ;
wire \Mux39~8_combout ;
wire \registerArray[28][24]~feeder_combout ;
wire \registerArray[28][24]~q ;
wire \registerArray[24][24]~feeder_combout ;
wire \registerArray[24][24]~q ;
wire \Mux39~4_combout ;
wire \Mux39~5_combout ;
wire \registerArray[22][24]~q ;
wire \registerArray[30][24]~q ;
wire \registerArray[18][24]~q ;
wire \Mux39~2_combout ;
wire \Mux39~3_combout ;
wire \Mux39~6_combout ;
wire \registerArray[14][24]~feeder_combout ;
wire \registerArray[14][24]~q ;
wire \registerArray[15][24]~q ;
wire \registerArray[13][24]~q ;
wire \Mux39~17_combout ;
wire \Mux39~18_combout ;
wire \registerArray[9][24]~q ;
wire \registerArray[11][24]~q ;
wire \registerArray[8][24]~q ;
wire \Mux39~10_combout ;
wire \Mux39~11_combout ;
wire \registerArray[6][24]~q ;
wire \registerArray[4][24]~q ;
wire \Mux39~12_combout ;
wire \Mux39~13_combout ;
wire \registerArray[2][24]~q ;
wire \registerArray[1][24]~q ;
wire \Mux39~14_combout ;
wire \Mux39~15_combout ;
wire \Mux39~16_combout ;
wire \registerArray[14][23]~feeder_combout ;
wire \registerArray[14][23]~q ;
wire \registerArray[15][23]~q ;
wire \registerArray[12][23]~q ;
wire \registerArray[13][23]~feeder_combout ;
wire \registerArray[13][23]~q ;
wire \Mux40~7_combout ;
wire \Mux40~8_combout ;
wire \registerArray[6][23]~q ;
wire \registerArray[7][23]~q ;
wire \registerArray[4][23]~q ;
wire \Mux40~0_combout ;
wire \Mux40~1_combout ;
wire \registerArray[2][23]~q ;
wire \registerArray[1][23]~q ;
wire \Mux40~4_combout ;
wire \Mux40~5_combout ;
wire \registerArray[9][23]~q ;
wire \registerArray[11][23]~q ;
wire \registerArray[8][23]~q ;
wire \Mux40~2_combout ;
wire \Mux40~3_combout ;
wire \Mux40~6_combout ;
wire \registerArray[22][23]~q ;
wire \registerArray[18][23]~q ;
wire \Mux40~12_combout ;
wire \registerArray[30][23]~q ;
wire \Mux40~13_combout ;
wire \registerArray[28][23]~q ;
wire \registerArray[16][23]~q ;
wire \Mux40~14_combout ;
wire \Mux40~15_combout ;
wire \Mux40~16_combout ;
wire \registerArray[21][23]~q ;
wire \registerArray[29][23]~q ;
wire \registerArray[17][23]~q ;
wire \registerArray[25][23]~q ;
wire \Mux40~10_combout ;
wire \Mux40~11_combout ;
wire \registerArray[19][23]~feeder_combout ;
wire \registerArray[19][23]~q ;
wire \Mux40~17_combout ;
wire \registerArray[31][23]~q ;
wire \registerArray[23][23]~feeder_combout ;
wire \registerArray[23][23]~q ;
wire \Mux40~18_combout ;
wire \registerArray[14][22]~q ;
wire \registerArray[15][22]~q ;
wire \registerArray[12][22]~q ;
wire \registerArray[13][22]~feeder_combout ;
wire \registerArray[13][22]~q ;
wire \Mux41~7_combout ;
wire \Mux41~8_combout ;
wire \registerArray[9][22]~feeder_combout ;
wire \registerArray[9][22]~q ;
wire \registerArray[11][22]~q ;
wire \registerArray[8][22]~q ;
wire \Mux41~0_combout ;
wire \Mux41~1_combout ;
wire \registerArray[2][22]~q ;
wire \registerArray[1][22]~q ;
wire \Mux41~4_combout ;
wire \Mux41~5_combout ;
wire \registerArray[7][22]~q ;
wire \registerArray[4][22]~q ;
wire \registerArray[5][22]~q ;
wire \Mux41~2_combout ;
wire \Mux41~3_combout ;
wire \Mux41~6_combout ;
wire \registerArray[31][22]~feeder_combout ;
wire \registerArray[31][22]~q ;
wire \registerArray[27][22]~q ;
wire \registerArray[19][22]~q ;
wire \Mux41~17_combout ;
wire \Mux41~18_combout ;
wire \registerArray[25][22]~q ;
wire \registerArray[29][22]~q ;
wire \registerArray[17][22]~q ;
wire \registerArray[21][22]~q ;
wire \Mux41~10_combout ;
wire \Mux41~11_combout ;
wire \registerArray[22][22]~q ;
wire \registerArray[30][22]~q ;
wire \registerArray[26][22]~q ;
wire \registerArray[18][22]~q ;
wire \Mux41~12_combout ;
wire \Mux41~13_combout ;
wire \registerArray[16][22]~q ;
wire \registerArray[24][22]~q ;
wire \Mux41~14_combout ;
wire \registerArray[28][22]~feeder_combout ;
wire \registerArray[28][22]~q ;
wire \Mux41~15_combout ;
wire \Mux41~16_combout ;
wire \registerArray[14][21]~q ;
wire \registerArray[15][21]~q ;
wire \registerArray[12][21]~q ;
wire \registerArray[13][21]~q ;
wire \Mux42~7_combout ;
wire \Mux42~8_combout ;
wire \registerArray[2][21]~q ;
wire \registerArray[1][21]~feeder_combout ;
wire \registerArray[1][21]~q ;
wire \Mux42~4_combout ;
wire \Mux42~5_combout ;
wire \registerArray[9][21]~q ;
wire \registerArray[8][21]~q ;
wire \Mux42~2_combout ;
wire \Mux42~3_combout ;
wire \Mux42~6_combout ;
wire \registerArray[6][21]~feeder_combout ;
wire \registerArray[6][21]~q ;
wire \registerArray[7][21]~q ;
wire \registerArray[4][21]~q ;
wire \Mux42~0_combout ;
wire \Mux42~1_combout ;
wire \registerArray[21][21]~feeder_combout ;
wire \registerArray[21][21]~q ;
wire \registerArray[29][21]~q ;
wire \registerArray[17][21]~feeder_combout ;
wire \registerArray[17][21]~q ;
wire \registerArray[25][21]~feeder_combout ;
wire \registerArray[25][21]~q ;
wire \Mux42~10_combout ;
wire \Mux42~11_combout ;
wire \registerArray[31][21]~feeder_combout ;
wire \registerArray[31][21]~q ;
wire \registerArray[23][21]~q ;
wire \registerArray[19][21]~q ;
wire \Mux42~17_combout ;
wire \Mux42~18_combout ;
wire \registerArray[28][21]~q ;
wire \registerArray[20][21]~q ;
wire \Mux42~14_combout ;
wire \Mux42~15_combout ;
wire \registerArray[30][21]~q ;
wire \registerArray[18][21]~q ;
wire \Mux42~12_combout ;
wire \Mux42~13_combout ;
wire \Mux42~16_combout ;
wire \registerArray[14][20]~q ;
wire \registerArray[15][20]~q ;
wire \registerArray[12][20]~q ;
wire \registerArray[13][20]~q ;
wire \Mux43~7_combout ;
wire \Mux43~8_combout ;
wire \registerArray[11][20]~feeder_combout ;
wire \registerArray[11][20]~q ;
wire \registerArray[9][20]~feeder_combout ;
wire \registerArray[9][20]~q ;
wire \registerArray[8][20]~q ;
wire \Mux43~0_combout ;
wire \Mux43~1_combout ;
wire \registerArray[7][20]~q ;
wire \registerArray[4][20]~q ;
wire \Mux43~2_combout ;
wire \Mux43~3_combout ;
wire \registerArray[2][20]~q ;
wire \registerArray[1][20]~q ;
wire \Mux43~4_combout ;
wire \Mux43~5_combout ;
wire \Mux43~6_combout ;
wire \registerArray[16][20]~feeder_combout ;
wire \registerArray[16][20]~q ;
wire \registerArray[24][20]~q ;
wire \Mux43~14_combout ;
wire \registerArray[28][20]~q ;
wire \Mux43~15_combout ;
wire \registerArray[22][20]~q ;
wire \registerArray[30][20]~q ;
wire \registerArray[26][20]~feeder_combout ;
wire \registerArray[26][20]~q ;
wire \registerArray[18][20]~q ;
wire \Mux43~12_combout ;
wire \Mux43~13_combout ;
wire \Mux43~16_combout ;
wire \registerArray[25][20]~q ;
wire \registerArray[29][20]~q ;
wire \registerArray[17][20]~q ;
wire \Mux43~10_combout ;
wire \Mux43~11_combout ;
wire \registerArray[27][20]~q ;
wire \registerArray[31][20]~q ;
wire \registerArray[19][20]~feeder_combout ;
wire \registerArray[19][20]~q ;
wire \Mux43~17_combout ;
wire \Mux43~18_combout ;
wire \registerArray[14][5]~feeder_combout ;
wire \registerArray[14][5]~q ;
wire \registerArray[15][5]~q ;
wire \registerArray[12][5]~q ;
wire \Mux58~7_combout ;
wire \Mux58~8_combout ;
wire \registerArray[6][5]~feeder_combout ;
wire \registerArray[6][5]~q ;
wire \registerArray[7][5]~q ;
wire \registerArray[4][5]~feeder_combout ;
wire \registerArray[4][5]~q ;
wire \Mux58~0_combout ;
wire \Mux58~1_combout ;
wire \registerArray[3][5]~q ;
wire \Mux58~4_combout ;
wire \Mux58~5_combout ;
wire \registerArray[9][5]~q ;
wire \registerArray[8][5]~q ;
wire \Mux58~2_combout ;
wire \Mux58~3_combout ;
wire \Mux58~6_combout ;
wire \registerArray[23][5]~q ;
wire \registerArray[27][5]~q ;
wire \registerArray[19][5]~q ;
wire \Mux58~17_combout ;
wire \registerArray[31][5]~q ;
wire \Mux58~18_combout ;
wire \registerArray[28][5]~feeder_combout ;
wire \registerArray[28][5]~q ;
wire \registerArray[16][5]~feeder_combout ;
wire \registerArray[16][5]~q ;
wire \registerArray[20][5]~q ;
wire \Mux58~14_combout ;
wire \Mux58~15_combout ;
wire \registerArray[30][5]~q ;
wire \registerArray[18][5]~q ;
wire \Mux58~12_combout ;
wire \Mux58~13_combout ;
wire \Mux58~16_combout ;
wire \registerArray[21][5]~q ;
wire \registerArray[17][5]~q ;
wire \Mux58~10_combout ;
wire \registerArray[29][5]~q ;
wire \Mux58~11_combout ;
wire \registerArray[15][19]~feeder_combout ;
wire \registerArray[15][19]~q ;
wire \registerArray[14][19]~feeder_combout ;
wire \registerArray[14][19]~q ;
wire \registerArray[12][19]~q ;
wire \Mux44~7_combout ;
wire \Mux44~8_combout ;
wire \registerArray[6][19]~q ;
wire \registerArray[7][19]~q ;
wire \registerArray[4][19]~q ;
wire \Mux44~0_combout ;
wire \Mux44~1_combout ;
wire \registerArray[11][19]~q ;
wire \registerArray[8][19]~feeder_combout ;
wire \registerArray[8][19]~q ;
wire \Mux44~2_combout ;
wire \Mux44~3_combout ;
wire \registerArray[2][19]~q ;
wire \registerArray[3][19]~q ;
wire \Mux44~4_combout ;
wire \Mux44~5_combout ;
wire \Mux44~6_combout ;
wire \registerArray[28][19]~q ;
wire \registerArray[16][19]~q ;
wire \Mux44~14_combout ;
wire \Mux44~15_combout ;
wire \registerArray[26][19]~feeder_combout ;
wire \registerArray[26][19]~q ;
wire \registerArray[30][19]~q ;
wire \registerArray[22][19]~feeder_combout ;
wire \registerArray[22][19]~q ;
wire \registerArray[18][19]~q ;
wire \Mux44~12_combout ;
wire \Mux44~13_combout ;
wire \Mux44~16_combout ;
wire \registerArray[23][19]~q ;
wire \registerArray[31][19]~q ;
wire \registerArray[27][19]~q ;
wire \registerArray[19][19]~q ;
wire \Mux44~17_combout ;
wire \Mux44~18_combout ;
wire \registerArray[21][19]~q ;
wire \registerArray[29][19]~q ;
wire \registerArray[25][19]~feeder_combout ;
wire \registerArray[25][19]~q ;
wire \registerArray[17][19]~q ;
wire \Mux44~10_combout ;
wire \Mux44~11_combout ;
wire \registerArray[9][18]~feeder_combout ;
wire \registerArray[9][18]~q ;
wire \registerArray[11][18]~q ;
wire \registerArray[8][18]~q ;
wire \Mux45~0_combout ;
wire \Mux45~1_combout ;
wire \registerArray[14][18]~feeder_combout ;
wire \registerArray[14][18]~q ;
wire \registerArray[15][18]~q ;
wire \registerArray[12][18]~q ;
wire \Mux45~7_combout ;
wire \Mux45~8_combout ;
wire \registerArray[7][18]~q ;
wire \registerArray[4][18]~q ;
wire \Mux45~2_combout ;
wire \Mux45~3_combout ;
wire \registerArray[1][18]~q ;
wire \Mux45~4_combout ;
wire \Mux45~5_combout ;
wire \Mux45~6_combout ;
wire \registerArray[22][18]~q ;
wire \registerArray[30][18]~q ;
wire \registerArray[18][18]~q ;
wire \Mux45~12_combout ;
wire \Mux45~13_combout ;
wire \registerArray[28][18]~q ;
wire \registerArray[24][18]~q ;
wire \registerArray[16][18]~q ;
wire \Mux45~14_combout ;
wire \Mux45~15_combout ;
wire \Mux45~16_combout ;
wire \registerArray[27][18]~feeder_combout ;
wire \registerArray[27][18]~q ;
wire \registerArray[31][18]~q ;
wire \registerArray[19][18]~q ;
wire \Mux45~17_combout ;
wire \Mux45~18_combout ;
wire \registerArray[25][18]~feeder_combout ;
wire \registerArray[25][18]~q ;
wire \registerArray[29][18]~q ;
wire \registerArray[21][18]~feeder_combout ;
wire \registerArray[21][18]~q ;
wire \Mux45~10_combout ;
wire \Mux45~11_combout ;
wire \registerArray[14][17]~feeder_combout ;
wire \registerArray[14][17]~q ;
wire \registerArray[15][17]~q ;
wire \registerArray[12][17]~q ;
wire \Mux46~7_combout ;
wire \Mux46~8_combout ;
wire \registerArray[6][17]~q ;
wire \registerArray[7][17]~q ;
wire \registerArray[5][17]~q ;
wire \Mux46~0_combout ;
wire \Mux46~1_combout ;
wire \registerArray[9][17]~q ;
wire \registerArray[11][17]~q ;
wire \registerArray[8][17]~q ;
wire \Mux46~2_combout ;
wire \Mux46~3_combout ;
wire \registerArray[2][17]~q ;
wire \registerArray[1][17]~q ;
wire \Mux46~4_combout ;
wire \Mux46~5_combout ;
wire \Mux46~6_combout ;
wire \registerArray[24][17]~q ;
wire \registerArray[28][17]~q ;
wire \registerArray[16][17]~q ;
wire \Mux46~14_combout ;
wire \Mux46~15_combout ;
wire \registerArray[30][17]~q ;
wire \registerArray[18][17]~q ;
wire \Mux46~12_combout ;
wire \Mux46~13_combout ;
wire \Mux46~16_combout ;
wire \registerArray[21][17]~q ;
wire \registerArray[29][17]~q ;
wire \registerArray[25][17]~q ;
wire \Mux46~10_combout ;
wire \Mux46~11_combout ;
wire \registerArray[31][17]~q ;
wire \registerArray[23][17]~q ;
wire \registerArray[19][17]~q ;
wire \Mux46~17_combout ;
wire \Mux46~18_combout ;
wire \registerArray[27][16]~feeder_combout ;
wire \registerArray[27][16]~q ;
wire \registerArray[31][16]~q ;
wire \registerArray[19][16]~feeder_combout ;
wire \registerArray[19][16]~q ;
wire \Mux47~7_combout ;
wire \Mux47~8_combout ;
wire \registerArray[29][16]~feeder_combout ;
wire \registerArray[29][16]~q ;
wire \registerArray[25][16]~q ;
wire \registerArray[17][16]~feeder_combout ;
wire \registerArray[17][16]~q ;
wire \Mux47~0_combout ;
wire \Mux47~1_combout ;
wire \registerArray[20][16]~q ;
wire \registerArray[28][16]~q ;
wire \Mux47~5_combout ;
wire \registerArray[30][16]~q ;
wire \registerArray[26][16]~q ;
wire \registerArray[18][16]~q ;
wire \Mux47~2_combout ;
wire \Mux47~3_combout ;
wire \Mux47~6_combout ;
wire \registerArray[14][16]~feeder_combout ;
wire \registerArray[14][16]~q ;
wire \registerArray[15][16]~q ;
wire \registerArray[12][16]~q ;
wire \Mux47~17_combout ;
wire \Mux47~18_combout ;
wire \registerArray[2][16]~q ;
wire \registerArray[1][16]~q ;
wire \Mux47~14_combout ;
wire \Mux47~15_combout ;
wire \registerArray[6][16]~q ;
wire \registerArray[4][16]~q ;
wire \Mux47~12_combout ;
wire \Mux47~13_combout ;
wire \Mux47~16_combout ;
wire \registerArray[9][16]~q ;
wire \registerArray[8][16]~q ;
wire \Mux47~10_combout ;
wire \registerArray[11][16]~q ;
wire \Mux47~11_combout ;
wire \registerArray[6][15]~feeder_combout ;
wire \registerArray[6][15]~q ;
wire \registerArray[7][15]~q ;
wire \registerArray[4][15]~q ;
wire \Mux48~0_combout ;
wire \Mux48~1_combout ;
wire \registerArray[14][15]~feeder_combout ;
wire \registerArray[14][15]~q ;
wire \registerArray[15][15]~q ;
wire \registerArray[12][15]~q ;
wire \Mux48~7_combout ;
wire \Mux48~8_combout ;
wire \registerArray[2][15]~q ;
wire \registerArray[1][15]~q ;
wire \registerArray[3][15]~feeder_combout ;
wire \registerArray[3][15]~q ;
wire \Mux48~4_combout ;
wire \Mux48~5_combout ;
wire \registerArray[11][15]~q ;
wire \registerArray[8][15]~q ;
wire \Mux48~2_combout ;
wire \Mux48~3_combout ;
wire \Mux48~6_combout ;
wire \registerArray[21][15]~q ;
wire \registerArray[29][15]~q ;
wire \registerArray[17][15]~q ;
wire \Mux48~10_combout ;
wire \Mux48~11_combout ;
wire \registerArray[23][15]~feeder_combout ;
wire \registerArray[23][15]~q ;
wire \registerArray[31][15]~q ;
wire \registerArray[27][15]~feeder_combout ;
wire \registerArray[27][15]~q ;
wire \Mux48~17_combout ;
wire \Mux48~18_combout ;
wire \registerArray[28][15]~feeder_combout ;
wire \registerArray[28][15]~q ;
wire \registerArray[16][15]~feeder_combout ;
wire \registerArray[16][15]~q ;
wire \Mux48~14_combout ;
wire \Mux48~15_combout ;
wire \registerArray[26][15]~feeder_combout ;
wire \registerArray[26][15]~q ;
wire \registerArray[30][15]~q ;
wire \registerArray[18][15]~q ;
wire \registerArray[22][15]~q ;
wire \Mux48~12_combout ;
wire \Mux48~13_combout ;
wire \Mux48~16_combout ;
wire \registerArray[12][14]~q ;
wire \Mux49~7_combout ;
wire \registerArray[15][14]~q ;
wire \registerArray[14][14]~feeder_combout ;
wire \registerArray[14][14]~q ;
wire \Mux49~8_combout ;
wire \registerArray[9][14]~q ;
wire \registerArray[11][14]~q ;
wire \registerArray[8][14]~q ;
wire \Mux49~0_combout ;
wire \Mux49~1_combout ;
wire \registerArray[7][14]~q ;
wire \registerArray[4][14]~q ;
wire \Mux49~2_combout ;
wire \Mux49~3_combout ;
wire \registerArray[2][14]~q ;
wire \registerArray[3][14]~q ;
wire \registerArray[1][14]~q ;
wire \Mux49~4_combout ;
wire \Mux49~5_combout ;
wire \Mux49~6_combout ;
wire \registerArray[27][14]~feeder_combout ;
wire \registerArray[27][14]~q ;
wire \registerArray[31][14]~q ;
wire \registerArray[19][14]~q ;
wire \Mux49~17_combout ;
wire \Mux49~18_combout ;
wire \registerArray[20][14]~q ;
wire \registerArray[28][14]~q ;
wire \registerArray[16][14]~feeder_combout ;
wire \registerArray[16][14]~q ;
wire \registerArray[24][14]~q ;
wire \Mux49~14_combout ;
wire \Mux49~15_combout ;
wire \registerArray[30][14]~q ;
wire \registerArray[18][14]~q ;
wire \registerArray[26][14]~q ;
wire \Mux49~12_combout ;
wire \Mux49~13_combout ;
wire \Mux49~16_combout ;
wire \registerArray[25][14]~q ;
wire \registerArray[29][14]~q ;
wire \registerArray[17][14]~q ;
wire \Mux49~10_combout ;
wire \Mux49~11_combout ;
wire \registerArray[14][13]~feeder_combout ;
wire \registerArray[14][13]~q ;
wire \registerArray[15][13]~feeder_combout ;
wire \registerArray[15][13]~q ;
wire \registerArray[12][13]~feeder_combout ;
wire \registerArray[12][13]~q ;
wire \registerArray[13][13]~q ;
wire \Mux50~7_combout ;
wire \Mux50~8_combout ;
wire \registerArray[6][13]~q ;
wire \registerArray[4][13]~q ;
wire \Mux50~0_combout ;
wire \registerArray[7][13]~q ;
wire \Mux50~1_combout ;
wire \registerArray[2][13]~q ;
wire \registerArray[3][13]~feeder_combout ;
wire \registerArray[3][13]~q ;
wire \registerArray[1][13]~q ;
wire \Mux50~4_combout ;
wire \Mux50~5_combout ;
wire \registerArray[8][13]~q ;
wire \Mux50~2_combout ;
wire \registerArray[11][13]~q ;
wire \Mux50~3_combout ;
wire \Mux50~6_combout ;
wire \registerArray[27][13]~q ;
wire \registerArray[19][13]~q ;
wire \Mux50~17_combout ;
wire \registerArray[23][13]~q ;
wire \registerArray[31][13]~q ;
wire \Mux50~18_combout ;
wire \registerArray[18][13]~q ;
wire \registerArray[22][13]~q ;
wire \Mux50~12_combout ;
wire \registerArray[30][13]~q ;
wire \registerArray[26][13]~q ;
wire \Mux50~13_combout ;
wire \registerArray[28][13]~q ;
wire \registerArray[16][13]~q ;
wire \Mux50~14_combout ;
wire \Mux50~15_combout ;
wire \Mux50~16_combout ;
wire \registerArray[21][13]~q ;
wire \registerArray[29][13]~feeder_combout ;
wire \registerArray[29][13]~q ;
wire \registerArray[25][13]~q ;
wire \registerArray[17][13]~feeder_combout ;
wire \registerArray[17][13]~q ;
wire \Mux50~10_combout ;
wire \Mux50~11_combout ;
wire \registerArray[14][12]~feeder_combout ;
wire \registerArray[14][12]~q ;
wire \registerArray[15][12]~q ;
wire \registerArray[12][12]~q ;
wire \Mux51~7_combout ;
wire \Mux51~8_combout ;
wire \registerArray[9][12]~feeder_combout ;
wire \registerArray[9][12]~q ;
wire \registerArray[11][12]~q ;
wire \registerArray[8][12]~feeder_combout ;
wire \registerArray[8][12]~q ;
wire \registerArray[10][12]~q ;
wire \Mux51~0_combout ;
wire \Mux51~1_combout ;
wire \registerArray[7][12]~feeder_combout ;
wire \registerArray[7][12]~q ;
wire \registerArray[6][12]~q ;
wire \registerArray[5][12]~q ;
wire \registerArray[4][12]~q ;
wire \Mux51~2_combout ;
wire \Mux51~3_combout ;
wire \registerArray[2][12]~feeder_combout ;
wire \registerArray[2][12]~q ;
wire \registerArray[3][12]~q ;
wire \Mux51~4_combout ;
wire \Mux51~5_combout ;
wire \Mux51~6_combout ;
wire \registerArray[29][12]~feeder_combout ;
wire \registerArray[29][12]~q ;
wire \registerArray[25][12]~q ;
wire \registerArray[17][12]~q ;
wire \Mux51~10_combout ;
wire \Mux51~11_combout ;
wire \registerArray[30][12]~q ;
wire \registerArray[26][12]~feeder_combout ;
wire \registerArray[26][12]~q ;
wire \registerArray[18][12]~q ;
wire \Mux51~12_combout ;
wire \Mux51~13_combout ;
wire \registerArray[20][12]~q ;
wire \registerArray[28][12]~q ;
wire \registerArray[16][12]~feeder_combout ;
wire \registerArray[16][12]~q ;
wire \Mux51~14_combout ;
wire \Mux51~15_combout ;
wire \Mux51~16_combout ;
wire \registerArray[27][12]~feeder_combout ;
wire \registerArray[27][12]~q ;
wire \registerArray[31][12]~q ;
wire \registerArray[19][12]~q ;
wire \registerArray[23][12]~feeder_combout ;
wire \registerArray[23][12]~q ;
wire \Mux51~17_combout ;
wire \Mux51~18_combout ;
wire \registerArray[12][11]~q ;
wire \Mux52~7_combout ;
wire \registerArray[15][11]~q ;
wire \registerArray[14][11]~q ;
wire \Mux52~8_combout ;
wire \registerArray[2][11]~q ;
wire \registerArray[3][11]~feeder_combout ;
wire \registerArray[3][11]~q ;
wire \registerArray[1][11]~q ;
wire \Mux52~4_combout ;
wire \Mux52~5_combout ;
wire \registerArray[11][11]~q ;
wire \registerArray[8][11]~q ;
wire \Mux52~2_combout ;
wire \Mux52~3_combout ;
wire \Mux52~6_combout ;
wire \registerArray[5][11]~q ;
wire \registerArray[4][11]~q ;
wire \Mux52~0_combout ;
wire \registerArray[7][11]~q ;
wire \registerArray[6][11]~q ;
wire \Mux52~1_combout ;
wire \registerArray[23][11]~feeder_combout ;
wire \registerArray[23][11]~q ;
wire \registerArray[31][11]~q ;
wire \registerArray[19][11]~q ;
wire \registerArray[27][11]~feeder_combout ;
wire \registerArray[27][11]~q ;
wire \Mux52~17_combout ;
wire \Mux52~18_combout ;
wire \registerArray[21][11]~q ;
wire \registerArray[29][11]~q ;
wire \registerArray[17][11]~feeder_combout ;
wire \registerArray[17][11]~q ;
wire \registerArray[25][11]~q ;
wire \Mux52~10_combout ;
wire \Mux52~11_combout ;
wire \registerArray[26][11]~q ;
wire \registerArray[30][11]~q ;
wire \registerArray[22][11]~q ;
wire \registerArray[18][11]~q ;
wire \Mux52~12_combout ;
wire \Mux52~13_combout ;
wire \registerArray[28][11]~q ;
wire \registerArray[20][11]~q ;
wire \registerArray[16][11]~q ;
wire \Mux52~14_combout ;
wire \Mux52~15_combout ;
wire \Mux52~16_combout ;
wire \registerArray[14][10]~feeder_combout ;
wire \registerArray[14][10]~q ;
wire \registerArray[15][10]~q ;
wire \registerArray[13][10]~feeder_combout ;
wire \registerArray[13][10]~q ;
wire \Mux53~7_combout ;
wire \Mux53~8_combout ;
wire \registerArray[9][10]~q ;
wire \registerArray[11][10]~q ;
wire \registerArray[8][10]~q ;
wire \Mux53~0_combout ;
wire \Mux53~1_combout ;
wire \registerArray[2][10]~feeder_combout ;
wire \registerArray[2][10]~q ;
wire \registerArray[1][10]~feeder_combout ;
wire \registerArray[1][10]~q ;
wire \Mux53~4_combout ;
wire \Mux53~5_combout ;
wire \registerArray[6][10]~feeder_combout ;
wire \registerArray[6][10]~q ;
wire \registerArray[7][10]~feeder_combout ;
wire \registerArray[7][10]~q ;
wire \registerArray[4][10]~q ;
wire \Mux53~2_combout ;
wire \Mux53~3_combout ;
wire \Mux53~6_combout ;
wire \registerArray[27][10]~feeder_combout ;
wire \registerArray[27][10]~q ;
wire \registerArray[31][10]~q ;
wire \registerArray[19][10]~q ;
wire \Mux53~17_combout ;
wire \Mux53~18_combout ;
wire \registerArray[25][10]~q ;
wire \registerArray[29][10]~q ;
wire \registerArray[17][10]~feeder_combout ;
wire \registerArray[17][10]~q ;
wire \Mux53~10_combout ;
wire \Mux53~11_combout ;
wire \registerArray[30][10]~q ;
wire \registerArray[26][10]~q ;
wire \registerArray[18][10]~q ;
wire \Mux53~12_combout ;
wire \Mux53~13_combout ;
wire \registerArray[20][10]~q ;
wire \registerArray[28][10]~q ;
wire \registerArray[16][10]~feeder_combout ;
wire \registerArray[16][10]~q ;
wire \Mux53~14_combout ;
wire \Mux53~15_combout ;
wire \Mux53~16_combout ;
wire \registerArray[14][9]~q ;
wire \registerArray[12][9]~q ;
wire \Mux54~7_combout ;
wire \registerArray[15][9]~q ;
wire \Mux54~8_combout ;
wire \registerArray[6][9]~q ;
wire \registerArray[7][9]~q ;
wire \registerArray[5][9]~q ;
wire \registerArray[4][9]~q ;
wire \Mux54~0_combout ;
wire \Mux54~1_combout ;
wire \registerArray[2][9]~feeder_combout ;
wire \registerArray[2][9]~q ;
wire \registerArray[1][9]~feeder_combout ;
wire \registerArray[1][9]~q ;
wire \Mux54~4_combout ;
wire \Mux54~5_combout ;
wire \registerArray[9][9]~q ;
wire \registerArray[11][9]~q ;
wire \registerArray[8][9]~q ;
wire \Mux54~2_combout ;
wire \Mux54~3_combout ;
wire \Mux54~6_combout ;
wire \registerArray[24][9]~q ;
wire \registerArray[28][9]~q ;
wire \Mux54~15_combout ;
wire \registerArray[22][9]~q ;
wire \registerArray[18][9]~q ;
wire \Mux54~12_combout ;
wire \registerArray[30][9]~q ;
wire \registerArray[26][9]~q ;
wire \Mux54~13_combout ;
wire \Mux54~16_combout ;
wire \registerArray[21][9]~q ;
wire \registerArray[29][9]~feeder_combout ;
wire \registerArray[29][9]~q ;
wire \registerArray[25][9]~feeder_combout ;
wire \registerArray[25][9]~q ;
wire \registerArray[17][9]~q ;
wire \Mux54~10_combout ;
wire \Mux54~11_combout ;
wire \registerArray[23][9]~q ;
wire \registerArray[31][9]~q ;
wire \registerArray[19][9]~q ;
wire \Mux54~17_combout ;
wire \Mux54~18_combout ;
wire \registerArray[9][8]~q ;
wire \registerArray[8][8]~q ;
wire \Mux55~0_combout ;
wire \registerArray[11][8]~q ;
wire \Mux55~1_combout ;
wire \registerArray[14][8]~feeder_combout ;
wire \registerArray[14][8]~q ;
wire \registerArray[15][8]~q ;
wire \registerArray[12][8]~q ;
wire \Mux55~7_combout ;
wire \Mux55~8_combout ;
wire \registerArray[6][8]~feeder_combout ;
wire \registerArray[6][8]~q ;
wire \registerArray[7][8]~q ;
wire \registerArray[4][8]~q ;
wire \Mux55~2_combout ;
wire \Mux55~3_combout ;
wire \registerArray[2][8]~q ;
wire \registerArray[1][8]~q ;
wire \Mux55~4_combout ;
wire \Mux55~5_combout ;
wire \Mux55~6_combout ;
wire \registerArray[19][8]~feeder_combout ;
wire \registerArray[19][8]~q ;
wire \registerArray[23][8]~feeder_combout ;
wire \registerArray[23][8]~q ;
wire \Mux55~17_combout ;
wire \registerArray[27][8]~q ;
wire \registerArray[31][8]~q ;
wire \Mux55~18_combout ;
wire \registerArray[30][8]~q ;
wire \registerArray[18][8]~q ;
wire \Mux55~12_combout ;
wire \Mux55~13_combout ;
wire \registerArray[20][8]~q ;
wire \registerArray[28][8]~q ;
wire \Mux55~15_combout ;
wire \Mux55~16_combout ;
wire \registerArray[29][8]~feeder_combout ;
wire \registerArray[29][8]~q ;
wire \registerArray[25][8]~feeder_combout ;
wire \registerArray[25][8]~q ;
wire \registerArray[17][8]~feeder_combout ;
wire \registerArray[17][8]~q ;
wire \Mux55~10_combout ;
wire \Mux55~11_combout ;
wire \registerArray[14][7]~feeder_combout ;
wire \registerArray[14][7]~q ;
wire \registerArray[15][7]~q ;
wire \registerArray[13][7]~q ;
wire \registerArray[12][7]~q ;
wire \Mux56~7_combout ;
wire \Mux56~8_combout ;
wire \registerArray[6][7]~q ;
wire \registerArray[7][7]~q ;
wire \registerArray[4][7]~feeder_combout ;
wire \registerArray[4][7]~q ;
wire \Mux56~0_combout ;
wire \Mux56~1_combout ;
wire \registerArray[2][7]~q ;
wire \Mux56~5_combout ;
wire \registerArray[11][7]~q ;
wire \registerArray[8][7]~q ;
wire \Mux56~2_combout ;
wire \Mux56~3_combout ;
wire \Mux56~6_combout ;
wire \registerArray[23][7]~q ;
wire \registerArray[31][7]~q ;
wire \registerArray[19][7]~q ;
wire \Mux56~17_combout ;
wire \Mux56~18_combout ;
wire \registerArray[21][7]~q ;
wire \registerArray[29][7]~q ;
wire \registerArray[25][7]~q ;
wire \registerArray[17][7]~q ;
wire \Mux56~10_combout ;
wire \Mux56~11_combout ;
wire \registerArray[28][7]~q ;
wire \registerArray[16][7]~q ;
wire \Mux56~14_combout ;
wire \Mux56~15_combout ;
wire \registerArray[30][7]~q ;
wire \registerArray[18][7]~q ;
wire \Mux56~12_combout ;
wire \Mux56~13_combout ;
wire \Mux56~16_combout ;
wire \registerArray[9][6]~q ;
wire \registerArray[11][6]~q ;
wire \registerArray[8][6]~q ;
wire \Mux57~0_combout ;
wire \Mux57~1_combout ;
wire \registerArray[2][6]~q ;
wire \registerArray[3][6]~feeder_combout ;
wire \registerArray[3][6]~q ;
wire \registerArray[1][6]~q ;
wire \Mux57~4_combout ;
wire \Mux57~5_combout ;
wire \registerArray[7][6]~q ;
wire \registerArray[5][6]~feeder_combout ;
wire \registerArray[5][6]~q ;
wire \Mux57~2_combout ;
wire \Mux57~3_combout ;
wire \Mux57~6_combout ;
wire \registerArray[14][6]~q ;
wire \registerArray[15][6]~q ;
wire \registerArray[12][6]~q ;
wire \registerArray[13][6]~q ;
wire \Mux57~7_combout ;
wire \Mux57~8_combout ;
wire \registerArray[25][6]~q ;
wire \registerArray[29][6]~q ;
wire \registerArray[21][6]~q ;
wire \registerArray[17][6]~q ;
wire \Mux57~10_combout ;
wire \Mux57~11_combout ;
wire \registerArray[27][6]~feeder_combout ;
wire \registerArray[27][6]~q ;
wire \registerArray[31][6]~q ;
wire \registerArray[23][6]~q ;
wire \Mux57~17_combout ;
wire \Mux57~18_combout ;
wire \registerArray[22][6]~q ;
wire \registerArray[30][6]~q ;
wire \registerArray[18][6]~q ;
wire \Mux57~12_combout ;
wire \Mux57~13_combout ;
wire \registerArray[28][6]~q ;
wire \registerArray[24][6]~q ;
wire \Mux57~14_combout ;
wire \Mux57~15_combout ;
wire \Mux57~16_combout ;
wire \registerArray[31][2]~q ;
wire \registerArray[19][2]~q ;
wire \registerArray[27][2]~q ;
wire \Mux29~7_combout ;
wire \Mux29~8_combout ;
wire \registerArray[30][2]~q ;
wire \registerArray[26][2]~q ;
wire \registerArray[22][2]~q ;
wire \Mux29~2_combout ;
wire \Mux29~3_combout ;
wire \registerArray[28][2]~q ;
wire \registerArray[24][2]~q ;
wire \registerArray[16][2]~q ;
wire \registerArray[20][2]~q ;
wire \Mux29~4_combout ;
wire \Mux29~5_combout ;
wire \Mux29~6_combout ;
wire \registerArray[21][2]~feeder_combout ;
wire \registerArray[21][2]~q ;
wire \registerArray[17][2]~q ;
wire \Mux29~0_combout ;
wire \Mux29~1_combout ;
wire \Mux29~9_combout ;
wire \registerArray[7][2]~feeder_combout ;
wire \registerArray[7][2]~q ;
wire \registerArray[6][2]~q ;
wire \registerArray[5][2]~q ;
wire \Mux29~10_combout ;
wire \Mux29~11_combout ;
wire \registerArray[12][2]~feeder_combout ;
wire \registerArray[12][2]~q ;
wire \registerArray[13][2]~q ;
wire \Mux29~17_combout ;
wire \registerArray[14][2]~q ;
wire \Mux29~18_combout ;
wire \registerArray[2][2]~q ;
wire \registerArray[1][2]~feeder_combout ;
wire \registerArray[1][2]~q ;
wire \Mux29~14_combout ;
wire \Mux29~15_combout ;
wire \registerArray[9][2]~q ;
wire \registerArray[11][2]~q ;
wire \registerArray[8][2]~q ;
wire \Mux29~12_combout ;
wire \Mux29~13_combout ;
wire \Mux29~16_combout ;
wire \Mux29~19_combout ;
wire \registerArray[25][1]~q ;
wire \registerArray[21][1]~feeder_combout ;
wire \registerArray[21][1]~q ;
wire \Mux30~0_combout ;
wire \Mux30~1_combout ;
wire \registerArray[30][1]~q ;
wire \registerArray[22][1]~q ;
wire \registerArray[18][1]~feeder_combout ;
wire \registerArray[18][1]~q ;
wire \registerArray[26][1]~q ;
wire \Mux30~2_combout ;
wire \Mux30~3_combout ;
wire \registerArray[28][1]~q ;
wire \registerArray[20][1]~q ;
wire \registerArray[16][1]~q ;
wire \registerArray[24][1]~q ;
wire \Mux30~4_combout ;
wire \Mux30~5_combout ;
wire \Mux30~6_combout ;
wire \registerArray[31][1]~q ;
wire \registerArray[27][1]~feeder_combout ;
wire \registerArray[27][1]~q ;
wire \Mux30~8_combout ;
wire \Mux30~9_combout ;
wire \registerArray[9][1]~q ;
wire \registerArray[11][1]~q ;
wire \Mux30~11_combout ;
wire \registerArray[14][1]~feeder_combout ;
wire \registerArray[14][1]~q ;
wire \registerArray[15][1]~q ;
wire \registerArray[13][1]~feeder_combout ;
wire \registerArray[13][1]~q ;
wire \registerArray[12][1]~feeder_combout ;
wire \registerArray[12][1]~q ;
wire \Mux30~17_combout ;
wire \Mux30~18_combout ;
wire \registerArray[1][1]~q ;
wire \registerArray[3][1]~feeder_combout ;
wire \registerArray[3][1]~q ;
wire \Mux30~14_combout ;
wire \Mux30~15_combout ;
wire \registerArray[6][1]~feeder_combout ;
wire \registerArray[6][1]~q ;
wire \registerArray[7][1]~q ;
wire \registerArray[5][1]~q ;
wire \Mux30~12_combout ;
wire \Mux30~13_combout ;
wire \Mux30~16_combout ;
wire \Mux30~19_combout ;
wire \Mux62~7_combout ;
wire \Mux62~8_combout ;
wire \registerArray[4][1]~q ;
wire \Mux62~0_combout ;
wire \Mux62~1_combout ;
wire \registerArray[8][1]~q ;
wire \Mux62~2_combout ;
wire \Mux62~3_combout ;
wire \registerArray[2][1]~q ;
wire \Mux62~4_combout ;
wire \Mux62~5_combout ;
wire \Mux62~6_combout ;
wire \registerArray[23][1]~q ;
wire \registerArray[19][1]~q ;
wire \Mux62~17_combout ;
wire \Mux62~18_combout ;
wire \Mux62~14_combout ;
wire \Mux62~15_combout ;
wire \Mux62~12_combout ;
wire \Mux62~13_combout ;
wire \Mux62~16_combout ;
wire \registerArray[29][1]~feeder_combout ;
wire \registerArray[29][1]~q ;
wire \registerArray[17][1]~q ;
wire \Mux62~10_combout ;
wire \Mux62~11_combout ;
wire \registerArray[7][4]~q ;
wire \registerArray[6][4]~q ;
wire \registerArray[5][4]~q ;
wire \Mux27~10_combout ;
wire \Mux27~11_combout ;
wire \registerArray[9][4]~q ;
wire \registerArray[11][4]~q ;
wire \registerArray[8][4]~q ;
wire \Mux27~12_combout ;
wire \Mux27~13_combout ;
wire \registerArray[2][4]~q ;
wire \registerArray[3][4]~feeder_combout ;
wire \registerArray[3][4]~q ;
wire \Mux27~14_combout ;
wire \Mux27~15_combout ;
wire \Mux27~16_combout ;
wire \registerArray[15][4]~feeder_combout ;
wire \registerArray[15][4]~q ;
wire \registerArray[13][4]~q ;
wire \Mux27~17_combout ;
wire \Mux27~18_combout ;
wire \Mux27~19_combout ;
wire \registerArray[21][4]~feeder_combout ;
wire \registerArray[21][4]~q ;
wire \registerArray[17][4]~q ;
wire \Mux27~0_combout ;
wire \Mux27~1_combout ;
wire \registerArray[30][4]~q ;
wire \registerArray[26][4]~q ;
wire \registerArray[18][4]~q ;
wire \registerArray[22][4]~q ;
wire \Mux27~2_combout ;
wire \Mux27~3_combout ;
wire \registerArray[28][4]~q ;
wire \registerArray[24][4]~q ;
wire \registerArray[16][4]~q ;
wire \registerArray[20][4]~q ;
wire \Mux27~4_combout ;
wire \Mux27~5_combout ;
wire \Mux27~6_combout ;
wire \registerArray[23][4]~feeder_combout ;
wire \registerArray[23][4]~q ;
wire \registerArray[19][4]~q ;
wire \registerArray[27][4]~q ;
wire \Mux27~7_combout ;
wire \Mux27~8_combout ;
wire \Mux27~9_combout ;
wire \registerArray[29][3]~q ;
wire \registerArray[21][3]~q ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \registerArray[30][3]~q ;
wire \registerArray[22][3]~q ;
wire \Mux28~3_combout ;
wire \registerArray[16][3]~q ;
wire \registerArray[24][3]~q ;
wire \Mux28~4_combout ;
wire \registerArray[20][3]~q ;
wire \Mux28~5_combout ;
wire \Mux28~6_combout ;
wire \registerArray[27][3]~feeder_combout ;
wire \registerArray[27][3]~q ;
wire \registerArray[23][3]~q ;
wire \Mux28~7_combout ;
wire \Mux28~8_combout ;
wire \Mux28~9_combout ;
wire \registerArray[10][3]~q ;
wire \registerArray[8][3]~feeder_combout ;
wire \registerArray[8][3]~q ;
wire \Mux28~10_combout ;
wire \registerArray[9][3]~q ;
wire \Mux28~11_combout ;
wire \registerArray[15][3]~feeder_combout ;
wire \registerArray[15][3]~q ;
wire \registerArray[13][3]~q ;
wire \Mux28~17_combout ;
wire \Mux28~18_combout ;
wire \registerArray[6][3]~q ;
wire \registerArray[7][3]~q ;
wire \registerArray[4][3]~q ;
wire \Mux28~12_combout ;
wire \Mux28~13_combout ;
wire \registerArray[1][3]~q ;
wire \registerArray[3][3]~q ;
wire \Mux28~14_combout ;
wire \Mux28~15_combout ;
wire \Mux28~16_combout ;
wire \Mux28~19_combout ;
wire \Mux61~4_combout ;
wire \Mux61~5_combout ;
wire \registerArray[18][2]~q ;
wire \Mux61~2_combout ;
wire \Mux61~3_combout ;
wire \Mux61~6_combout ;
wire \registerArray[23][2]~feeder_combout ;
wire \registerArray[23][2]~q ;
wire \Mux61~7_combout ;
wire \Mux61~8_combout ;
wire \registerArray[29][2]~feeder_combout ;
wire \registerArray[29][2]~q ;
wire \registerArray[25][2]~feeder_combout ;
wire \registerArray[25][2]~q ;
wire \Mux61~0_combout ;
wire \Mux61~1_combout ;
wire \registerArray[10][2]~feeder_combout ;
wire \registerArray[10][2]~q ;
wire \Mux61~10_combout ;
wire \Mux61~11_combout ;
wire \registerArray[15][2]~q ;
wire \Mux61~17_combout ;
wire \Mux61~18_combout ;
wire \registerArray[4][2]~q ;
wire \Mux61~12_combout ;
wire \Mux61~13_combout ;
wire \registerArray[3][2]~feeder_combout ;
wire \registerArray[3][2]~q ;
wire \Mux61~14_combout ;
wire \Mux61~15_combout ;
wire \Mux61~16_combout ;
wire \registerArray[21][8]~feeder_combout ;
wire \registerArray[21][8]~q ;
wire \Mux23~0_combout ;
wire \Mux23~1_combout ;
wire \registerArray[16][8]~q ;
wire \Mux23~4_combout ;
wire \Mux23~5_combout ;
wire \Mux23~6_combout ;
wire \Mux23~7_combout ;
wire \Mux23~8_combout ;
wire \Mux23~9_combout ;
wire \registerArray[3][8]~q ;
wire \Mux23~14_combout ;
wire \Mux23~15_combout ;
wire \registerArray[10][8]~q ;
wire \Mux23~12_combout ;
wire \Mux23~13_combout ;
wire \Mux23~16_combout ;
wire \registerArray[13][8]~q ;
wire \Mux23~17_combout ;
wire \Mux23~18_combout ;
wire \Mux23~10_combout ;
wire \Mux23~11_combout ;
wire \Mux23~19_combout ;
wire \Mux24~0_combout ;
wire \Mux24~1_combout ;
wire \registerArray[27][7]~q ;
wire \Mux24~7_combout ;
wire \Mux24~8_combout ;
wire \registerArray[26][7]~feeder_combout ;
wire \registerArray[26][7]~q ;
wire \Mux24~2_combout ;
wire \Mux24~3_combout ;
wire \registerArray[20][7]~q ;
wire \registerArray[24][7]~q ;
wire \Mux24~4_combout ;
wire \Mux24~5_combout ;
wire \Mux24~6_combout ;
wire \Mux24~9_combout ;
wire \Mux24~17_combout ;
wire \Mux24~18_combout ;
wire \registerArray[9][7]~q ;
wire \Mux24~11_combout ;
wire \registerArray[5][7]~q ;
wire \Mux24~12_combout ;
wire \Mux24~13_combout ;
wire \Mux24~16_combout ;
wire \Mux24~19_combout ;
wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \registerArray[19][6]~q ;
wire \Mux25~7_combout ;
wire \Mux25~8_combout ;
wire \registerArray[16][6]~feeder_combout ;
wire \registerArray[16][6]~q ;
wire \registerArray[20][6]~q ;
wire \Mux25~4_combout ;
wire \Mux25~5_combout ;
wire \registerArray[26][6]~q ;
wire \Mux25~2_combout ;
wire \Mux25~3_combout ;
wire \Mux25~6_combout ;
wire \Mux25~9_combout ;
wire \Mux25~10_combout ;
wire \Mux25~11_combout ;
wire \Mux25~17_combout ;
wire \Mux25~18_combout ;
wire \registerArray[10][6]~q ;
wire \Mux25~12_combout ;
wire \Mux25~13_combout ;
wire \Mux25~14_combout ;
wire \Mux25~15_combout ;
wire \Mux25~16_combout ;
wire \Mux25~19_combout ;
wire \Mux26~7_combout ;
wire \Mux26~8_combout ;
wire \registerArray[24][5]~q ;
wire \Mux26~4_combout ;
wire \Mux26~5_combout ;
wire \registerArray[22][5]~q ;
wire \registerArray[26][5]~q ;
wire \Mux26~2_combout ;
wire \Mux26~3_combout ;
wire \Mux26~6_combout ;
wire \registerArray[25][5]~q ;
wire \Mux26~0_combout ;
wire \Mux26~1_combout ;
wire \Mux26~9_combout ;
wire \registerArray[10][5]~q ;
wire \Mux26~10_combout ;
wire \Mux26~11_combout ;
wire \registerArray[13][5]~feeder_combout ;
wire \registerArray[13][5]~q ;
wire \Mux26~17_combout ;
wire \Mux26~18_combout ;
wire \registerArray[1][5]~q ;
wire \Mux26~14_combout ;
wire \registerArray[2][5]~feeder_combout ;
wire \registerArray[2][5]~q ;
wire \Mux26~15_combout ;
wire \Mux26~16_combout ;
wire \Mux26~19_combout ;
wire \registerArray[28][3]~q ;
wire \Mux60~4_combout ;
wire \Mux60~5_combout ;
wire \registerArray[18][3]~q ;
wire \Mux60~2_combout ;
wire \Mux60~3_combout ;
wire \Mux60~6_combout ;
wire \registerArray[25][3]~feeder_combout ;
wire \registerArray[25][3]~q ;
wire \Mux60~0_combout ;
wire \Mux60~1_combout ;
wire \registerArray[19][3]~q ;
wire \Mux60~7_combout ;
wire \registerArray[31][3]~q ;
wire \Mux60~8_combout ;
wire \registerArray[14][3]~q ;
wire \registerArray[12][3]~feeder_combout ;
wire \registerArray[12][3]~q ;
wire \Mux60~17_combout ;
wire \Mux60~18_combout ;
wire \registerArray[5][3]~q ;
wire \Mux60~10_combout ;
wire \Mux60~11_combout ;
wire \registerArray[2][3]~feeder_combout ;
wire \registerArray[2][3]~q ;
wire \Mux60~14_combout ;
wire \Mux60~15_combout ;
wire \registerArray[11][3]~feeder_combout ;
wire \registerArray[11][3]~q ;
wire \Mux60~12_combout ;
wire \Mux60~13_combout ;
wire \Mux60~16_combout ;
wire \registerArray[7][16]~feeder_combout ;
wire \registerArray[7][16]~q ;
wire \Mux15~10_combout ;
wire \Mux15~11_combout ;
wire \Mux15~14_combout ;
wire \Mux15~15_combout ;
wire \registerArray[10][16]~q ;
wire \Mux15~12_combout ;
wire \Mux15~13_combout ;
wire \Mux15~16_combout ;
wire \registerArray[13][16]~feeder_combout ;
wire \registerArray[13][16]~q ;
wire \Mux15~17_combout ;
wire \Mux15~18_combout ;
wire \Mux15~19_combout ;
wire \registerArray[22][16]~q ;
wire \Mux15~2_combout ;
wire \Mux15~3_combout ;
wire \Mux15~6_combout ;
wire \Mux15~7_combout ;
wire \Mux15~8_combout ;
wire \Mux15~0_combout ;
wire \Mux15~1_combout ;
wire \Mux15~9_combout ;
wire \Mux16~2_combout ;
wire \Mux16~3_combout ;
wire \registerArray[20][15]~q ;
wire \registerArray[24][15]~q ;
wire \Mux16~4_combout ;
wire \Mux16~5_combout ;
wire \Mux16~6_combout ;
wire \Mux16~7_combout ;
wire \Mux16~8_combout ;
wire \registerArray[25][15]~q ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \Mux16~9_combout ;
wire \registerArray[5][15]~feeder_combout ;
wire \registerArray[5][15]~q ;
wire \Mux16~12_combout ;
wire \Mux16~13_combout ;
wire \Mux16~16_combout ;
wire \registerArray[13][15]~feeder_combout ;
wire \registerArray[13][15]~q ;
wire \Mux16~17_combout ;
wire \Mux16~18_combout ;
wire \Mux16~10_combout ;
wire \Mux16~11_combout ;
wire \Mux16~19_combout ;
wire \Mux17~14_combout ;
wire \Mux17~15_combout ;
wire \Mux17~13_combout ;
wire \Mux17~16_combout ;
wire \registerArray[13][14]~q ;
wire \Mux17~17_combout ;
wire \Mux17~18_combout ;
wire \registerArray[6][14]~feeder_combout ;
wire \registerArray[6][14]~q ;
wire \Mux17~10_combout ;
wire \Mux17~11_combout ;
wire \Mux17~19_combout ;
wire \registerArray[21][14]~q ;
wire \Mux17~0_combout ;
wire \Mux17~1_combout ;
wire \registerArray[23][14]~feeder_combout ;
wire \registerArray[23][14]~q ;
wire \Mux17~7_combout ;
wire \Mux17~8_combout ;
wire \Mux17~4_combout ;
wire \Mux17~5_combout ;
wire \registerArray[22][14]~q ;
wire \Mux17~2_combout ;
wire \Mux17~3_combout ;
wire \Mux17~6_combout ;
wire \Mux17~9_combout ;
wire \Mux18~0_combout ;
wire \Mux18~1_combout ;
wire \Mux18~7_combout ;
wire \Mux18~8_combout ;
wire \Mux18~2_combout ;
wire \Mux18~3_combout ;
wire \Mux18~4_combout ;
wire \Mux18~5_combout ;
wire \Mux18~6_combout ;
wire \Mux18~9_combout ;
wire \registerArray[9][13]~q ;
wire \registerArray[10][13]~q ;
wire \Mux18~10_combout ;
wire \Mux18~11_combout ;
wire \Mux18~17_combout ;
wire \Mux18~18_combout ;
wire \Mux18~14_combout ;
wire \Mux18~15_combout ;
wire \Mux18~12_combout ;
wire \Mux18~13_combout ;
wire \Mux18~16_combout ;
wire \Mux18~19_combout ;
wire \Mux19~7_combout ;
wire \Mux19~8_combout ;
wire \Mux19~0_combout ;
wire \Mux19~1_combout ;
wire \registerArray[24][12]~q ;
wire \Mux19~4_combout ;
wire \Mux19~5_combout ;
wire \Mux19~2_combout ;
wire \Mux19~3_combout ;
wire \Mux19~6_combout ;
wire \Mux19~9_combout ;
wire \Mux19~10_combout ;
wire \Mux19~11_combout ;
wire \registerArray[13][12]~feeder_combout ;
wire \registerArray[13][12]~q ;
wire \Mux19~17_combout ;
wire \Mux19~18_combout ;
wire \Mux19~15_combout ;
wire \Mux19~12_combout ;
wire \Mux19~13_combout ;
wire \Mux19~16_combout ;
wire \Mux19~19_combout ;
wire \Mux20~2_combout ;
wire \Mux20~3_combout ;
wire \registerArray[24][11]~q ;
wire \Mux20~4_combout ;
wire \Mux20~5_combout ;
wire \Mux20~6_combout ;
wire \Mux20~0_combout ;
wire \Mux20~1_combout ;
wire \Mux20~7_combout ;
wire \Mux20~8_combout ;
wire \Mux20~9_combout ;
wire \registerArray[9][11]~feeder_combout ;
wire \registerArray[9][11]~q ;
wire \registerArray[10][11]~q ;
wire \Mux20~10_combout ;
wire \Mux20~11_combout ;
wire \registerArray[13][11]~q ;
wire \Mux20~17_combout ;
wire \Mux20~18_combout ;
wire \Mux20~12_combout ;
wire \Mux20~13_combout ;
wire \Mux20~14_combout ;
wire \Mux20~15_combout ;
wire \Mux20~16_combout ;
wire \Mux20~19_combout ;
wire \Mux21~7_combout ;
wire \Mux21~8_combout ;
wire \Mux21~0_combout ;
wire \Mux21~1_combout ;
wire \registerArray[24][10]~q ;
wire \Mux21~4_combout ;
wire \Mux21~5_combout ;
wire \registerArray[22][10]~q ;
wire \Mux21~2_combout ;
wire \Mux21~3_combout ;
wire \Mux21~6_combout ;
wire \Mux21~9_combout ;
wire \registerArray[12][10]~q ;
wire \Mux21~17_combout ;
wire \Mux21~18_combout ;
wire \registerArray[5][10]~q ;
wire \Mux21~10_combout ;
wire \Mux21~11_combout ;
wire \Mux21~13_combout ;
wire \Mux21~16_combout ;
wire \Mux21~19_combout ;
wire \Mux22~0_combout ;
wire \Mux22~1_combout ;
wire \Mux22~2_combout ;
wire \Mux22~3_combout ;
wire \Mux22~4_combout ;
wire \registerArray[20][9]~q ;
wire \Mux22~5_combout ;
wire \Mux22~6_combout ;
wire \registerArray[27][9]~q ;
wire \Mux22~7_combout ;
wire \Mux22~8_combout ;
wire \Mux22~9_combout ;
wire \registerArray[13][9]~q ;
wire \Mux22~17_combout ;
wire \Mux22~18_combout ;
wire \registerArray[10][9]~q ;
wire \Mux22~10_combout ;
wire \Mux22~11_combout ;
wire \Mux22~12_combout ;
wire \Mux22~13_combout ;
wire \registerArray[3][9]~q ;
wire \Mux22~14_combout ;
wire \Mux22~15_combout ;
wire \Mux22~16_combout ;
wire \Mux22~19_combout ;
wire \Mux59~4_combout ;
wire \Mux59~5_combout ;
wire \Mux59~2_combout ;
wire \Mux59~3_combout ;
wire \Mux59~6_combout ;
wire \Mux59~0_combout ;
wire \registerArray[25][4]~feeder_combout ;
wire \registerArray[25][4]~q ;
wire \registerArray[29][4]~q ;
wire \Mux59~1_combout ;
wire \registerArray[31][4]~q ;
wire \Mux59~7_combout ;
wire \Mux59~8_combout ;
wire \registerArray[10][4]~feeder_combout ;
wire \registerArray[10][4]~q ;
wire \Mux59~10_combout ;
wire \Mux59~11_combout ;
wire \registerArray[14][4]~feeder_combout ;
wire \registerArray[14][4]~q ;
wire \registerArray[12][4]~feeder_combout ;
wire \registerArray[12][4]~q ;
wire \Mux59~17_combout ;
wire \Mux59~18_combout ;
wire \registerArray[1][4]~feeder_combout ;
wire \registerArray[1][4]~q ;
wire \Mux59~14_combout ;
wire \Mux59~15_combout ;
wire \registerArray[4][4]~q ;
wire \Mux59~12_combout ;
wire \Mux59~13_combout ;
wire \Mux59~16_combout ;
wire \registerArray[10][31]~q ;
wire \Mux0~10_combout ;
wire \Mux0~11_combout ;
wire \registerArray[4][31]~q ;
wire \Mux0~12_combout ;
wire \Mux0~13_combout ;
wire \Mux0~14_combout ;
wire \Mux0~15_combout ;
wire \Mux0~16_combout ;
wire \Mux0~17_combout ;
wire \Mux0~18_combout ;
wire \Mux0~19_combout ;
wire \Mux0~7_combout ;
wire \Mux0~8_combout ;
wire \registerArray[24][31]~q ;
wire \Mux0~4_combout ;
wire \Mux0~5_combout ;
wire \registerArray[22][31]~q ;
wire \registerArray[26][31]~q ;
wire \Mux0~2_combout ;
wire \Mux0~3_combout ;
wire \Mux0~6_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \Mux0~9_combout ;
wire \registerArray[26][29]~feeder_combout ;
wire \registerArray[26][29]~q ;
wire \Mux2~2_combout ;
wire \Mux2~3_combout ;
wire \Mux2~6_combout ;
wire \Mux2~7_combout ;
wire \Mux2~8_combout ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \Mux2~9_combout ;
wire \Mux2~17_combout ;
wire \Mux2~18_combout ;
wire \Mux2~14_combout ;
wire \Mux2~15_combout ;
wire \registerArray[5][29]~q ;
wire \Mux2~12_combout ;
wire \Mux2~13_combout ;
wire \Mux2~16_combout ;
wire \Mux2~10_combout ;
wire \Mux2~11_combout ;
wire \Mux2~19_combout ;
wire \registerArray[13][30]~q ;
wire \Mux1~17_combout ;
wire \Mux1~18_combout ;
wire \registerArray[5][30]~feeder_combout ;
wire \registerArray[5][30]~q ;
wire \Mux1~10_combout ;
wire \Mux1~11_combout ;
wire \registerArray[3][30]~q ;
wire \Mux1~14_combout ;
wire \Mux1~15_combout ;
wire \Mux1~13_combout ;
wire \Mux1~16_combout ;
wire \Mux1~19_combout ;
wire \registerArray[24][30]~feeder_combout ;
wire \registerArray[24][30]~q ;
wire \registerArray[28][30]~feeder_combout ;
wire \registerArray[28][30]~q ;
wire \Mux1~4_combout ;
wire \Mux1~5_combout ;
wire \Mux1~6_combout ;
wire \Mux1~7_combout ;
wire \registerArray[23][30]~q ;
wire \Mux1~8_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Mux1~9_combout ;
wire \Mux3~7_combout ;
wire \Mux3~8_combout ;
wire \registerArray[17][28]~feeder_combout ;
wire \registerArray[17][28]~q ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \registerArray[24][28]~q ;
wire \registerArray[16][28]~feeder_combout ;
wire \registerArray[16][28]~q ;
wire \Mux3~4_combout ;
wire \Mux3~5_combout ;
wire \registerArray[22][28]~q ;
wire \Mux3~2_combout ;
wire \Mux3~3_combout ;
wire \Mux3~6_combout ;
wire \Mux3~9_combout ;
wire \Mux3~17_combout ;
wire \Mux3~18_combout ;
wire \registerArray[6][28]~q ;
wire \Mux3~10_combout ;
wire \Mux3~11_combout ;
wire \Mux3~14_combout ;
wire \Mux3~15_combout ;
wire \Mux3~12_combout ;
wire \Mux3~13_combout ;
wire \Mux3~16_combout ;
wire \Mux3~19_combout ;
wire \Mux4~0_combout ;
wire \Mux4~1_combout ;
wire \Mux4~7_combout ;
wire \Mux4~8_combout ;
wire \registerArray[22][27]~q ;
wire \registerArray[26][27]~q ;
wire \Mux4~2_combout ;
wire \Mux4~3_combout ;
wire \registerArray[20][27]~q ;
wire \Mux4~4_combout ;
wire \Mux4~5_combout ;
wire \Mux4~6_combout ;
wire \Mux4~9_combout ;
wire \Mux4~17_combout ;
wire \Mux4~18_combout ;
wire \Mux4~12_combout ;
wire \Mux4~13_combout ;
wire \Mux4~14_combout ;
wire \Mux4~15_combout ;
wire \Mux4~16_combout ;
wire \registerArray[10][27]~q ;
wire \Mux4~10_combout ;
wire \Mux4~11_combout ;
wire \Mux4~19_combout ;
wire \Mux5~10_combout ;
wire \Mux5~11_combout ;
wire \Mux5~14_combout ;
wire \Mux5~15_combout ;
wire \Mux5~12_combout ;
wire \Mux5~13_combout ;
wire \Mux5~16_combout ;
wire \Mux5~17_combout ;
wire \Mux5~18_combout ;
wire \Mux5~19_combout ;
wire \Mux5~0_combout ;
wire \Mux5~1_combout ;
wire \Mux5~7_combout ;
wire \Mux5~8_combout ;
wire \Mux5~2_combout ;
wire \Mux5~3_combout ;
wire \registerArray[20][26]~feeder_combout ;
wire \registerArray[20][26]~q ;
wire \Mux5~4_combout ;
wire \Mux5~5_combout ;
wire \Mux5~6_combout ;
wire \Mux5~9_combout ;
wire \registerArray[27][25]~q ;
wire \Mux6~7_combout ;
wire \Mux6~8_combout ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \registerArray[24][25]~q ;
wire \Mux6~4_combout ;
wire \Mux6~5_combout ;
wire \Mux6~6_combout ;
wire \Mux6~9_combout ;
wire \registerArray[9][25]~q ;
wire \registerArray[10][25]~q ;
wire \Mux6~10_combout ;
wire \Mux6~11_combout ;
wire \Mux6~17_combout ;
wire \Mux6~18_combout ;
wire \Mux6~14_combout ;
wire \Mux6~15_combout ;
wire \Mux6~12_combout ;
wire \Mux6~13_combout ;
wire \Mux6~16_combout ;
wire \Mux6~19_combout ;
wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \registerArray[16][24]~feeder_combout ;
wire \registerArray[16][24]~q ;
wire \Mux7~4_combout ;
wire \Mux7~5_combout ;
wire \Mux7~2_combout ;
wire \registerArray[26][24]~q ;
wire \Mux7~3_combout ;
wire \Mux7~6_combout ;
wire \registerArray[23][24]~q ;
wire \Mux7~7_combout ;
wire \Mux7~8_combout ;
wire \Mux7~9_combout ;
wire \Mux7~17_combout ;
wire \Mux7~18_combout ;
wire \registerArray[3][24]~q ;
wire \Mux7~14_combout ;
wire \Mux7~15_combout ;
wire \registerArray[10][24]~q ;
wire \Mux7~12_combout ;
wire \Mux7~13_combout ;
wire \Mux7~16_combout ;
wire \registerArray[7][24]~q ;
wire \Mux7~11_combout ;
wire \Mux7~19_combout ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \registerArray[24][23]~feeder_combout ;
wire \registerArray[24][23]~q ;
wire \Mux8~4_combout ;
wire \Mux8~5_combout ;
wire \Mux8~6_combout ;
wire \registerArray[27][23]~q ;
wire \Mux8~7_combout ;
wire \Mux8~8_combout ;
wire \Mux8~9_combout ;
wire \registerArray[3][23]~q ;
wire \Mux8~14_combout ;
wire \Mux8~15_combout ;
wire \registerArray[5][23]~q ;
wire \Mux8~12_combout ;
wire \Mux8~13_combout ;
wire \Mux8~16_combout ;
wire \Mux8~17_combout ;
wire \Mux8~18_combout ;
wire \registerArray[10][23]~q ;
wire \Mux8~10_combout ;
wire \Mux8~11_combout ;
wire \Mux8~19_combout ;
wire \registerArray[3][22]~q ;
wire \Mux9~14_combout ;
wire \Mux9~15_combout ;
wire \registerArray[10][22]~feeder_combout ;
wire \registerArray[10][22]~q ;
wire \Mux9~12_combout ;
wire \Mux9~13_combout ;
wire \Mux9~16_combout ;
wire \Mux9~17_combout ;
wire \Mux9~18_combout ;
wire \registerArray[6][22]~q ;
wire \Mux9~10_combout ;
wire \Mux9~11_combout ;
wire \Mux9~19_combout ;
wire \registerArray[23][22]~q ;
wire \Mux9~7_combout ;
wire \Mux9~8_combout ;
wire \Mux9~0_combout ;
wire \Mux9~1_combout ;
wire \Mux9~2_combout ;
wire \Mux9~3_combout ;
wire \registerArray[20][22]~q ;
wire \Mux9~4_combout ;
wire \Mux9~5_combout ;
wire \Mux9~6_combout ;
wire \Mux9~9_combout ;
wire \Mux10~17_combout ;
wire \Mux10~18_combout ;
wire \registerArray[3][21]~q ;
wire \Mux10~14_combout ;
wire \Mux10~15_combout ;
wire \registerArray[5][21]~q ;
wire \Mux10~12_combout ;
wire \Mux10~13_combout ;
wire \Mux10~16_combout ;
wire \registerArray[11][21]~feeder_combout ;
wire \registerArray[11][21]~q ;
wire \Mux10~11_combout ;
wire \Mux10~19_combout ;
wire \Mux10~0_combout ;
wire \Mux10~1_combout ;
wire \Mux10~7_combout ;
wire \Mux10~8_combout ;
wire \registerArray[24][21]~q ;
wire \registerArray[16][21]~feeder_combout ;
wire \registerArray[16][21]~q ;
wire \Mux10~4_combout ;
wire \Mux10~5_combout ;
wire \Mux10~6_combout ;
wire \Mux10~9_combout ;
wire \Mux11~17_combout ;
wire \Mux11~18_combout ;
wire \Mux11~12_combout ;
wire \Mux11~13_combout ;
wire \Mux11~16_combout ;
wire \registerArray[6][20]~q ;
wire \registerArray[5][20]~q ;
wire \Mux11~10_combout ;
wire \Mux11~11_combout ;
wire \Mux11~19_combout ;
wire \registerArray[21][20]~q ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \registerArray[20][20]~q ;
wire \Mux11~4_combout ;
wire \Mux11~5_combout ;
wire \Mux11~2_combout ;
wire \Mux11~3_combout ;
wire \Mux11~6_combout ;
wire \registerArray[23][20]~q ;
wire \Mux11~7_combout ;
wire \Mux11~8_combout ;
wire \Mux11~9_combout ;
wire \Mux12~7_combout ;
wire \Mux12~8_combout ;
wire \Mux12~2_combout ;
wire \Mux12~3_combout ;
wire \Mux12~6_combout ;
wire \Mux12~0_combout ;
wire \Mux12~1_combout ;
wire \Mux12~9_combout ;
wire \registerArray[1][19]~feeder_combout ;
wire \registerArray[1][19]~q ;
wire \Mux12~14_combout ;
wire \Mux12~15_combout ;
wire \Mux12~12_combout ;
wire \Mux12~13_combout ;
wire \Mux12~16_combout ;
wire \registerArray[9][19]~q ;
wire \registerArray[10][19]~q ;
wire \Mux12~10_combout ;
wire \Mux12~11_combout ;
wire \Mux12~17_combout ;
wire \Mux12~18_combout ;
wire \Mux12~19_combout ;
wire \registerArray[20][18]~feeder_combout ;
wire \registerArray[20][18]~q ;
wire \Mux13~4_combout ;
wire \Mux13~5_combout ;
wire \Mux13~6_combout ;
wire \registerArray[23][18]~feeder_combout ;
wire \registerArray[23][18]~q ;
wire \Mux13~7_combout ;
wire \Mux13~8_combout ;
wire \registerArray[17][18]~feeder_combout ;
wire \registerArray[17][18]~q ;
wire \Mux13~0_combout ;
wire \Mux13~1_combout ;
wire \Mux13~9_combout ;
wire \Mux13~17_combout ;
wire \Mux13~18_combout ;
wire \registerArray[6][18]~q ;
wire \Mux13~10_combout ;
wire \Mux13~11_combout ;
wire \Mux13~14_combout ;
wire \Mux13~15_combout ;
wire \registerArray[10][18]~feeder_combout ;
wire \registerArray[10][18]~q ;
wire \Mux13~12_combout ;
wire \Mux13~13_combout ;
wire \Mux13~16_combout ;
wire \Mux13~19_combout ;
wire \registerArray[13][17]~feeder_combout ;
wire \registerArray[13][17]~q ;
wire \Mux14~17_combout ;
wire \Mux14~18_combout ;
wire \Mux14~11_combout ;
wire \registerArray[3][17]~q ;
wire \Mux14~14_combout ;
wire \Mux14~15_combout ;
wire \registerArray[4][17]~feeder_combout ;
wire \registerArray[4][17]~q ;
wire \Mux14~12_combout ;
wire \Mux14~13_combout ;
wire \Mux14~16_combout ;
wire \Mux14~19_combout ;
wire \registerArray[27][17]~q ;
wire \Mux14~7_combout ;
wire \Mux14~8_combout ;
wire \registerArray[17][17]~feeder_combout ;
wire \registerArray[17][17]~q ;
wire \Mux14~0_combout ;
wire \Mux14~1_combout ;
wire \registerArray[22][17]~q ;
wire \registerArray[26][17]~feeder_combout ;
wire \registerArray[26][17]~q ;
wire \Mux14~2_combout ;
wire \Mux14~3_combout ;
wire \Mux14~6_combout ;
wire \Mux14~9_combout ;
wire \registerArray[6][0]~q ;
wire \registerArray[5][0]~feeder_combout ;
wire \registerArray[5][0]~q ;
wire \Mux31~10_combout ;
wire \Mux31~11_combout ;
wire \registerArray[8][0]~q ;
wire \Mux31~12_combout ;
wire \Mux31~13_combout ;
wire \Mux31~14_combout ;
wire \Mux31~15_combout ;
wire \Mux31~16_combout ;
wire \Mux31~17_combout ;
wire \Mux31~18_combout ;
wire \Mux31~19_combout ;
wire \registerArray[23][0]~feeder_combout ;
wire \registerArray[23][0]~q ;
wire \Mux31~7_combout ;
wire \Mux31~8_combout ;
wire \registerArray[20][0]~feeder_combout ;
wire \registerArray[20][0]~q ;
wire \Mux31~4_combout ;
wire \Mux31~5_combout ;
wire \Mux31~2_combout ;
wire \registerArray[26][0]~feeder_combout ;
wire \registerArray[26][0]~q ;
wire \Mux31~3_combout ;
wire \Mux31~6_combout ;
wire \registerArray[21][0]~feeder_combout ;
wire \registerArray[21][0]~q ;
wire \Mux31~0_combout ;
wire \Mux31~1_combout ;
wire \Mux31~9_combout ;


// Location: FF_X66_Y38_N25
dffeas \registerArray[9][31] (
	.clk(clk),
	.d(\registerArray[9][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][31] .is_wysiwyg = "true";
defparam \registerArray[9][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y43_N23
dffeas \registerArray[1][31] (
	.clk(clk),
	.d(\registerArray[1][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][31] .is_wysiwyg = "true";
defparam \registerArray[1][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N27
dffeas \registerArray[10][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][30] .is_wysiwyg = "true";
defparam \registerArray[10][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N23
dffeas \registerArray[6][30] (
	.clk(clk),
	.d(\registerArray[6][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][30] .is_wysiwyg = "true";
defparam \registerArray[6][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N21
dffeas \registerArray[26][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][30] .is_wysiwyg = "true";
defparam \registerArray[26][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N17
dffeas \registerArray[24][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][29] .is_wysiwyg = "true";
defparam \registerArray[24][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N3
dffeas \registerArray[20][29] (
	.clk(clk),
	.d(\registerArray[20][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][29] .is_wysiwyg = "true";
defparam \registerArray[20][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y38_N15
dffeas \registerArray[9][29] (
	.clk(clk),
	.d(\registerArray[9][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][29] .is_wysiwyg = "true";
defparam \registerArray[9][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N1
dffeas \registerArray[10][29] (
	.clk(clk),
	.d(\registerArray[10][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][29] .is_wysiwyg = "true";
defparam \registerArray[10][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N21
dffeas \registerArray[5][28] (
	.clk(clk),
	.d(\registerArray[5][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][28] .is_wysiwyg = "true";
defparam \registerArray[5][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N12
cycloneive_lcell_comb \Mux35~14 (
// Equation(s):
// \Mux35~14_combout  = (cuifregT_3 & (((\registerArray[24][28]~q ) # (cuifregT_2)))) # (!cuifregT_3 & (\registerArray[16][28]~q  & ((!cuifregT_2))))

	.dataa(\registerArray[16][28]~q ),
	.datab(\registerArray[24][28]~q ),
	.datac(cuifregT_3),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux35~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~14 .lut_mask = 16'hF0CA;
defparam \Mux35~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y34_N23
dffeas \registerArray[16][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][27] .is_wysiwyg = "true";
defparam \registerArray[16][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N22
cycloneive_lcell_comb \Mux36~14 (
// Equation(s):
// \Mux36~14_combout  = (cuifregT_2 & ((\registerArray[20][27]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[16][27]~q  & !cuifregT_3))))

	.dataa(cuifregT_2),
	.datab(\registerArray[20][27]~q ),
	.datac(\registerArray[16][27]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux36~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~14 .lut_mask = 16'hAAD8;
defparam \Mux36~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N17
dffeas \registerArray[3][26] (
	.clk(clk),
	.d(\registerArray[3][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][26] .is_wysiwyg = "true";
defparam \registerArray[3][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y37_N27
dffeas \registerArray[23][26] (
	.clk(clk),
	.d(\registerArray[23][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][26] .is_wysiwyg = "true";
defparam \registerArray[23][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N9
dffeas \registerArray[26][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][25] .is_wysiwyg = "true";
defparam \registerArray[26][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N15
dffeas \registerArray[22][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][25] .is_wysiwyg = "true";
defparam \registerArray[22][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N25
dffeas \registerArray[20][24] (
	.clk(clk),
	.d(\registerArray[20][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][24] .is_wysiwyg = "true";
defparam \registerArray[20][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N21
dffeas \registerArray[5][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][24] .is_wysiwyg = "true";
defparam \registerArray[5][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N9
dffeas \registerArray[12][24] (
	.clk(clk),
	.d(\registerArray[12][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][24] .is_wysiwyg = "true";
defparam \registerArray[12][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N29
dffeas \registerArray[26][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][23] .is_wysiwyg = "true";
defparam \registerArray[26][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N13
dffeas \registerArray[20][23] (
	.clk(clk),
	.d(\registerArray[20][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][23] .is_wysiwyg = "true";
defparam \registerArray[20][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y43_N31
dffeas \registerArray[10][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][21] .is_wysiwyg = "true";
defparam \registerArray[10][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y40_N17
dffeas \registerArray[26][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][21] .is_wysiwyg = "true";
defparam \registerArray[26][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y40_N7
dffeas \registerArray[22][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][21] .is_wysiwyg = "true";
defparam \registerArray[22][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y41_N5
dffeas \registerArray[27][21] (
	.clk(clk),
	.d(\registerArray[27][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][21] .is_wysiwyg = "true";
defparam \registerArray[27][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y44_N9
dffeas \registerArray[10][20] (
	.clk(clk),
	.d(\registerArray[10][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][20] .is_wysiwyg = "true";
defparam \registerArray[10][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y42_N23
dffeas \registerArray[3][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][20] .is_wysiwyg = "true";
defparam \registerArray[3][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N29
dffeas \registerArray[5][5] (
	.clk(clk),
	.d(\registerArray[5][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][5] .is_wysiwyg = "true";
defparam \registerArray[5][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y42_N9
dffeas \registerArray[11][5] (
	.clk(clk),
	.d(\registerArray[11][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][5] .is_wysiwyg = "true";
defparam \registerArray[11][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N19
dffeas \registerArray[5][19] (
	.clk(clk),
	.d(\registerArray[5][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][19] .is_wysiwyg = "true";
defparam \registerArray[5][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y43_N21
dffeas \registerArray[13][19] (
	.clk(clk),
	.d(\registerArray[13][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][19] .is_wysiwyg = "true";
defparam \registerArray[13][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y40_N3
dffeas \registerArray[24][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][19] .is_wysiwyg = "true";
defparam \registerArray[24][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N23
dffeas \registerArray[20][19] (
	.clk(clk),
	.d(\registerArray[20][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][19] .is_wysiwyg = "true";
defparam \registerArray[20][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y31_N9
dffeas \registerArray[5][18] (
	.clk(clk),
	.d(\registerArray[5][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][18] .is_wysiwyg = "true";
defparam \registerArray[5][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y42_N5
dffeas \registerArray[3][18] (
	.clk(clk),
	.d(Mux502),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][18] .is_wysiwyg = "true";
defparam \registerArray[3][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y42_N3
dffeas \registerArray[2][18] (
	.clk(clk),
	.d(\registerArray[2][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][18] .is_wysiwyg = "true";
defparam \registerArray[2][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y42_N15
dffeas \registerArray[13][18] (
	.clk(clk),
	.d(\registerArray[13][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][18] .is_wysiwyg = "true";
defparam \registerArray[13][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N13
dffeas \registerArray[26][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][18] .is_wysiwyg = "true";
defparam \registerArray[26][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N31
dffeas \registerArray[10][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][17] .is_wysiwyg = "true";
defparam \registerArray[10][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N31
dffeas \registerArray[20][17] (
	.clk(clk),
	.d(\registerArray[20][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][17] .is_wysiwyg = "true";
defparam \registerArray[20][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y40_N23
dffeas \registerArray[21][16] (
	.clk(clk),
	.d(\registerArray[21][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][16] .is_wysiwyg = "true";
defparam \registerArray[21][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y43_N19
dffeas \registerArray[24][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][16] .is_wysiwyg = "true";
defparam \registerArray[24][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N23
dffeas \registerArray[16][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][16] .is_wysiwyg = "true";
defparam \registerArray[16][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N22
cycloneive_lcell_comb \Mux47~4 (
// Equation(s):
// \Mux47~4_combout  = (cuifregT_3 & ((\registerArray[24][16]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[16][16]~q  & !cuifregT_2))))

	.dataa(\registerArray[24][16]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[16][16]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux47~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~4 .lut_mask = 16'hCCB8;
defparam \Mux47~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y40_N31
dffeas \registerArray[23][16] (
	.clk(clk),
	.d(\registerArray[23][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][16] .is_wysiwyg = "true";
defparam \registerArray[23][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y31_N15
dffeas \registerArray[5][16] (
	.clk(clk),
	.d(\registerArray[5][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][16] .is_wysiwyg = "true";
defparam \registerArray[5][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N21
dffeas \registerArray[3][16] (
	.clk(clk),
	.d(\registerArray[3][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][16] .is_wysiwyg = "true";
defparam \registerArray[3][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y37_N27
dffeas \registerArray[9][15] (
	.clk(clk),
	.d(\registerArray[9][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][15] .is_wysiwyg = "true";
defparam \registerArray[9][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N7
dffeas \registerArray[10][15] (
	.clk(clk),
	.d(\registerArray[10][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][15] .is_wysiwyg = "true";
defparam \registerArray[10][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N31
dffeas \registerArray[19][15] (
	.clk(clk),
	.d(\registerArray[19][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][15] .is_wysiwyg = "true";
defparam \registerArray[19][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N27
dffeas \registerArray[10][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][14] .is_wysiwyg = "true";
defparam \registerArray[10][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y31_N7
dffeas \registerArray[5][14] (
	.clk(clk),
	.d(\registerArray[5][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][14] .is_wysiwyg = "true";
defparam \registerArray[5][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y31_N13
dffeas \registerArray[5][13] (
	.clk(clk),
	.d(\registerArray[5][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][13] .is_wysiwyg = "true";
defparam \registerArray[5][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y37_N1
dffeas \registerArray[24][13] (
	.clk(clk),
	.d(\registerArray[24][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][13] .is_wysiwyg = "true";
defparam \registerArray[24][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y39_N5
dffeas \registerArray[20][13] (
	.clk(clk),
	.d(\registerArray[20][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][13] .is_wysiwyg = "true";
defparam \registerArray[20][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y42_N13
dffeas \registerArray[1][12] (
	.clk(clk),
	.d(\registerArray[1][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][12] .is_wysiwyg = "true";
defparam \registerArray[1][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y42_N27
dffeas \registerArray[21][12] (
	.clk(clk),
	.d(\registerArray[21][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][12] .is_wysiwyg = "true";
defparam \registerArray[21][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N1
dffeas \registerArray[22][12] (
	.clk(clk),
	.d(\registerArray[22][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][12] .is_wysiwyg = "true";
defparam \registerArray[22][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N7
dffeas \registerArray[10][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][10] .is_wysiwyg = "true";
defparam \registerArray[10][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y43_N27
dffeas \registerArray[3][10] (
	.clk(clk),
	.d(\registerArray[3][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][10] .is_wysiwyg = "true";
defparam \registerArray[3][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y40_N17
dffeas \registerArray[21][10] (
	.clk(clk),
	.d(Mux582),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][10] .is_wysiwyg = "true";
defparam \registerArray[21][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y43_N31
dffeas \registerArray[23][10] (
	.clk(clk),
	.d(\registerArray[23][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][10] .is_wysiwyg = "true";
defparam \registerArray[23][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N27
dffeas \registerArray[16][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][9] .is_wysiwyg = "true";
defparam \registerArray[16][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N26
cycloneive_lcell_comb \Mux54~14 (
// Equation(s):
// \Mux54~14_combout  = (cuifregT_2 & ((\registerArray[20][9]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[16][9]~q  & !cuifregT_3))))

	.dataa(cuifregT_2),
	.datab(\registerArray[20][9]~q ),
	.datac(\registerArray[16][9]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux54~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~14 .lut_mask = 16'hAAD8;
defparam \Mux54~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y30_N13
dffeas \registerArray[5][8] (
	.clk(clk),
	.d(\registerArray[5][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][8] .is_wysiwyg = "true";
defparam \registerArray[5][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N25
dffeas \registerArray[22][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][8] .is_wysiwyg = "true";
defparam \registerArray[22][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N31
dffeas \registerArray[26][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][8] .is_wysiwyg = "true";
defparam \registerArray[26][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N23
dffeas \registerArray[24][8] (
	.clk(clk),
	.d(\registerArray[24][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][8] .is_wysiwyg = "true";
defparam \registerArray[24][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N26
cycloneive_lcell_comb \Mux55~14 (
// Equation(s):
// \Mux55~14_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[24][8]~q )) # (!cuifregT_3 & ((\registerArray[16][8]~q )))))

	.dataa(\registerArray[24][8]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[16][8]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux55~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~14 .lut_mask = 16'hEE30;
defparam \Mux55~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N23
dffeas \registerArray[10][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][7] .is_wysiwyg = "true";
defparam \registerArray[10][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N7
dffeas \registerArray[3][7] (
	.clk(clk),
	.d(\registerArray[3][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][7] .is_wysiwyg = "true";
defparam \registerArray[3][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y35_N27
dffeas \registerArray[1][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][7] .is_wysiwyg = "true";
defparam \registerArray[1][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N26
cycloneive_lcell_comb \Mux56~4 (
// Equation(s):
// \Mux56~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][7]~q )) # (!cuifregT_1 & ((\registerArray[1][7]~q )))))

	.dataa(\registerArray[3][7]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[1][7]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux56~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~4 .lut_mask = 16'hB800;
defparam \Mux56~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N27
dffeas \registerArray[22][7] (
	.clk(clk),
	.d(\registerArray[22][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][7] .is_wysiwyg = "true";
defparam \registerArray[22][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y30_N31
dffeas \registerArray[6][6] (
	.clk(clk),
	.d(\registerArray[6][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][6] .is_wysiwyg = "true";
defparam \registerArray[6][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N23
dffeas \registerArray[4][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][6] .is_wysiwyg = "true";
defparam \registerArray[4][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N8
cycloneive_lcell_comb \Mux30~7 (
// Equation(s):
// \Mux30~7_combout  = (cuifregS_2 & (((\registerArray[23][1]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[19][1]~q  & ((!cuifregS_3))))

	.dataa(\registerArray[19][1]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[23][1]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux30~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~7 .lut_mask = 16'hCCE2;
defparam \Mux30~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N31
dffeas \registerArray[10][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][1] .is_wysiwyg = "true";
defparam \registerArray[10][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N30
cycloneive_lcell_comb \Mux30~10 (
// Equation(s):
// \Mux30~10_combout  = (cuifregS_1 & ((cuifregS_0) # ((\registerArray[10][1]~q )))) # (!cuifregS_1 & (!cuifregS_0 & ((\registerArray[8][1]~q ))))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\registerArray[10][1]~q ),
	.datad(\registerArray[8][1]~q ),
	.cin(gnd),
	.combout(\Mux30~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~10 .lut_mask = 16'hB9A8;
defparam \Mux30~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N1
dffeas \registerArray[17][3] (
	.clk(clk),
	.d(\registerArray[17][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][3] .is_wysiwyg = "true";
defparam \registerArray[17][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N27
dffeas \registerArray[26][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][3] .is_wysiwyg = "true";
defparam \registerArray[26][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N26
cycloneive_lcell_comb \Mux28~2 (
// Equation(s):
// \Mux28~2_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & ((\registerArray[26][3]~q ))) # (!cuifregS_3 & (\registerArray[18][3]~q ))))

	.dataa(\registerArray[18][3]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[26][3]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux28~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~2 .lut_mask = 16'hFC22;
defparam \Mux28~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N24
cycloneive_lcell_comb \Mux23~2 (
// Equation(s):
// \Mux23~2_combout  = (cuifregS_2 & (((\registerArray[22][8]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[18][8]~q  & ((!cuifregS_3))))

	.dataa(\registerArray[18][8]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[22][8]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux23~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~2 .lut_mask = 16'hCCE2;
defparam \Mux23~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N30
cycloneive_lcell_comb \Mux23~3 (
// Equation(s):
// \Mux23~3_combout  = (cuifregS_3 & ((\Mux23~2_combout  & (\registerArray[30][8]~q )) # (!\Mux23~2_combout  & ((\registerArray[26][8]~q ))))) # (!cuifregS_3 & (((\Mux23~2_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[30][8]~q ),
	.datac(\registerArray[26][8]~q ),
	.datad(\Mux23~2_combout ),
	.cin(gnd),
	.combout(\Mux23~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~3 .lut_mask = 16'hDDA0;
defparam \Mux23~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N22
cycloneive_lcell_comb \Mux24~10 (
// Equation(s):
// \Mux24~10_combout  = (cuifregS_1 & ((cuifregS_0) # ((\registerArray[10][7]~q )))) # (!cuifregS_1 & (!cuifregS_0 & ((\registerArray[8][7]~q ))))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\registerArray[10][7]~q ),
	.datad(\registerArray[8][7]~q ),
	.cin(gnd),
	.combout(\Mux24~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~10 .lut_mask = 16'hB9A8;
defparam \Mux24~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N24
cycloneive_lcell_comb \Mux24~14 (
// Equation(s):
// \Mux24~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][7]~q ))) # (!cuifregS_1 & (\registerArray[1][7]~q ))))

	.dataa(\registerArray[1][7]~q ),
	.datab(\registerArray[3][7]~q ),
	.datac(cuifregS_1),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux24~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~14 .lut_mask = 16'hCA00;
defparam \Mux24~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N10
cycloneive_lcell_comb \Mux24~15 (
// Equation(s):
// \Mux24~15_combout  = (\Mux24~14_combout ) # ((\registerArray[2][7]~q  & (!cuifregS_0 & cuifregS_1)))

	.dataa(\registerArray[2][7]~q ),
	.datab(cuifregS_0),
	.datac(cuifregS_1),
	.datad(\Mux24~14_combout ),
	.cin(gnd),
	.combout(\Mux24~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~15 .lut_mask = 16'hFF20;
defparam \Mux24~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N22
cycloneive_lcell_comb \Mux26~12 (
// Equation(s):
// \Mux26~12_combout  = (cuifregS_0 & ((\registerArray[5][5]~q ) # ((cuifregS_1)))) # (!cuifregS_0 & (((\registerArray[4][5]~q  & !cuifregS_1))))

	.dataa(\registerArray[5][5]~q ),
	.datab(\registerArray[4][5]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux26~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~12 .lut_mask = 16'hF0AC;
defparam \Mux26~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N8
cycloneive_lcell_comb \Mux26~13 (
// Equation(s):
// \Mux26~13_combout  = (\Mux26~12_combout  & ((\registerArray[7][5]~q ) # ((!cuifregS_1)))) # (!\Mux26~12_combout  & (((\registerArray[6][5]~q  & cuifregS_1))))

	.dataa(\registerArray[7][5]~q ),
	.datab(\registerArray[6][5]~q ),
	.datac(\Mux26~12_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux26~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~13 .lut_mask = 16'hACF0;
defparam \Mux26~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N16
cycloneive_lcell_comb \Mux15~4 (
// Equation(s):
// \Mux15~4_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[20][16]~q ))) # (!cuifregS_2 & (\registerArray[16][16]~q ))))

	.dataa(\registerArray[16][16]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[20][16]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux15~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~4 .lut_mask = 16'hFC22;
defparam \Mux15~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N18
cycloneive_lcell_comb \Mux15~5 (
// Equation(s):
// \Mux15~5_combout  = (cuifregS_3 & ((\Mux15~4_combout  & (\registerArray[28][16]~q )) # (!\Mux15~4_combout  & ((\registerArray[24][16]~q ))))) # (!cuifregS_3 & (((\Mux15~4_combout ))))

	.dataa(\registerArray[28][16]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[24][16]~q ),
	.datad(\Mux15~4_combout ),
	.cin(gnd),
	.combout(\Mux15~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~5 .lut_mask = 16'hBBC0;
defparam \Mux15~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N4
cycloneive_lcell_comb \Mux16~14 (
// Equation(s):
// \Mux16~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][15]~q ))) # (!cuifregS_1 & (\registerArray[1][15]~q ))))

	.dataa(\registerArray[1][15]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[3][15]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux16~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~14 .lut_mask = 16'hC088;
defparam \Mux16~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N12
cycloneive_lcell_comb \Mux16~15 (
// Equation(s):
// \Mux16~15_combout  = (\Mux16~14_combout ) # ((\registerArray[2][15]~q  & (cuifregS_1 & !cuifregS_0)))

	.dataa(\Mux16~14_combout ),
	.datab(\registerArray[2][15]~q ),
	.datac(cuifregS_1),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux16~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~15 .lut_mask = 16'hAAEA;
defparam \Mux16~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N26
cycloneive_lcell_comb \Mux17~12 (
// Equation(s):
// \Mux17~12_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][14]~q ))) # (!cuifregS_1 & (\registerArray[8][14]~q ))))

	.dataa(\registerArray[8][14]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[10][14]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux17~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~12 .lut_mask = 16'hFC22;
defparam \Mux17~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N12
cycloneive_lcell_comb \Mux19~14 (
// Equation(s):
// \Mux19~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][12]~q ))) # (!cuifregS_1 & (\registerArray[1][12]~q ))))

	.dataa(\registerArray[1][12]~q ),
	.datab(cuifregS_1),
	.datac(\registerArray[3][12]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux19~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~14 .lut_mask = 16'hE200;
defparam \Mux19~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N6
cycloneive_lcell_comb \Mux21~12 (
// Equation(s):
// \Mux21~12_combout  = (cuifregS_1 & (((\registerArray[10][10]~q ) # (cuifregS_0)))) # (!cuifregS_1 & (\registerArray[8][10]~q  & ((!cuifregS_0))))

	.dataa(cuifregS_1),
	.datab(\registerArray[8][10]~q ),
	.datac(\registerArray[10][10]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux21~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~12 .lut_mask = 16'hAAE4;
defparam \Mux21~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N14
cycloneive_lcell_comb \Mux21~14 (
// Equation(s):
// \Mux21~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][10]~q ))) # (!cuifregS_1 & (\registerArray[1][10]~q ))))

	.dataa(\registerArray[1][10]~q ),
	.datab(\registerArray[3][10]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux21~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~14 .lut_mask = 16'hC0A0;
defparam \Mux21~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N12
cycloneive_lcell_comb \Mux21~15 (
// Equation(s):
// \Mux21~15_combout  = (\Mux21~14_combout ) # ((cuifregS_1 & (!cuifregS_0 & \registerArray[2][10]~q )))

	.dataa(cuifregS_1),
	.datab(\Mux21~14_combout ),
	.datac(cuifregS_0),
	.datad(\registerArray[2][10]~q ),
	.cin(gnd),
	.combout(\Mux21~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~15 .lut_mask = 16'hCECC;
defparam \Mux21~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N16
cycloneive_lcell_comb \Mux2~4 (
// Equation(s):
// \Mux2~4_combout  = (cuifregS_3 & ((cuifregS_2) # ((\registerArray[24][29]~q )))) # (!cuifregS_3 & (!cuifregS_2 & ((\registerArray[16][29]~q ))))

	.dataa(cuifregS_3),
	.datab(cuifregS_2),
	.datac(\registerArray[24][29]~q ),
	.datad(\registerArray[16][29]~q ),
	.cin(gnd),
	.combout(\Mux2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~4 .lut_mask = 16'hB9A8;
defparam \Mux2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N14
cycloneive_lcell_comb \Mux2~5 (
// Equation(s):
// \Mux2~5_combout  = (\Mux2~4_combout  & (((\registerArray[28][29]~q ) # (!cuifregS_2)))) # (!\Mux2~4_combout  & (\registerArray[20][29]~q  & ((cuifregS_2))))

	.dataa(\registerArray[20][29]~q ),
	.datab(\registerArray[28][29]~q ),
	.datac(\Mux2~4_combout ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~5 .lut_mask = 16'hCAF0;
defparam \Mux2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N18
cycloneive_lcell_comb \Mux1~2 (
// Equation(s):
// \Mux1~2_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[22][30]~q ))) # (!cuifregS_2 & (\registerArray[18][30]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[18][30]~q ),
	.datac(\registerArray[22][30]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~2 .lut_mask = 16'hFA44;
defparam \Mux1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N20
cycloneive_lcell_comb \Mux1~3 (
// Equation(s):
// \Mux1~3_combout  = (cuifregS_3 & ((\Mux1~2_combout  & (\registerArray[30][30]~q )) # (!\Mux1~2_combout  & ((\registerArray[26][30]~q ))))) # (!cuifregS_3 & (((\Mux1~2_combout ))))

	.dataa(\registerArray[30][30]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[26][30]~q ),
	.datad(\Mux1~2_combout ),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~3 .lut_mask = 16'hBBC0;
defparam \Mux1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N26
cycloneive_lcell_comb \Mux1~12 (
// Equation(s):
// \Mux1~12_combout  = (cuifregS_1 & (((\registerArray[10][30]~q ) # (cuifregS_0)))) # (!cuifregS_1 & (\registerArray[8][30]~q  & ((!cuifregS_0))))

	.dataa(cuifregS_1),
	.datab(\registerArray[8][30]~q ),
	.datac(\registerArray[10][30]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux1~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~12 .lut_mask = 16'hAAE4;
defparam \Mux1~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N8
cycloneive_lcell_comb \Mux6~2 (
// Equation(s):
// \Mux6~2_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & ((\registerArray[26][25]~q ))) # (!cuifregS_3 & (\registerArray[18][25]~q ))))

	.dataa(\registerArray[18][25]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[26][25]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~2 .lut_mask = 16'hFC22;
defparam \Mux6~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N14
cycloneive_lcell_comb \Mux6~3 (
// Equation(s):
// \Mux6~3_combout  = (\Mux6~2_combout  & ((\registerArray[30][25]~q ) # ((!cuifregS_2)))) # (!\Mux6~2_combout  & (((\registerArray[22][25]~q  & cuifregS_2))))

	.dataa(\registerArray[30][25]~q ),
	.datab(\Mux6~2_combout ),
	.datac(\registerArray[22][25]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux6~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~3 .lut_mask = 16'hB8CC;
defparam \Mux6~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N20
cycloneive_lcell_comb \Mux7~10 (
// Equation(s):
// \Mux7~10_combout  = (cuifregS_0 & (((\registerArray[5][24]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[4][24]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[4][24]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[5][24]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux7~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~10 .lut_mask = 16'hCCE2;
defparam \Mux7~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N28
cycloneive_lcell_comb \Mux8~2 (
// Equation(s):
// \Mux8~2_combout  = (cuifregS_3 & (((\registerArray[26][23]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[18][23]~q  & ((!cuifregS_2))))

	.dataa(\registerArray[18][23]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[26][23]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux8~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~2 .lut_mask = 16'hCCE2;
defparam \Mux8~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N10
cycloneive_lcell_comb \Mux8~3 (
// Equation(s):
// \Mux8~3_combout  = (cuifregS_2 & ((\Mux8~2_combout  & (\registerArray[30][23]~q )) # (!\Mux8~2_combout  & ((\registerArray[22][23]~q ))))) # (!cuifregS_2 & (((\Mux8~2_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[30][23]~q ),
	.datac(\registerArray[22][23]~q ),
	.datad(\Mux8~2_combout ),
	.cin(gnd),
	.combout(\Mux8~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~3 .lut_mask = 16'hDDA0;
defparam \Mux8~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N16
cycloneive_lcell_comb \Mux10~2 (
// Equation(s):
// \Mux10~2_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & ((\registerArray[26][21]~q ))) # (!cuifregS_3 & (\registerArray[18][21]~q ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[18][21]~q ),
	.datac(\registerArray[26][21]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~2 .lut_mask = 16'hFA44;
defparam \Mux10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y40_N6
cycloneive_lcell_comb \Mux10~3 (
// Equation(s):
// \Mux10~3_combout  = (cuifregS_2 & ((\Mux10~2_combout  & (\registerArray[30][21]~q )) # (!\Mux10~2_combout  & ((\registerArray[22][21]~q ))))) # (!cuifregS_2 & (((\Mux10~2_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[30][21]~q ),
	.datac(\registerArray[22][21]~q ),
	.datad(\Mux10~2_combout ),
	.cin(gnd),
	.combout(\Mux10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~3 .lut_mask = 16'hDDA0;
defparam \Mux10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N30
cycloneive_lcell_comb \Mux10~10 (
// Equation(s):
// \Mux10~10_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][21]~q ))) # (!cuifregS_1 & (\registerArray[8][21]~q ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[8][21]~q ),
	.datac(\registerArray[10][21]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux10~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~10 .lut_mask = 16'hFA44;
defparam \Mux10~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N22
cycloneive_lcell_comb \Mux11~14 (
// Equation(s):
// \Mux11~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][20]~q ))) # (!cuifregS_1 & (\registerArray[1][20]~q ))))

	.dataa(\registerArray[1][20]~q ),
	.datab(cuifregS_1),
	.datac(\registerArray[3][20]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux11~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~14 .lut_mask = 16'hE200;
defparam \Mux11~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N2
cycloneive_lcell_comb \Mux11~15 (
// Equation(s):
// \Mux11~15_combout  = (\Mux11~14_combout ) # ((\registerArray[2][20]~q  & (cuifregS_1 & !cuifregS_0)))

	.dataa(\Mux11~14_combout ),
	.datab(\registerArray[2][20]~q ),
	.datac(cuifregS_1),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux11~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~15 .lut_mask = 16'hAAEA;
defparam \Mux11~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N2
cycloneive_lcell_comb \Mux12~4 (
// Equation(s):
// \Mux12~4_combout  = (cuifregS_3 & ((cuifregS_2) # ((\registerArray[24][19]~q )))) # (!cuifregS_3 & (!cuifregS_2 & ((\registerArray[16][19]~q ))))

	.dataa(cuifregS_3),
	.datab(cuifregS_2),
	.datac(\registerArray[24][19]~q ),
	.datad(\registerArray[16][19]~q ),
	.cin(gnd),
	.combout(\Mux12~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~4 .lut_mask = 16'hB9A8;
defparam \Mux12~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N26
cycloneive_lcell_comb \Mux12~5 (
// Equation(s):
// \Mux12~5_combout  = (cuifregS_2 & ((\Mux12~4_combout  & ((\registerArray[28][19]~q ))) # (!\Mux12~4_combout  & (\registerArray[20][19]~q )))) # (!cuifregS_2 & (((\Mux12~4_combout ))))

	.dataa(\registerArray[20][19]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[28][19]~q ),
	.datad(\Mux12~4_combout ),
	.cin(gnd),
	.combout(\Mux12~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~5 .lut_mask = 16'hF388;
defparam \Mux12~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N14
cycloneive_lcell_comb \Mux13~2 (
// Equation(s):
// \Mux13~2_combout  = (cuifregS_2 & (((\registerArray[22][18]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[18][18]~q  & ((!cuifregS_3))))

	.dataa(cuifregS_2),
	.datab(\registerArray[18][18]~q ),
	.datac(\registerArray[22][18]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux13~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~2 .lut_mask = 16'hAAE4;
defparam \Mux13~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N12
cycloneive_lcell_comb \Mux13~3 (
// Equation(s):
// \Mux13~3_combout  = (cuifregS_3 & ((\Mux13~2_combout  & (\registerArray[30][18]~q )) # (!\Mux13~2_combout  & ((\registerArray[26][18]~q ))))) # (!cuifregS_3 & (((\Mux13~2_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[30][18]~q ),
	.datac(\registerArray[26][18]~q ),
	.datad(\Mux13~2_combout ),
	.cin(gnd),
	.combout(\Mux13~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~3 .lut_mask = 16'hDDA0;
defparam \Mux13~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N10
cycloneive_lcell_comb \Mux14~4 (
// Equation(s):
// \Mux14~4_combout  = (cuifregS_3 & ((cuifregS_2) # ((\registerArray[24][17]~q )))) # (!cuifregS_3 & (!cuifregS_2 & ((\registerArray[16][17]~q ))))

	.dataa(cuifregS_3),
	.datab(cuifregS_2),
	.datac(\registerArray[24][17]~q ),
	.datad(\registerArray[16][17]~q ),
	.cin(gnd),
	.combout(\Mux14~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~4 .lut_mask = 16'hB9A8;
defparam \Mux14~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N6
cycloneive_lcell_comb \Mux14~5 (
// Equation(s):
// \Mux14~5_combout  = (\Mux14~4_combout  & (((\registerArray[28][17]~q ) # (!cuifregS_2)))) # (!\Mux14~4_combout  & (\registerArray[20][17]~q  & ((cuifregS_2))))

	.dataa(\registerArray[20][17]~q ),
	.datab(\registerArray[28][17]~q ),
	.datac(\Mux14~4_combout ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux14~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~5 .lut_mask = 16'hCAF0;
defparam \Mux14~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N30
cycloneive_lcell_comb \Mux14~10 (
// Equation(s):
// \Mux14~10_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][17]~q ))) # (!cuifregS_1 & (\registerArray[8][17]~q ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[8][17]~q ),
	.datac(\registerArray[10][17]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux14~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~10 .lut_mask = 16'hFA44;
defparam \Mux14~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N24
cycloneive_lcell_comb \registerArray[9][31]~feeder (
// Equation(s):
// \registerArray[9][31]~feeder_combout  = \Mux37~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux372),
	.cin(gnd),
	.combout(\registerArray[9][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[9][31]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[9][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N22
cycloneive_lcell_comb \registerArray[1][31]~feeder (
// Equation(s):
// \registerArray[1][31]~feeder_combout  = \Mux37~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux372),
	.cin(gnd),
	.combout(\registerArray[1][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[1][31]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[1][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N22
cycloneive_lcell_comb \registerArray[6][30]~feeder (
// Equation(s):
// \registerArray[6][30]~feeder_combout  = \Mux38~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux382),
	.cin(gnd),
	.combout(\registerArray[6][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[6][30]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[6][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N0
cycloneive_lcell_comb \registerArray[10][29]~feeder (
// Equation(s):
// \registerArray[10][29]~feeder_combout  = \Mux39~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux392),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[10][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[10][29]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[10][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N14
cycloneive_lcell_comb \registerArray[9][29]~feeder (
// Equation(s):
// \registerArray[9][29]~feeder_combout  = \Mux39~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux392),
	.cin(gnd),
	.combout(\registerArray[9][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[9][29]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[9][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N2
cycloneive_lcell_comb \registerArray[20][29]~feeder (
// Equation(s):
// \registerArray[20][29]~feeder_combout  = \Mux39~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux392),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[20][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[20][29]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[20][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N20
cycloneive_lcell_comb \registerArray[5][28]~feeder (
// Equation(s):
// \registerArray[5][28]~feeder_combout  = \Mux40~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux402),
	.cin(gnd),
	.combout(\registerArray[5][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[5][28]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[5][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N26
cycloneive_lcell_comb \registerArray[23][26]~feeder (
// Equation(s):
// \registerArray[23][26]~feeder_combout  = \Mux42~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux422),
	.cin(gnd),
	.combout(\registerArray[23][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[23][26]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[23][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N16
cycloneive_lcell_comb \registerArray[3][26]~feeder (
// Equation(s):
// \registerArray[3][26]~feeder_combout  = \Mux42~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux422),
	.cin(gnd),
	.combout(\registerArray[3][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[3][26]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[3][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N8
cycloneive_lcell_comb \registerArray[12][24]~feeder (
// Equation(s):
// \registerArray[12][24]~feeder_combout  = \Mux44~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux442),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[12][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[12][24]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[12][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N24
cycloneive_lcell_comb \registerArray[20][24]~feeder (
// Equation(s):
// \registerArray[20][24]~feeder_combout  = \Mux44~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux442),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[20][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[20][24]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[20][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N12
cycloneive_lcell_comb \registerArray[20][23]~feeder (
// Equation(s):
// \registerArray[20][23]~feeder_combout  = \Mux45~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux452),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[20][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[20][23]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[20][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N4
cycloneive_lcell_comb \registerArray[27][21]~feeder (
// Equation(s):
// \registerArray[27][21]~feeder_combout  = \Mux47~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux472),
	.cin(gnd),
	.combout(\registerArray[27][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[27][21]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[27][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y44_N8
cycloneive_lcell_comb \registerArray[10][20]~feeder (
// Equation(s):
// \registerArray[10][20]~feeder_combout  = \Mux48~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux482),
	.cin(gnd),
	.combout(\registerArray[10][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[10][20]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[10][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N28
cycloneive_lcell_comb \registerArray[5][5]~feeder (
// Equation(s):
// \registerArray[5][5]~feeder_combout  = \Mux63~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux632),
	.cin(gnd),
	.combout(\registerArray[5][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[5][5]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[5][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N8
cycloneive_lcell_comb \registerArray[11][5]~feeder (
// Equation(s):
// \registerArray[11][5]~feeder_combout  = \Mux63~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux632),
	.cin(gnd),
	.combout(\registerArray[11][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[11][5]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[11][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N18
cycloneive_lcell_comb \registerArray[5][19]~feeder (
// Equation(s):
// \registerArray[5][19]~feeder_combout  = \Mux49~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux492),
	.cin(gnd),
	.combout(\registerArray[5][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[5][19]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[5][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N22
cycloneive_lcell_comb \registerArray[20][19]~feeder (
// Equation(s):
// \registerArray[20][19]~feeder_combout  = \Mux49~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux492),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[20][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[20][19]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[20][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y43_N20
cycloneive_lcell_comb \registerArray[13][19]~feeder (
// Equation(s):
// \registerArray[13][19]~feeder_combout  = \Mux49~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux492),
	.cin(gnd),
	.combout(\registerArray[13][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[13][19]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[13][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N2
cycloneive_lcell_comb \registerArray[2][18]~feeder (
// Equation(s):
// \registerArray[2][18]~feeder_combout  = \Mux50~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux502),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[2][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[2][18]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[2][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N14
cycloneive_lcell_comb \registerArray[13][18]~feeder (
// Equation(s):
// \registerArray[13][18]~feeder_combout  = \Mux50~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux502),
	.cin(gnd),
	.combout(\registerArray[13][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[13][18]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[13][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N8
cycloneive_lcell_comb \registerArray[5][18]~feeder (
// Equation(s):
// \registerArray[5][18]~feeder_combout  = \Mux50~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux502),
	.cin(gnd),
	.combout(\registerArray[5][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[5][18]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[5][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N30
cycloneive_lcell_comb \registerArray[20][17]~feeder (
// Equation(s):
// \registerArray[20][17]~feeder_combout  = \Mux51~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux512),
	.cin(gnd),
	.combout(\registerArray[20][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[20][17]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[20][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N30
cycloneive_lcell_comb \registerArray[23][16]~feeder (
// Equation(s):
// \registerArray[23][16]~feeder_combout  = \Mux52~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux522),
	.cin(gnd),
	.combout(\registerArray[23][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[23][16]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[23][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N22
cycloneive_lcell_comb \registerArray[21][16]~feeder (
// Equation(s):
// \registerArray[21][16]~feeder_combout  = \Mux52~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux522),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[21][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[21][16]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[21][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N14
cycloneive_lcell_comb \registerArray[5][16]~feeder (
// Equation(s):
// \registerArray[5][16]~feeder_combout  = \Mux52~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux522),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[5][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[5][16]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[5][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N20
cycloneive_lcell_comb \registerArray[3][16]~feeder (
// Equation(s):
// \registerArray[3][16]~feeder_combout  = \Mux52~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux522),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[3][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[3][16]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[3][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N30
cycloneive_lcell_comb \registerArray[19][15]~feeder (
// Equation(s):
// \registerArray[19][15]~feeder_combout  = \Mux53~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux532),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[19][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[19][15]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[19][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N26
cycloneive_lcell_comb \registerArray[9][15]~feeder (
// Equation(s):
// \registerArray[9][15]~feeder_combout  = \Mux53~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux532),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[9][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[9][15]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[9][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N6
cycloneive_lcell_comb \registerArray[10][15]~feeder (
// Equation(s):
// \registerArray[10][15]~feeder_combout  = \Mux53~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux532),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[10][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[10][15]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[10][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N6
cycloneive_lcell_comb \registerArray[5][14]~feeder (
// Equation(s):
// \registerArray[5][14]~feeder_combout  = \Mux54~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux542),
	.cin(gnd),
	.combout(\registerArray[5][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[5][14]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[5][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y37_N0
cycloneive_lcell_comb \registerArray[24][13]~feeder (
// Equation(s):
// \registerArray[24][13]~feeder_combout  = \Mux55~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux552),
	.cin(gnd),
	.combout(\registerArray[24][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[24][13]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[24][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N4
cycloneive_lcell_comb \registerArray[20][13]~feeder (
// Equation(s):
// \registerArray[20][13]~feeder_combout  = \Mux55~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux552),
	.cin(gnd),
	.combout(\registerArray[20][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[20][13]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[20][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N12
cycloneive_lcell_comb \registerArray[5][13]~feeder (
// Equation(s):
// \registerArray[5][13]~feeder_combout  = \Mux55~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux552),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[5][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[5][13]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[5][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y42_N12
cycloneive_lcell_comb \registerArray[1][12]~feeder (
// Equation(s):
// \registerArray[1][12]~feeder_combout  = \Mux56~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux562),
	.cin(gnd),
	.combout(\registerArray[1][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[1][12]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[1][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N0
cycloneive_lcell_comb \registerArray[22][12]~feeder (
// Equation(s):
// \registerArray[22][12]~feeder_combout  = \Mux56~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux562),
	.cin(gnd),
	.combout(\registerArray[22][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[22][12]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[22][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N26
cycloneive_lcell_comb \registerArray[21][12]~feeder (
// Equation(s):
// \registerArray[21][12]~feeder_combout  = \Mux56~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux562),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[21][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[21][12]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[21][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N30
cycloneive_lcell_comb \registerArray[23][10]~feeder (
// Equation(s):
// \registerArray[23][10]~feeder_combout  = \Mux58~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux582),
	.cin(gnd),
	.combout(\registerArray[23][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[23][10]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[23][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N26
cycloneive_lcell_comb \registerArray[3][10]~feeder (
// Equation(s):
// \registerArray[3][10]~feeder_combout  = \Mux58~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux582),
	.cin(gnd),
	.combout(\registerArray[3][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[3][10]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[3][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N12
cycloneive_lcell_comb \registerArray[5][8]~feeder (
// Equation(s):
// \registerArray[5][8]~feeder_combout  = \Mux60~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux602),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[5][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[5][8]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[5][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N22
cycloneive_lcell_comb \registerArray[24][8]~feeder (
// Equation(s):
// \registerArray[24][8]~feeder_combout  = \Mux60~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux602),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[24][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[24][8]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[24][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N6
cycloneive_lcell_comb \registerArray[3][7]~feeder (
// Equation(s):
// \registerArray[3][7]~feeder_combout  = \Mux61~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux612),
	.cin(gnd),
	.combout(\registerArray[3][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[3][7]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[3][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N26
cycloneive_lcell_comb \registerArray[22][7]~feeder (
// Equation(s):
// \registerArray[22][7]~feeder_combout  = \Mux61~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux612),
	.cin(gnd),
	.combout(\registerArray[22][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[22][7]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[22][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N30
cycloneive_lcell_comb \registerArray[6][6]~feeder (
// Equation(s):
// \registerArray[6][6]~feeder_combout  = \Mux62~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux622),
	.cin(gnd),
	.combout(\registerArray[6][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[6][6]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[6][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N0
cycloneive_lcell_comb \registerArray[17][3]~feeder (
// Equation(s):
// \registerArray[17][3]~feeder_combout  = \Mux65~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux65),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[17][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[17][3]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[17][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N18
cycloneive_lcell_comb \Mux63~9 (
// Equation(s):
// Mux63 = (cuifregT_01 & ((\Mux63~6_combout  & (\Mux63~8_combout )) # (!\Mux63~6_combout  & ((\Mux63~1_combout ))))) # (!cuifregT_01 & (((\Mux63~6_combout ))))

	.dataa(\Mux63~8_combout ),
	.datab(cuifregT_0),
	.datac(\Mux63~1_combout ),
	.datad(\Mux63~6_combout ),
	.cin(gnd),
	.combout(Mux63),
	.cout());
// synopsys translate_off
defparam \Mux63~9 .lut_mask = 16'hBBC0;
defparam \Mux63~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N6
cycloneive_lcell_comb \Mux63~19 (
// Equation(s):
// Mux631 = (cuifregT_3 & ((\Mux63~16_combout  & ((\Mux63~18_combout ))) # (!\Mux63~16_combout  & (\Mux63~11_combout )))) # (!cuifregT_3 & (((\Mux63~16_combout ))))

	.dataa(cuifregT_3),
	.datab(\Mux63~11_combout ),
	.datac(\Mux63~16_combout ),
	.datad(\Mux63~18_combout ),
	.cin(gnd),
	.combout(Mux631),
	.cout());
// synopsys translate_off
defparam \Mux63~19 .lut_mask = 16'hF858;
defparam \Mux63~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N26
cycloneive_lcell_comb \Mux32~9 (
// Equation(s):
// Mux32 = (cuifregT_01 & ((\Mux32~6_combout  & (\Mux32~8_combout )) # (!\Mux32~6_combout  & ((\Mux32~1_combout ))))) # (!cuifregT_01 & (((\Mux32~6_combout ))))

	.dataa(cuifregT_0),
	.datab(\Mux32~8_combout ),
	.datac(\Mux32~6_combout ),
	.datad(\Mux32~1_combout ),
	.cin(gnd),
	.combout(Mux32),
	.cout());
// synopsys translate_off
defparam \Mux32~9 .lut_mask = 16'hDAD0;
defparam \Mux32~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N2
cycloneive_lcell_comb \Mux32~19 (
// Equation(s):
// Mux321 = (cuifregT_2 & ((\Mux32~16_combout  & ((\Mux32~18_combout ))) # (!\Mux32~16_combout  & (\Mux32~11_combout )))) # (!cuifregT_2 & (((\Mux32~16_combout ))))

	.dataa(\Mux32~11_combout ),
	.datab(cuifregT_2),
	.datac(\Mux32~18_combout ),
	.datad(\Mux32~16_combout ),
	.cin(gnd),
	.combout(Mux321),
	.cout());
// synopsys translate_off
defparam \Mux32~19 .lut_mask = 16'hF388;
defparam \Mux32~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N26
cycloneive_lcell_comb \Mux33~9 (
// Equation(s):
// Mux33 = (cuifregT_3 & ((\Mux33~6_combout  & ((\Mux33~8_combout ))) # (!\Mux33~6_combout  & (\Mux33~1_combout )))) # (!cuifregT_3 & (\Mux33~6_combout ))

	.dataa(cuifregT_3),
	.datab(\Mux33~6_combout ),
	.datac(\Mux33~1_combout ),
	.datad(\Mux33~8_combout ),
	.cin(gnd),
	.combout(Mux33),
	.cout());
// synopsys translate_off
defparam \Mux33~9 .lut_mask = 16'hEC64;
defparam \Mux33~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N2
cycloneive_lcell_comb \Mux33~19 (
// Equation(s):
// Mux331 = (cuifregT_01 & ((\Mux33~16_combout  & (\Mux33~18_combout )) # (!\Mux33~16_combout  & ((\Mux33~11_combout ))))) # (!cuifregT_01 & (((\Mux33~16_combout ))))

	.dataa(\Mux33~18_combout ),
	.datab(cuifregT_0),
	.datac(\Mux33~11_combout ),
	.datad(\Mux33~16_combout ),
	.cin(gnd),
	.combout(Mux331),
	.cout());
// synopsys translate_off
defparam \Mux33~19 .lut_mask = 16'hBBC0;
defparam \Mux33~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N30
cycloneive_lcell_comb \Mux34~9 (
// Equation(s):
// Mux34 = (cuifregT_01 & ((\Mux34~6_combout  & (\Mux34~8_combout )) # (!\Mux34~6_combout  & ((\Mux34~1_combout ))))) # (!cuifregT_01 & (((\Mux34~6_combout ))))

	.dataa(cuifregT_0),
	.datab(\Mux34~8_combout ),
	.datac(\Mux34~1_combout ),
	.datad(\Mux34~6_combout ),
	.cin(gnd),
	.combout(Mux34),
	.cout());
// synopsys translate_off
defparam \Mux34~9 .lut_mask = 16'hDDA0;
defparam \Mux34~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N6
cycloneive_lcell_comb \Mux34~19 (
// Equation(s):
// Mux341 = (cuifregT_2 & ((\Mux34~16_combout  & ((\Mux34~18_combout ))) # (!\Mux34~16_combout  & (\Mux34~11_combout )))) # (!cuifregT_2 & (((\Mux34~16_combout ))))

	.dataa(\Mux34~11_combout ),
	.datab(cuifregT_2),
	.datac(\Mux34~18_combout ),
	.datad(\Mux34~16_combout ),
	.cin(gnd),
	.combout(Mux341),
	.cout());
// synopsys translate_off
defparam \Mux34~19 .lut_mask = 16'hF388;
defparam \Mux34~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N12
cycloneive_lcell_comb \Mux35~9 (
// Equation(s):
// Mux35 = (cuifregT_3 & ((\Mux35~6_combout  & ((\Mux35~8_combout ))) # (!\Mux35~6_combout  & (\Mux35~1_combout )))) # (!cuifregT_3 & (((\Mux35~6_combout ))))

	.dataa(\Mux35~1_combout ),
	.datab(cuifregT_3),
	.datac(\Mux35~8_combout ),
	.datad(\Mux35~6_combout ),
	.cin(gnd),
	.combout(Mux35),
	.cout());
// synopsys translate_off
defparam \Mux35~9 .lut_mask = 16'hF388;
defparam \Mux35~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N8
cycloneive_lcell_comb \Mux35~19 (
// Equation(s):
// Mux351 = (cuifregT_01 & ((\Mux35~16_combout  & (\Mux35~18_combout )) # (!\Mux35~16_combout  & ((\Mux35~11_combout ))))) # (!cuifregT_01 & (((\Mux35~16_combout ))))

	.dataa(\Mux35~18_combout ),
	.datab(cuifregT_0),
	.datac(\Mux35~16_combout ),
	.datad(\Mux35~11_combout ),
	.cin(gnd),
	.combout(Mux351),
	.cout());
// synopsys translate_off
defparam \Mux35~19 .lut_mask = 16'hBCB0;
defparam \Mux35~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N24
cycloneive_lcell_comb \Mux36~9 (
// Equation(s):
// Mux36 = (cuifregT_2 & ((\Mux36~6_combout  & ((\Mux36~8_combout ))) # (!\Mux36~6_combout  & (\Mux36~1_combout )))) # (!cuifregT_2 & (((\Mux36~6_combout ))))

	.dataa(cuifregT_2),
	.datab(\Mux36~1_combout ),
	.datac(\Mux36~8_combout ),
	.datad(\Mux36~6_combout ),
	.cin(gnd),
	.combout(Mux36),
	.cout());
// synopsys translate_off
defparam \Mux36~9 .lut_mask = 16'hF588;
defparam \Mux36~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N8
cycloneive_lcell_comb \Mux36~19 (
// Equation(s):
// Mux361 = (cuifregT_01 & ((\Mux36~16_combout  & ((\Mux36~18_combout ))) # (!\Mux36~16_combout  & (\Mux36~11_combout )))) # (!cuifregT_01 & (((\Mux36~16_combout ))))

	.dataa(\Mux36~11_combout ),
	.datab(cuifregT_0),
	.datac(\Mux36~16_combout ),
	.datad(\Mux36~18_combout ),
	.cin(gnd),
	.combout(Mux361),
	.cout());
// synopsys translate_off
defparam \Mux36~19 .lut_mask = 16'hF838;
defparam \Mux36~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N26
cycloneive_lcell_comb \Mux37~9 (
// Equation(s):
// Mux37 = (cuifregT_3 & ((\Mux37~6_combout  & (\Mux37~8_combout )) # (!\Mux37~6_combout  & ((\Mux37~1_combout ))))) # (!cuifregT_3 & (((\Mux37~6_combout ))))

	.dataa(cuifregT_3),
	.datab(\Mux37~8_combout ),
	.datac(\Mux37~6_combout ),
	.datad(\Mux37~1_combout ),
	.cin(gnd),
	.combout(Mux37),
	.cout());
// synopsys translate_off
defparam \Mux37~9 .lut_mask = 16'hDAD0;
defparam \Mux37~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N12
cycloneive_lcell_comb \Mux37~19 (
// Equation(s):
// Mux371 = (cuifregT_01 & ((\Mux37~16_combout  & ((\Mux37~18_combout ))) # (!\Mux37~16_combout  & (\Mux37~11_combout )))) # (!cuifregT_01 & (((\Mux37~16_combout ))))

	.dataa(\Mux37~11_combout ),
	.datab(\Mux37~18_combout ),
	.datac(cuifregT_0),
	.datad(\Mux37~16_combout ),
	.cin(gnd),
	.combout(Mux371),
	.cout());
// synopsys translate_off
defparam \Mux37~19 .lut_mask = 16'hCFA0;
defparam \Mux37~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N0
cycloneive_lcell_comb \Mux38~9 (
// Equation(s):
// Mux38 = (cuifregT_2 & ((\Mux38~6_combout  & (\Mux38~8_combout )) # (!\Mux38~6_combout  & ((\Mux38~1_combout ))))) # (!cuifregT_2 & (((\Mux38~6_combout ))))

	.dataa(\Mux38~8_combout ),
	.datab(cuifregT_2),
	.datac(\Mux38~1_combout ),
	.datad(\Mux38~6_combout ),
	.cin(gnd),
	.combout(Mux38),
	.cout());
// synopsys translate_off
defparam \Mux38~9 .lut_mask = 16'hBBC0;
defparam \Mux38~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N10
cycloneive_lcell_comb \Mux38~19 (
// Equation(s):
// Mux381 = (cuifregT_01 & ((\Mux38~16_combout  & (\Mux38~18_combout )) # (!\Mux38~16_combout  & ((\Mux38~11_combout ))))) # (!cuifregT_01 & (\Mux38~16_combout ))

	.dataa(cuifregT_0),
	.datab(\Mux38~16_combout ),
	.datac(\Mux38~18_combout ),
	.datad(\Mux38~11_combout ),
	.cin(gnd),
	.combout(Mux381),
	.cout());
// synopsys translate_off
defparam \Mux38~19 .lut_mask = 16'hE6C4;
defparam \Mux38~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N20
cycloneive_lcell_comb \Mux39~9 (
// Equation(s):
// Mux39 = (cuifregT_01 & ((\Mux39~6_combout  & ((\Mux39~8_combout ))) # (!\Mux39~6_combout  & (\Mux39~1_combout )))) # (!cuifregT_01 & (((\Mux39~6_combout ))))

	.dataa(\Mux39~1_combout ),
	.datab(cuifregT_0),
	.datac(\Mux39~8_combout ),
	.datad(\Mux39~6_combout ),
	.cin(gnd),
	.combout(Mux39),
	.cout());
// synopsys translate_off
defparam \Mux39~9 .lut_mask = 16'hF388;
defparam \Mux39~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N22
cycloneive_lcell_comb \Mux39~19 (
// Equation(s):
// Mux391 = (cuifregT_3 & ((\Mux39~16_combout  & (\Mux39~18_combout )) # (!\Mux39~16_combout  & ((\Mux39~11_combout ))))) # (!cuifregT_3 & (((\Mux39~16_combout ))))

	.dataa(\Mux39~18_combout ),
	.datab(cuifregT_3),
	.datac(\Mux39~11_combout ),
	.datad(\Mux39~16_combout ),
	.cin(gnd),
	.combout(Mux391),
	.cout());
// synopsys translate_off
defparam \Mux39~19 .lut_mask = 16'hBBC0;
defparam \Mux39~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N26
cycloneive_lcell_comb \Mux40~9 (
// Equation(s):
// Mux40 = (cuifregT_2 & ((\Mux40~6_combout  & (\Mux40~8_combout )) # (!\Mux40~6_combout  & ((\Mux40~1_combout ))))) # (!cuifregT_2 & (((\Mux40~6_combout ))))

	.dataa(\Mux40~8_combout ),
	.datab(cuifregT_2),
	.datac(\Mux40~1_combout ),
	.datad(\Mux40~6_combout ),
	.cin(gnd),
	.combout(Mux40),
	.cout());
// synopsys translate_off
defparam \Mux40~9 .lut_mask = 16'hBBC0;
defparam \Mux40~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N18
cycloneive_lcell_comb \Mux40~19 (
// Equation(s):
// Mux401 = (cuifregT_01 & ((\Mux40~16_combout  & ((\Mux40~18_combout ))) # (!\Mux40~16_combout  & (\Mux40~11_combout )))) # (!cuifregT_01 & (\Mux40~16_combout ))

	.dataa(cuifregT_0),
	.datab(\Mux40~16_combout ),
	.datac(\Mux40~11_combout ),
	.datad(\Mux40~18_combout ),
	.cin(gnd),
	.combout(Mux401),
	.cout());
// synopsys translate_off
defparam \Mux40~19 .lut_mask = 16'hEC64;
defparam \Mux40~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N18
cycloneive_lcell_comb \Mux41~9 (
// Equation(s):
// Mux41 = (cuifregT_3 & ((\Mux41~6_combout  & (\Mux41~8_combout )) # (!\Mux41~6_combout  & ((\Mux41~1_combout ))))) # (!cuifregT_3 & (((\Mux41~6_combout ))))

	.dataa(cuifregT_3),
	.datab(\Mux41~8_combout ),
	.datac(\Mux41~1_combout ),
	.datad(\Mux41~6_combout ),
	.cin(gnd),
	.combout(Mux41),
	.cout());
// synopsys translate_off
defparam \Mux41~9 .lut_mask = 16'hDDA0;
defparam \Mux41~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N30
cycloneive_lcell_comb \Mux41~19 (
// Equation(s):
// Mux411 = (cuifregT_01 & ((\Mux41~16_combout  & (\Mux41~18_combout )) # (!\Mux41~16_combout  & ((\Mux41~11_combout ))))) # (!cuifregT_01 & (((\Mux41~16_combout ))))

	.dataa(\Mux41~18_combout ),
	.datab(cuifregT_0),
	.datac(\Mux41~11_combout ),
	.datad(\Mux41~16_combout ),
	.cin(gnd),
	.combout(Mux411),
	.cout());
// synopsys translate_off
defparam \Mux41~19 .lut_mask = 16'hBBC0;
defparam \Mux41~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N8
cycloneive_lcell_comb \Mux42~9 (
// Equation(s):
// Mux42 = (cuifregT_2 & ((\Mux42~6_combout  & (\Mux42~8_combout )) # (!\Mux42~6_combout  & ((\Mux42~1_combout ))))) # (!cuifregT_2 & (((\Mux42~6_combout ))))

	.dataa(cuifregT_2),
	.datab(\Mux42~8_combout ),
	.datac(\Mux42~6_combout ),
	.datad(\Mux42~1_combout ),
	.cin(gnd),
	.combout(Mux42),
	.cout());
// synopsys translate_off
defparam \Mux42~9 .lut_mask = 16'hDAD0;
defparam \Mux42~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N10
cycloneive_lcell_comb \Mux42~19 (
// Equation(s):
// Mux421 = (cuifregT_01 & ((\Mux42~16_combout  & ((\Mux42~18_combout ))) # (!\Mux42~16_combout  & (\Mux42~11_combout )))) # (!cuifregT_01 & (((\Mux42~16_combout ))))

	.dataa(\Mux42~11_combout ),
	.datab(cuifregT_0),
	.datac(\Mux42~18_combout ),
	.datad(\Mux42~16_combout ),
	.cin(gnd),
	.combout(Mux421),
	.cout());
// synopsys translate_off
defparam \Mux42~19 .lut_mask = 16'hF388;
defparam \Mux42~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N2
cycloneive_lcell_comb \Mux43~9 (
// Equation(s):
// Mux43 = (cuifregT_3 & ((\Mux43~6_combout  & (\Mux43~8_combout )) # (!\Mux43~6_combout  & ((\Mux43~1_combout ))))) # (!cuifregT_3 & (((\Mux43~6_combout ))))

	.dataa(\Mux43~8_combout ),
	.datab(cuifregT_3),
	.datac(\Mux43~1_combout ),
	.datad(\Mux43~6_combout ),
	.cin(gnd),
	.combout(Mux43),
	.cout());
// synopsys translate_off
defparam \Mux43~9 .lut_mask = 16'hBBC0;
defparam \Mux43~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N4
cycloneive_lcell_comb \Mux43~19 (
// Equation(s):
// Mux431 = (\Mux43~16_combout  & (((\Mux43~18_combout )) # (!cuifregT_01))) # (!\Mux43~16_combout  & (cuifregT_01 & (\Mux43~11_combout )))

	.dataa(\Mux43~16_combout ),
	.datab(cuifregT_0),
	.datac(\Mux43~11_combout ),
	.datad(\Mux43~18_combout ),
	.cin(gnd),
	.combout(Mux431),
	.cout());
// synopsys translate_off
defparam \Mux43~19 .lut_mask = 16'hEA62;
defparam \Mux43~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N24
cycloneive_lcell_comb \Mux58~9 (
// Equation(s):
// Mux58 = (cuifregT_2 & ((\Mux58~6_combout  & (\Mux58~8_combout )) # (!\Mux58~6_combout  & ((\Mux58~1_combout ))))) # (!cuifregT_2 & (((\Mux58~6_combout ))))

	.dataa(cuifregT_2),
	.datab(\Mux58~8_combout ),
	.datac(\Mux58~1_combout ),
	.datad(\Mux58~6_combout ),
	.cin(gnd),
	.combout(Mux58),
	.cout());
// synopsys translate_off
defparam \Mux58~9 .lut_mask = 16'hDDA0;
defparam \Mux58~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N26
cycloneive_lcell_comb \Mux58~19 (
// Equation(s):
// Mux581 = (cuifregT_01 & ((\Mux58~16_combout  & (\Mux58~18_combout )) # (!\Mux58~16_combout  & ((\Mux58~11_combout ))))) # (!cuifregT_01 & (((\Mux58~16_combout ))))

	.dataa(\Mux58~18_combout ),
	.datab(cuifregT_0),
	.datac(\Mux58~16_combout ),
	.datad(\Mux58~11_combout ),
	.cin(gnd),
	.combout(Mux581),
	.cout());
// synopsys translate_off
defparam \Mux58~19 .lut_mask = 16'hBCB0;
defparam \Mux58~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N14
cycloneive_lcell_comb \Mux44~9 (
// Equation(s):
// Mux44 = (cuifregT_2 & ((\Mux44~6_combout  & (\Mux44~8_combout )) # (!\Mux44~6_combout  & ((\Mux44~1_combout ))))) # (!cuifregT_2 & (((\Mux44~6_combout ))))

	.dataa(cuifregT_2),
	.datab(\Mux44~8_combout ),
	.datac(\Mux44~1_combout ),
	.datad(\Mux44~6_combout ),
	.cin(gnd),
	.combout(Mux44),
	.cout());
// synopsys translate_off
defparam \Mux44~9 .lut_mask = 16'hDDA0;
defparam \Mux44~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N10
cycloneive_lcell_comb \Mux44~19 (
// Equation(s):
// Mux441 = (cuifregT_01 & ((\Mux44~16_combout  & (\Mux44~18_combout )) # (!\Mux44~16_combout  & ((\Mux44~11_combout ))))) # (!cuifregT_01 & (\Mux44~16_combout ))

	.dataa(cuifregT_0),
	.datab(\Mux44~16_combout ),
	.datac(\Mux44~18_combout ),
	.datad(\Mux44~11_combout ),
	.cin(gnd),
	.combout(Mux441),
	.cout());
// synopsys translate_off
defparam \Mux44~19 .lut_mask = 16'hE6C4;
defparam \Mux44~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N0
cycloneive_lcell_comb \Mux45~9 (
// Equation(s):
// Mux45 = (cuifregT_3 & ((\Mux45~6_combout  & ((\Mux45~8_combout ))) # (!\Mux45~6_combout  & (\Mux45~1_combout )))) # (!cuifregT_3 & (((\Mux45~6_combout ))))

	.dataa(\Mux45~1_combout ),
	.datab(\Mux45~8_combout ),
	.datac(cuifregT_3),
	.datad(\Mux45~6_combout ),
	.cin(gnd),
	.combout(Mux45),
	.cout());
// synopsys translate_off
defparam \Mux45~9 .lut_mask = 16'hCFA0;
defparam \Mux45~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N30
cycloneive_lcell_comb \Mux45~19 (
// Equation(s):
// Mux451 = (cuifregT_01 & ((\Mux45~16_combout  & (\Mux45~18_combout )) # (!\Mux45~16_combout  & ((\Mux45~11_combout ))))) # (!cuifregT_01 & (\Mux45~16_combout ))

	.dataa(cuifregT_0),
	.datab(\Mux45~16_combout ),
	.datac(\Mux45~18_combout ),
	.datad(\Mux45~11_combout ),
	.cin(gnd),
	.combout(Mux451),
	.cout());
// synopsys translate_off
defparam \Mux45~19 .lut_mask = 16'hE6C4;
defparam \Mux45~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N20
cycloneive_lcell_comb \Mux46~9 (
// Equation(s):
// Mux46 = (cuifregT_2 & ((\Mux46~6_combout  & (\Mux46~8_combout )) # (!\Mux46~6_combout  & ((\Mux46~1_combout ))))) # (!cuifregT_2 & (((\Mux46~6_combout ))))

	.dataa(cuifregT_2),
	.datab(\Mux46~8_combout ),
	.datac(\Mux46~1_combout ),
	.datad(\Mux46~6_combout ),
	.cin(gnd),
	.combout(Mux46),
	.cout());
// synopsys translate_off
defparam \Mux46~9 .lut_mask = 16'hDDA0;
defparam \Mux46~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N26
cycloneive_lcell_comb \Mux46~19 (
// Equation(s):
// Mux461 = (cuifregT_01 & ((\Mux46~16_combout  & ((\Mux46~18_combout ))) # (!\Mux46~16_combout  & (\Mux46~11_combout )))) # (!cuifregT_01 & (\Mux46~16_combout ))

	.dataa(cuifregT_0),
	.datab(\Mux46~16_combout ),
	.datac(\Mux46~11_combout ),
	.datad(\Mux46~18_combout ),
	.cin(gnd),
	.combout(Mux461),
	.cout());
// synopsys translate_off
defparam \Mux46~19 .lut_mask = 16'hEC64;
defparam \Mux46~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N24
cycloneive_lcell_comb \Mux47~9 (
// Equation(s):
// Mux47 = (cuifregT_01 & ((\Mux47~6_combout  & (\Mux47~8_combout )) # (!\Mux47~6_combout  & ((\Mux47~1_combout ))))) # (!cuifregT_01 & (((\Mux47~6_combout ))))

	.dataa(cuifregT_0),
	.datab(\Mux47~8_combout ),
	.datac(\Mux47~1_combout ),
	.datad(\Mux47~6_combout ),
	.cin(gnd),
	.combout(Mux47),
	.cout());
// synopsys translate_off
defparam \Mux47~9 .lut_mask = 16'hDDA0;
defparam \Mux47~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N2
cycloneive_lcell_comb \Mux47~19 (
// Equation(s):
// Mux471 = (cuifregT_3 & ((\Mux47~16_combout  & (\Mux47~18_combout )) # (!\Mux47~16_combout  & ((\Mux47~11_combout ))))) # (!cuifregT_3 & (((\Mux47~16_combout ))))

	.dataa(cuifregT_3),
	.datab(\Mux47~18_combout ),
	.datac(\Mux47~16_combout ),
	.datad(\Mux47~11_combout ),
	.cin(gnd),
	.combout(Mux471),
	.cout());
// synopsys translate_off
defparam \Mux47~19 .lut_mask = 16'hDAD0;
defparam \Mux47~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N2
cycloneive_lcell_comb \Mux48~9 (
// Equation(s):
// Mux48 = (cuifregT_2 & ((\Mux48~6_combout  & ((\Mux48~8_combout ))) # (!\Mux48~6_combout  & (\Mux48~1_combout )))) # (!cuifregT_2 & (((\Mux48~6_combout ))))

	.dataa(cuifregT_2),
	.datab(\Mux48~1_combout ),
	.datac(\Mux48~8_combout ),
	.datad(\Mux48~6_combout ),
	.cin(gnd),
	.combout(Mux48),
	.cout());
// synopsys translate_off
defparam \Mux48~9 .lut_mask = 16'hF588;
defparam \Mux48~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N6
cycloneive_lcell_comb \Mux48~19 (
// Equation(s):
// Mux481 = (cuifregT_01 & ((\Mux48~16_combout  & ((\Mux48~18_combout ))) # (!\Mux48~16_combout  & (\Mux48~11_combout )))) # (!cuifregT_01 & (((\Mux48~16_combout ))))

	.dataa(\Mux48~11_combout ),
	.datab(cuifregT_0),
	.datac(\Mux48~18_combout ),
	.datad(\Mux48~16_combout ),
	.cin(gnd),
	.combout(Mux481),
	.cout());
// synopsys translate_off
defparam \Mux48~19 .lut_mask = 16'hF388;
defparam \Mux48~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N10
cycloneive_lcell_comb \Mux49~9 (
// Equation(s):
// Mux49 = (cuifregT_3 & ((\Mux49~6_combout  & (\Mux49~8_combout )) # (!\Mux49~6_combout  & ((\Mux49~1_combout ))))) # (!cuifregT_3 & (((\Mux49~6_combout ))))

	.dataa(cuifregT_3),
	.datab(\Mux49~8_combout ),
	.datac(\Mux49~1_combout ),
	.datad(\Mux49~6_combout ),
	.cin(gnd),
	.combout(Mux49),
	.cout());
// synopsys translate_off
defparam \Mux49~9 .lut_mask = 16'hDDA0;
defparam \Mux49~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N22
cycloneive_lcell_comb \Mux49~19 (
// Equation(s):
// Mux491 = (cuifregT_01 & ((\Mux49~16_combout  & (\Mux49~18_combout )) # (!\Mux49~16_combout  & ((\Mux49~11_combout ))))) # (!cuifregT_01 & (((\Mux49~16_combout ))))

	.dataa(cuifregT_0),
	.datab(\Mux49~18_combout ),
	.datac(\Mux49~16_combout ),
	.datad(\Mux49~11_combout ),
	.cin(gnd),
	.combout(Mux491),
	.cout());
// synopsys translate_off
defparam \Mux49~19 .lut_mask = 16'hDAD0;
defparam \Mux49~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N2
cycloneive_lcell_comb \Mux50~9 (
// Equation(s):
// Mux50 = (cuifregT_2 & ((\Mux50~6_combout  & (\Mux50~8_combout )) # (!\Mux50~6_combout  & ((\Mux50~1_combout ))))) # (!cuifregT_2 & (((\Mux50~6_combout ))))

	.dataa(\Mux50~8_combout ),
	.datab(cuifregT_2),
	.datac(\Mux50~1_combout ),
	.datad(\Mux50~6_combout ),
	.cin(gnd),
	.combout(Mux50),
	.cout());
// synopsys translate_off
defparam \Mux50~9 .lut_mask = 16'hBBC0;
defparam \Mux50~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N24
cycloneive_lcell_comb \Mux50~19 (
// Equation(s):
// Mux501 = (cuifregT_01 & ((\Mux50~16_combout  & (\Mux50~18_combout )) # (!\Mux50~16_combout  & ((\Mux50~11_combout ))))) # (!cuifregT_01 & (((\Mux50~16_combout ))))

	.dataa(\Mux50~18_combout ),
	.datab(cuifregT_0),
	.datac(\Mux50~16_combout ),
	.datad(\Mux50~11_combout ),
	.cin(gnd),
	.combout(Mux501),
	.cout());
// synopsys translate_off
defparam \Mux50~19 .lut_mask = 16'hBCB0;
defparam \Mux50~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N2
cycloneive_lcell_comb \Mux51~9 (
// Equation(s):
// Mux51 = (cuifregT_3 & ((\Mux51~6_combout  & (\Mux51~8_combout )) # (!\Mux51~6_combout  & ((\Mux51~1_combout ))))) # (!cuifregT_3 & (((\Mux51~6_combout ))))

	.dataa(cuifregT_3),
	.datab(\Mux51~8_combout ),
	.datac(\Mux51~1_combout ),
	.datad(\Mux51~6_combout ),
	.cin(gnd),
	.combout(Mux51),
	.cout());
// synopsys translate_off
defparam \Mux51~9 .lut_mask = 16'hDDA0;
defparam \Mux51~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N4
cycloneive_lcell_comb \Mux51~19 (
// Equation(s):
// Mux511 = (\Mux51~16_combout  & (((\Mux51~18_combout ) # (!cuifregT_01)))) # (!\Mux51~16_combout  & (\Mux51~11_combout  & ((cuifregT_01))))

	.dataa(\Mux51~11_combout ),
	.datab(\Mux51~16_combout ),
	.datac(\Mux51~18_combout ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(Mux511),
	.cout());
// synopsys translate_off
defparam \Mux51~19 .lut_mask = 16'hE2CC;
defparam \Mux51~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N14
cycloneive_lcell_comb \Mux52~9 (
// Equation(s):
// Mux52 = (cuifregT_2 & ((\Mux52~6_combout  & (\Mux52~8_combout )) # (!\Mux52~6_combout  & ((\Mux52~1_combout ))))) # (!cuifregT_2 & (((\Mux52~6_combout ))))

	.dataa(\Mux52~8_combout ),
	.datab(cuifregT_2),
	.datac(\Mux52~6_combout ),
	.datad(\Mux52~1_combout ),
	.cin(gnd),
	.combout(Mux52),
	.cout());
// synopsys translate_off
defparam \Mux52~9 .lut_mask = 16'hBCB0;
defparam \Mux52~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N6
cycloneive_lcell_comb \Mux52~19 (
// Equation(s):
// Mux521 = (cuifregT_01 & ((\Mux52~16_combout  & (\Mux52~18_combout )) # (!\Mux52~16_combout  & ((\Mux52~11_combout ))))) # (!cuifregT_01 & (((\Mux52~16_combout ))))

	.dataa(\Mux52~18_combout ),
	.datab(cuifregT_0),
	.datac(\Mux52~11_combout ),
	.datad(\Mux52~16_combout ),
	.cin(gnd),
	.combout(Mux521),
	.cout());
// synopsys translate_off
defparam \Mux52~19 .lut_mask = 16'hBBC0;
defparam \Mux52~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N2
cycloneive_lcell_comb \Mux53~9 (
// Equation(s):
// Mux53 = (cuifregT_3 & ((\Mux53~6_combout  & (\Mux53~8_combout )) # (!\Mux53~6_combout  & ((\Mux53~1_combout ))))) # (!cuifregT_3 & (((\Mux53~6_combout ))))

	.dataa(\Mux53~8_combout ),
	.datab(cuifregT_3),
	.datac(\Mux53~1_combout ),
	.datad(\Mux53~6_combout ),
	.cin(gnd),
	.combout(Mux53),
	.cout());
// synopsys translate_off
defparam \Mux53~9 .lut_mask = 16'hBBC0;
defparam \Mux53~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N4
cycloneive_lcell_comb \Mux53~19 (
// Equation(s):
// Mux531 = (cuifregT_01 & ((\Mux53~16_combout  & (\Mux53~18_combout )) # (!\Mux53~16_combout  & ((\Mux53~11_combout ))))) # (!cuifregT_01 & (((\Mux53~16_combout ))))

	.dataa(cuifregT_0),
	.datab(\Mux53~18_combout ),
	.datac(\Mux53~11_combout ),
	.datad(\Mux53~16_combout ),
	.cin(gnd),
	.combout(Mux531),
	.cout());
// synopsys translate_off
defparam \Mux53~19 .lut_mask = 16'hDDA0;
defparam \Mux53~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N2
cycloneive_lcell_comb \Mux54~9 (
// Equation(s):
// Mux54 = (cuifregT_2 & ((\Mux54~6_combout  & (\Mux54~8_combout )) # (!\Mux54~6_combout  & ((\Mux54~1_combout ))))) # (!cuifregT_2 & (((\Mux54~6_combout ))))

	.dataa(cuifregT_2),
	.datab(\Mux54~8_combout ),
	.datac(\Mux54~1_combout ),
	.datad(\Mux54~6_combout ),
	.cin(gnd),
	.combout(Mux54),
	.cout());
// synopsys translate_off
defparam \Mux54~9 .lut_mask = 16'hDDA0;
defparam \Mux54~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N16
cycloneive_lcell_comb \Mux54~19 (
// Equation(s):
// Mux541 = (\Mux54~16_combout  & (((\Mux54~18_combout )) # (!cuifregT_01))) # (!\Mux54~16_combout  & (cuifregT_01 & (\Mux54~11_combout )))

	.dataa(\Mux54~16_combout ),
	.datab(cuifregT_0),
	.datac(\Mux54~11_combout ),
	.datad(\Mux54~18_combout ),
	.cin(gnd),
	.combout(Mux541),
	.cout());
// synopsys translate_off
defparam \Mux54~19 .lut_mask = 16'hEA62;
defparam \Mux54~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N6
cycloneive_lcell_comb \Mux55~9 (
// Equation(s):
// Mux55 = (cuifregT_3 & ((\Mux55~6_combout  & ((\Mux55~8_combout ))) # (!\Mux55~6_combout  & (\Mux55~1_combout )))) # (!cuifregT_3 & (((\Mux55~6_combout ))))

	.dataa(cuifregT_3),
	.datab(\Mux55~1_combout ),
	.datac(\Mux55~8_combout ),
	.datad(\Mux55~6_combout ),
	.cin(gnd),
	.combout(Mux55),
	.cout());
// synopsys translate_off
defparam \Mux55~9 .lut_mask = 16'hF588;
defparam \Mux55~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N24
cycloneive_lcell_comb \Mux55~19 (
// Equation(s):
// Mux551 = (\Mux55~16_combout  & ((\Mux55~18_combout ) # ((!cuifregT_01)))) # (!\Mux55~16_combout  & (((\Mux55~11_combout  & cuifregT_01))))

	.dataa(\Mux55~18_combout ),
	.datab(\Mux55~16_combout ),
	.datac(\Mux55~11_combout ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(Mux551),
	.cout());
// synopsys translate_off
defparam \Mux55~19 .lut_mask = 16'hB8CC;
defparam \Mux55~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N24
cycloneive_lcell_comb \Mux56~9 (
// Equation(s):
// Mux56 = (cuifregT_2 & ((\Mux56~6_combout  & (\Mux56~8_combout )) # (!\Mux56~6_combout  & ((\Mux56~1_combout ))))) # (!cuifregT_2 & (((\Mux56~6_combout ))))

	.dataa(cuifregT_2),
	.datab(\Mux56~8_combout ),
	.datac(\Mux56~1_combout ),
	.datad(\Mux56~6_combout ),
	.cin(gnd),
	.combout(Mux56),
	.cout());
// synopsys translate_off
defparam \Mux56~9 .lut_mask = 16'hDDA0;
defparam \Mux56~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N30
cycloneive_lcell_comb \Mux56~19 (
// Equation(s):
// Mux561 = (cuifregT_01 & ((\Mux56~16_combout  & (\Mux56~18_combout )) # (!\Mux56~16_combout  & ((\Mux56~11_combout ))))) # (!cuifregT_01 & (((\Mux56~16_combout ))))

	.dataa(cuifregT_0),
	.datab(\Mux56~18_combout ),
	.datac(\Mux56~11_combout ),
	.datad(\Mux56~16_combout ),
	.cin(gnd),
	.combout(Mux561),
	.cout());
// synopsys translate_off
defparam \Mux56~19 .lut_mask = 16'hDDA0;
defparam \Mux56~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N4
cycloneive_lcell_comb \Mux57~9 (
// Equation(s):
// Mux57 = (cuifregT_3 & ((\Mux57~6_combout  & ((\Mux57~8_combout ))) # (!\Mux57~6_combout  & (\Mux57~1_combout )))) # (!cuifregT_3 & (((\Mux57~6_combout ))))

	.dataa(cuifregT_3),
	.datab(\Mux57~1_combout ),
	.datac(\Mux57~6_combout ),
	.datad(\Mux57~8_combout ),
	.cin(gnd),
	.combout(Mux57),
	.cout());
// synopsys translate_off
defparam \Mux57~9 .lut_mask = 16'hF858;
defparam \Mux57~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N6
cycloneive_lcell_comb \Mux57~19 (
// Equation(s):
// Mux571 = (cuifregT_01 & ((\Mux57~16_combout  & ((\Mux57~18_combout ))) # (!\Mux57~16_combout  & (\Mux57~11_combout )))) # (!cuifregT_01 & (((\Mux57~16_combout ))))

	.dataa(cuifregT_0),
	.datab(\Mux57~11_combout ),
	.datac(\Mux57~18_combout ),
	.datad(\Mux57~16_combout ),
	.cin(gnd),
	.combout(Mux571),
	.cout());
// synopsys translate_off
defparam \Mux57~19 .lut_mask = 16'hF588;
defparam \Mux57~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N28
cycloneive_lcell_comb \Mux29~20 (
// Equation(s):
// Mux29 = (cuifregS_4 & (\Mux29~9_combout )) # (!cuifregS_4 & ((\Mux29~19_combout )))

	.dataa(cuifregS_4),
	.datab(gnd),
	.datac(\Mux29~9_combout ),
	.datad(\Mux29~19_combout ),
	.cin(gnd),
	.combout(Mux29),
	.cout());
// synopsys translate_off
defparam \Mux29~20 .lut_mask = 16'hF5A0;
defparam \Mux29~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N4
cycloneive_lcell_comb \Mux30~20 (
// Equation(s):
// Mux30 = (cuifregS_4 & (\Mux30~9_combout )) # (!cuifregS_4 & ((\Mux30~19_combout )))

	.dataa(gnd),
	.datab(\Mux30~9_combout ),
	.datac(cuifregS_4),
	.datad(\Mux30~19_combout ),
	.cin(gnd),
	.combout(Mux30),
	.cout());
// synopsys translate_off
defparam \Mux30~20 .lut_mask = 16'hCFC0;
defparam \Mux30~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N0
cycloneive_lcell_comb \Mux62~9 (
// Equation(s):
// Mux62 = (cuifregT_2 & ((\Mux62~6_combout  & (\Mux62~8_combout )) # (!\Mux62~6_combout  & ((\Mux62~1_combout ))))) # (!cuifregT_2 & (((\Mux62~6_combout ))))

	.dataa(cuifregT_2),
	.datab(\Mux62~8_combout ),
	.datac(\Mux62~1_combout ),
	.datad(\Mux62~6_combout ),
	.cin(gnd),
	.combout(Mux62),
	.cout());
// synopsys translate_off
defparam \Mux62~9 .lut_mask = 16'hDDA0;
defparam \Mux62~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N22
cycloneive_lcell_comb \Mux62~19 (
// Equation(s):
// Mux621 = (cuifregT_01 & ((\Mux62~16_combout  & (\Mux62~18_combout )) # (!\Mux62~16_combout  & ((\Mux62~11_combout ))))) # (!cuifregT_01 & (((\Mux62~16_combout ))))

	.dataa(\Mux62~18_combout ),
	.datab(cuifregT_0),
	.datac(\Mux62~16_combout ),
	.datad(\Mux62~11_combout ),
	.cin(gnd),
	.combout(Mux621),
	.cout());
// synopsys translate_off
defparam \Mux62~19 .lut_mask = 16'hBCB0;
defparam \Mux62~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N6
cycloneive_lcell_comb \Mux27~20 (
// Equation(s):
// Mux27 = (cuifregS_4 & ((\Mux27~9_combout ))) # (!cuifregS_4 & (\Mux27~19_combout ))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux27~19_combout ),
	.datad(\Mux27~9_combout ),
	.cin(gnd),
	.combout(Mux27),
	.cout());
// synopsys translate_off
defparam \Mux27~20 .lut_mask = 16'hFC30;
defparam \Mux27~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y43_N2
cycloneive_lcell_comb \Mux28~20 (
// Equation(s):
// Mux28 = (cuifregS_4 & (\Mux28~9_combout )) # (!cuifregS_4 & ((\Mux28~19_combout )))

	.dataa(cuifregS_4),
	.datab(gnd),
	.datac(\Mux28~9_combout ),
	.datad(\Mux28~19_combout ),
	.cin(gnd),
	.combout(Mux28),
	.cout());
// synopsys translate_off
defparam \Mux28~20 .lut_mask = 16'hF5A0;
defparam \Mux28~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N30
cycloneive_lcell_comb \Mux61~9 (
// Equation(s):
// Mux61 = (cuifregT_01 & ((\Mux61~6_combout  & (\Mux61~8_combout )) # (!\Mux61~6_combout  & ((\Mux61~1_combout ))))) # (!cuifregT_01 & (\Mux61~6_combout ))

	.dataa(cuifregT_0),
	.datab(\Mux61~6_combout ),
	.datac(\Mux61~8_combout ),
	.datad(\Mux61~1_combout ),
	.cin(gnd),
	.combout(Mux61),
	.cout());
// synopsys translate_off
defparam \Mux61~9 .lut_mask = 16'hE6C4;
defparam \Mux61~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N20
cycloneive_lcell_comb \Mux61~19 (
// Equation(s):
// Mux611 = (cuifregT_3 & ((\Mux61~16_combout  & ((\Mux61~18_combout ))) # (!\Mux61~16_combout  & (\Mux61~11_combout )))) # (!cuifregT_3 & (((\Mux61~16_combout ))))

	.dataa(cuifregT_3),
	.datab(\Mux61~11_combout ),
	.datac(\Mux61~18_combout ),
	.datad(\Mux61~16_combout ),
	.cin(gnd),
	.combout(Mux611),
	.cout());
// synopsys translate_off
defparam \Mux61~19 .lut_mask = 16'hF588;
defparam \Mux61~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N16
cycloneive_lcell_comb \Mux23~20 (
// Equation(s):
// Mux23 = (cuifregS_4 & (\Mux23~9_combout )) # (!cuifregS_4 & ((\Mux23~19_combout )))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux23~9_combout ),
	.datad(\Mux23~19_combout ),
	.cin(gnd),
	.combout(Mux23),
	.cout());
// synopsys translate_off
defparam \Mux23~20 .lut_mask = 16'hF3C0;
defparam \Mux23~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N14
cycloneive_lcell_comb \Mux24~20 (
// Equation(s):
// Mux24 = (cuifregS_4 & (\Mux24~9_combout )) # (!cuifregS_4 & ((\Mux24~19_combout )))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux24~9_combout ),
	.datad(\Mux24~19_combout ),
	.cin(gnd),
	.combout(Mux24),
	.cout());
// synopsys translate_off
defparam \Mux24~20 .lut_mask = 16'hF3C0;
defparam \Mux24~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N0
cycloneive_lcell_comb \Mux25~20 (
// Equation(s):
// Mux25 = (cuifregS_4 & (\Mux25~9_combout )) # (!cuifregS_4 & ((\Mux25~19_combout )))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux25~9_combout ),
	.datad(\Mux25~19_combout ),
	.cin(gnd),
	.combout(Mux25),
	.cout());
// synopsys translate_off
defparam \Mux25~20 .lut_mask = 16'hF3C0;
defparam \Mux25~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N12
cycloneive_lcell_comb \Mux26~20 (
// Equation(s):
// Mux26 = (cuifregS_4 & (\Mux26~9_combout )) # (!cuifregS_4 & ((\Mux26~19_combout )))

	.dataa(cuifregS_4),
	.datab(gnd),
	.datac(\Mux26~9_combout ),
	.datad(\Mux26~19_combout ),
	.cin(gnd),
	.combout(Mux26),
	.cout());
// synopsys translate_off
defparam \Mux26~20 .lut_mask = 16'hF5A0;
defparam \Mux26~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N18
cycloneive_lcell_comb \Mux60~9 (
// Equation(s):
// Mux60 = (cuifregT_01 & ((\Mux60~6_combout  & ((\Mux60~8_combout ))) # (!\Mux60~6_combout  & (\Mux60~1_combout )))) # (!cuifregT_01 & (\Mux60~6_combout ))

	.dataa(cuifregT_0),
	.datab(\Mux60~6_combout ),
	.datac(\Mux60~1_combout ),
	.datad(\Mux60~8_combout ),
	.cin(gnd),
	.combout(Mux60),
	.cout());
// synopsys translate_off
defparam \Mux60~9 .lut_mask = 16'hEC64;
defparam \Mux60~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N2
cycloneive_lcell_comb \Mux60~19 (
// Equation(s):
// Mux601 = (cuifregT_2 & ((\Mux60~16_combout  & (\Mux60~18_combout )) # (!\Mux60~16_combout  & ((\Mux60~11_combout ))))) # (!cuifregT_2 & (((\Mux60~16_combout ))))

	.dataa(\Mux60~18_combout ),
	.datab(cuifregT_2),
	.datac(\Mux60~11_combout ),
	.datad(\Mux60~16_combout ),
	.cin(gnd),
	.combout(Mux601),
	.cout());
// synopsys translate_off
defparam \Mux60~19 .lut_mask = 16'hBBC0;
defparam \Mux60~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N16
cycloneive_lcell_comb \Mux15~20 (
// Equation(s):
// Mux15 = (cuifregS_4 & ((\Mux15~9_combout ))) # (!cuifregS_4 & (\Mux15~19_combout ))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux15~19_combout ),
	.datad(\Mux15~9_combout ),
	.cin(gnd),
	.combout(Mux15),
	.cout());
// synopsys translate_off
defparam \Mux15~20 .lut_mask = 16'hFC30;
defparam \Mux15~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N30
cycloneive_lcell_comb \Mux16~20 (
// Equation(s):
// Mux16 = (cuifregS_4 & (\Mux16~9_combout )) # (!cuifregS_4 & ((\Mux16~19_combout )))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux16~9_combout ),
	.datad(\Mux16~19_combout ),
	.cin(gnd),
	.combout(Mux16),
	.cout());
// synopsys translate_off
defparam \Mux16~20 .lut_mask = 16'hF3C0;
defparam \Mux16~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N22
cycloneive_lcell_comb \Mux17~20 (
// Equation(s):
// Mux17 = (cuifregS_4 & ((\Mux17~9_combout ))) # (!cuifregS_4 & (\Mux17~19_combout ))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux17~19_combout ),
	.datad(\Mux17~9_combout ),
	.cin(gnd),
	.combout(Mux17),
	.cout());
// synopsys translate_off
defparam \Mux17~20 .lut_mask = 16'hFC30;
defparam \Mux17~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N30
cycloneive_lcell_comb \Mux18~20 (
// Equation(s):
// Mux18 = (cuifregS_4 & (\Mux18~9_combout )) # (!cuifregS_4 & ((\Mux18~19_combout )))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux18~9_combout ),
	.datad(\Mux18~19_combout ),
	.cin(gnd),
	.combout(Mux18),
	.cout());
// synopsys translate_off
defparam \Mux18~20 .lut_mask = 16'hF3C0;
defparam \Mux18~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N22
cycloneive_lcell_comb \Mux19~20 (
// Equation(s):
// Mux19 = (cuifregS_4 & (\Mux19~9_combout )) # (!cuifregS_4 & ((\Mux19~19_combout )))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux19~9_combout ),
	.datad(\Mux19~19_combout ),
	.cin(gnd),
	.combout(Mux19),
	.cout());
// synopsys translate_off
defparam \Mux19~20 .lut_mask = 16'hF3C0;
defparam \Mux19~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N30
cycloneive_lcell_comb \Mux20~20 (
// Equation(s):
// Mux20 = (cuifregS_4 & (\Mux20~9_combout )) # (!cuifregS_4 & ((\Mux20~19_combout )))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux20~9_combout ),
	.datad(\Mux20~19_combout ),
	.cin(gnd),
	.combout(Mux20),
	.cout());
// synopsys translate_off
defparam \Mux20~20 .lut_mask = 16'hF3C0;
defparam \Mux20~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N26
cycloneive_lcell_comb \Mux21~20 (
// Equation(s):
// Mux21 = (cuifregS_4 & (\Mux21~9_combout )) # (!cuifregS_4 & ((\Mux21~19_combout )))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux21~9_combout ),
	.datad(\Mux21~19_combout ),
	.cin(gnd),
	.combout(Mux21),
	.cout());
// synopsys translate_off
defparam \Mux21~20 .lut_mask = 16'hF3C0;
defparam \Mux21~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N10
cycloneive_lcell_comb \Mux22~20 (
// Equation(s):
// Mux22 = (cuifregS_4 & (\Mux22~9_combout )) # (!cuifregS_4 & ((\Mux22~19_combout )))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux22~9_combout ),
	.datad(\Mux22~19_combout ),
	.cin(gnd),
	.combout(Mux22),
	.cout());
// synopsys translate_off
defparam \Mux22~20 .lut_mask = 16'hF3C0;
defparam \Mux22~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N10
cycloneive_lcell_comb \Mux59~9 (
// Equation(s):
// Mux59 = (cuifregT_01 & ((\Mux59~6_combout  & ((\Mux59~8_combout ))) # (!\Mux59~6_combout  & (\Mux59~1_combout )))) # (!cuifregT_01 & (\Mux59~6_combout ))

	.dataa(cuifregT_0),
	.datab(\Mux59~6_combout ),
	.datac(\Mux59~1_combout ),
	.datad(\Mux59~8_combout ),
	.cin(gnd),
	.combout(Mux59),
	.cout());
// synopsys translate_off
defparam \Mux59~9 .lut_mask = 16'hEC64;
defparam \Mux59~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N24
cycloneive_lcell_comb \Mux59~19 (
// Equation(s):
// Mux591 = (cuifregT_3 & ((\Mux59~16_combout  & ((\Mux59~18_combout ))) # (!\Mux59~16_combout  & (\Mux59~11_combout )))) # (!cuifregT_3 & (((\Mux59~16_combout ))))

	.dataa(\Mux59~11_combout ),
	.datab(cuifregT_3),
	.datac(\Mux59~18_combout ),
	.datad(\Mux59~16_combout ),
	.cin(gnd),
	.combout(Mux591),
	.cout());
// synopsys translate_off
defparam \Mux59~19 .lut_mask = 16'hF388;
defparam \Mux59~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N6
cycloneive_lcell_comb \Mux0~20 (
// Equation(s):
// Mux0 = (cuifregS_4 & ((\Mux0~9_combout ))) # (!cuifregS_4 & (\Mux0~19_combout ))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux0~19_combout ),
	.datad(\Mux0~9_combout ),
	.cin(gnd),
	.combout(Mux0),
	.cout());
// synopsys translate_off
defparam \Mux0~20 .lut_mask = 16'hFC30;
defparam \Mux0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N12
cycloneive_lcell_comb \Mux2~20 (
// Equation(s):
// Mux2 = (cuifregS_4 & (\Mux2~9_combout )) # (!cuifregS_4 & ((\Mux2~19_combout )))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux2~9_combout ),
	.datad(\Mux2~19_combout ),
	.cin(gnd),
	.combout(Mux2),
	.cout());
// synopsys translate_off
defparam \Mux2~20 .lut_mask = 16'hF3C0;
defparam \Mux2~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N12
cycloneive_lcell_comb \Mux1~20 (
// Equation(s):
// Mux1 = (cuifregS_4 & ((\Mux1~9_combout ))) # (!cuifregS_4 & (\Mux1~19_combout ))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux1~19_combout ),
	.datad(\Mux1~9_combout ),
	.cin(gnd),
	.combout(Mux1),
	.cout());
// synopsys translate_off
defparam \Mux1~20 .lut_mask = 16'hFC30;
defparam \Mux1~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N10
cycloneive_lcell_comb \Mux3~20 (
// Equation(s):
// Mux3 = (cuifregS_4 & (\Mux3~9_combout )) # (!cuifregS_4 & ((\Mux3~19_combout )))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux3~9_combout ),
	.datad(\Mux3~19_combout ),
	.cin(gnd),
	.combout(Mux3),
	.cout());
// synopsys translate_off
defparam \Mux3~20 .lut_mask = 16'hF3C0;
defparam \Mux3~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N0
cycloneive_lcell_comb \Mux4~20 (
// Equation(s):
// Mux4 = (cuifregS_4 & (\Mux4~9_combout )) # (!cuifregS_4 & ((\Mux4~19_combout )))

	.dataa(\Mux4~9_combout ),
	.datab(gnd),
	.datac(cuifregS_4),
	.datad(\Mux4~19_combout ),
	.cin(gnd),
	.combout(Mux4),
	.cout());
// synopsys translate_off
defparam \Mux4~20 .lut_mask = 16'hAFA0;
defparam \Mux4~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N30
cycloneive_lcell_comb \Mux5~20 (
// Equation(s):
// Mux5 = (cuifregS_4 & ((\Mux5~9_combout ))) # (!cuifregS_4 & (\Mux5~19_combout ))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux5~19_combout ),
	.datad(\Mux5~9_combout ),
	.cin(gnd),
	.combout(Mux5),
	.cout());
// synopsys translate_off
defparam \Mux5~20 .lut_mask = 16'hFC30;
defparam \Mux5~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N14
cycloneive_lcell_comb \Mux6~20 (
// Equation(s):
// Mux6 = (cuifregS_4 & (\Mux6~9_combout )) # (!cuifregS_4 & ((\Mux6~19_combout )))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux6~9_combout ),
	.datad(\Mux6~19_combout ),
	.cin(gnd),
	.combout(Mux6),
	.cout());
// synopsys translate_off
defparam \Mux6~20 .lut_mask = 16'hF3C0;
defparam \Mux6~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N2
cycloneive_lcell_comb \Mux7~20 (
// Equation(s):
// Mux7 = (cuifregS_4 & (\Mux7~9_combout )) # (!cuifregS_4 & ((\Mux7~19_combout )))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux7~9_combout ),
	.datad(\Mux7~19_combout ),
	.cin(gnd),
	.combout(Mux7),
	.cout());
// synopsys translate_off
defparam \Mux7~20 .lut_mask = 16'hF3C0;
defparam \Mux7~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N26
cycloneive_lcell_comb \Mux8~20 (
// Equation(s):
// Mux8 = (cuifregS_4 & (\Mux8~9_combout )) # (!cuifregS_4 & ((\Mux8~19_combout )))

	.dataa(cuifregS_4),
	.datab(gnd),
	.datac(\Mux8~9_combout ),
	.datad(\Mux8~19_combout ),
	.cin(gnd),
	.combout(Mux8),
	.cout());
// synopsys translate_off
defparam \Mux8~20 .lut_mask = 16'hF5A0;
defparam \Mux8~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N6
cycloneive_lcell_comb \Mux9~20 (
// Equation(s):
// Mux9 = (cuifregS_4 & ((\Mux9~9_combout ))) # (!cuifregS_4 & (\Mux9~19_combout ))

	.dataa(cuifregS_4),
	.datab(gnd),
	.datac(\Mux9~19_combout ),
	.datad(\Mux9~9_combout ),
	.cin(gnd),
	.combout(Mux9),
	.cout());
// synopsys translate_off
defparam \Mux9~20 .lut_mask = 16'hFA50;
defparam \Mux9~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N0
cycloneive_lcell_comb \Mux10~20 (
// Equation(s):
// Mux10 = (cuifregS_4 & ((\Mux10~9_combout ))) # (!cuifregS_4 & (\Mux10~19_combout ))

	.dataa(cuifregS_4),
	.datab(gnd),
	.datac(\Mux10~19_combout ),
	.datad(\Mux10~9_combout ),
	.cin(gnd),
	.combout(Mux10),
	.cout());
// synopsys translate_off
defparam \Mux10~20 .lut_mask = 16'hFA50;
defparam \Mux10~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N28
cycloneive_lcell_comb \Mux11~20 (
// Equation(s):
// Mux11 = (cuifregS_4 & ((\Mux11~9_combout ))) # (!cuifregS_4 & (\Mux11~19_combout ))

	.dataa(cuifregS_4),
	.datab(\Mux11~19_combout ),
	.datac(gnd),
	.datad(\Mux11~9_combout ),
	.cin(gnd),
	.combout(Mux11),
	.cout());
// synopsys translate_off
defparam \Mux11~20 .lut_mask = 16'hEE44;
defparam \Mux11~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N6
cycloneive_lcell_comb \Mux12~20 (
// Equation(s):
// Mux12 = (cuifregS_4 & (\Mux12~9_combout )) # (!cuifregS_4 & ((\Mux12~19_combout )))

	.dataa(cuifregS_4),
	.datab(gnd),
	.datac(\Mux12~9_combout ),
	.datad(\Mux12~19_combout ),
	.cin(gnd),
	.combout(Mux12),
	.cout());
// synopsys translate_off
defparam \Mux12~20 .lut_mask = 16'hF5A0;
defparam \Mux12~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N14
cycloneive_lcell_comb \Mux13~20 (
// Equation(s):
// Mux13 = (cuifregS_4 & (\Mux13~9_combout )) # (!cuifregS_4 & ((\Mux13~19_combout )))

	.dataa(gnd),
	.datab(\Mux13~9_combout ),
	.datac(cuifregS_4),
	.datad(\Mux13~19_combout ),
	.cin(gnd),
	.combout(Mux13),
	.cout());
// synopsys translate_off
defparam \Mux13~20 .lut_mask = 16'hCFC0;
defparam \Mux13~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N26
cycloneive_lcell_comb \Mux14~20 (
// Equation(s):
// Mux14 = (cuifregS_4 & ((\Mux14~9_combout ))) # (!cuifregS_4 & (\Mux14~19_combout ))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux14~19_combout ),
	.datad(\Mux14~9_combout ),
	.cin(gnd),
	.combout(Mux14),
	.cout());
// synopsys translate_off
defparam \Mux14~20 .lut_mask = 16'hFC30;
defparam \Mux14~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N18
cycloneive_lcell_comb \Mux31~20 (
// Equation(s):
// Mux31 = (cuifregS_4 & ((\Mux31~9_combout ))) # (!cuifregS_4 & (\Mux31~19_combout ))

	.dataa(gnd),
	.datab(cuifregS_4),
	.datac(\Mux31~19_combout ),
	.datad(\Mux31~9_combout ),
	.cin(gnd),
	.combout(Mux31),
	.cout());
// synopsys translate_off
defparam \Mux31~20 .lut_mask = 16'hFC30;
defparam \Mux31~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N4
cycloneive_lcell_comb \Decoder0~50 (
// Equation(s):
// \Decoder0~50_combout  = (\Mux1~1_combout  & (\Mux0~2_combout  & (\WEN~5_combout  & always1)))

	.dataa(Mux110),
	.datab(Mux01),
	.datac(WEN),
	.datad(always1),
	.cin(gnd),
	.combout(\Decoder0~50_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~50 .lut_mask = 16'h8000;
defparam \Decoder0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N28
cycloneive_lcell_comb \Decoder0~68 (
// Equation(s):
// \Decoder0~68_combout  = (\Mux3~1_combout  & (\Decoder0~50_combout  & (\Mux4~1_combout  & !\Mux2~1_combout )))

	.dataa(Mux310),
	.datab(\Decoder0~50_combout ),
	.datac(Mux410),
	.datad(Mux210),
	.cin(gnd),
	.combout(\Decoder0~68_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~68 .lut_mask = 16'h0080;
defparam \Decoder0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N21
dffeas \registerArray[27][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][0] .is_wysiwyg = "true";
defparam \registerArray[27][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N10
cycloneive_lcell_comb \Decoder0~71 (
// Equation(s):
// \Decoder0~71_combout  = (\Mux2~1_combout  & (\Mux3~1_combout  & (\Decoder0~50_combout  & \Mux4~1_combout )))

	.dataa(Mux210),
	.datab(Mux310),
	.datac(\Decoder0~50_combout ),
	.datad(Mux410),
	.cin(gnd),
	.combout(\Decoder0~71_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~71 .lut_mask = 16'h8000;
defparam \Decoder0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N27
dffeas \registerArray[31][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][0] .is_wysiwyg = "true";
defparam \registerArray[31][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N10
cycloneive_lcell_comb \Decoder0~54 (
// Equation(s):
// \Decoder0~54_combout  = (!\Mux1~1_combout  & (\Mux3~1_combout  & (\WEN~5_combout  & always1)))

	.dataa(Mux110),
	.datab(Mux310),
	.datac(WEN),
	.datad(always1),
	.cin(gnd),
	.combout(\Decoder0~54_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~54 .lut_mask = 16'h4000;
defparam \Decoder0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N24
cycloneive_lcell_comb \Decoder0~70 (
// Equation(s):
// \Decoder0~70_combout  = (\Mux4~1_combout  & (!\Mux2~1_combout  & (\Mux0~2_combout  & \Decoder0~54_combout )))

	.dataa(Mux410),
	.datab(Mux210),
	.datac(Mux01),
	.datad(\Decoder0~54_combout ),
	.cin(gnd),
	.combout(\Decoder0~70_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~70 .lut_mask = 16'h2000;
defparam \Decoder0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N17
dffeas \registerArray[19][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][0] .is_wysiwyg = "true";
defparam \registerArray[19][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N16
cycloneive_lcell_comb \Mux63~7 (
// Equation(s):
// \Mux63~7_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[23][0]~q )) # (!cuifregT_2 & ((\registerArray[19][0]~q )))))

	.dataa(\registerArray[23][0]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[19][0]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux63~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~7 .lut_mask = 16'hEE30;
defparam \Mux63~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N26
cycloneive_lcell_comb \Mux63~8 (
// Equation(s):
// \Mux63~8_combout  = (cuifregT_3 & ((\Mux63~7_combout  & ((\registerArray[31][0]~q ))) # (!\Mux63~7_combout  & (\registerArray[27][0]~q )))) # (!cuifregT_3 & (((\Mux63~7_combout ))))

	.dataa(\registerArray[27][0]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[31][0]~q ),
	.datad(\Mux63~7_combout ),
	.cin(gnd),
	.combout(\Mux63~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~8 .lut_mask = 16'hF388;
defparam \Mux63~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N12
cycloneive_lcell_comb \registerArray[25][0]~feeder (
// Equation(s):
// \registerArray[25][0]~feeder_combout  = \Mux68~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux68),
	.cin(gnd),
	.combout(\registerArray[25][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[25][0]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[25][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N2
cycloneive_lcell_comb \Decoder0~60 (
// Equation(s):
// \Decoder0~60_combout  = (!\Mux3~1_combout  & (\Decoder0~50_combout  & (\Mux4~1_combout  & !\Mux2~1_combout )))

	.dataa(Mux310),
	.datab(\Decoder0~50_combout ),
	.datac(Mux410),
	.datad(Mux210),
	.cin(gnd),
	.combout(\Decoder0~60_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~60 .lut_mask = 16'h0040;
defparam \Decoder0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y40_N13
dffeas \registerArray[25][0] (
	.clk(clk),
	.d(\registerArray[25][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][0] .is_wysiwyg = "true";
defparam \registerArray[25][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N16
cycloneive_lcell_comb \Decoder0~61 (
// Equation(s):
// \Decoder0~61_combout  = (!\Mux3~1_combout  & (\Decoder0~50_combout  & (\Mux4~1_combout  & \Mux2~1_combout )))

	.dataa(Mux310),
	.datab(\Decoder0~50_combout ),
	.datac(Mux410),
	.datad(Mux210),
	.cin(gnd),
	.combout(\Decoder0~61_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~61 .lut_mask = 16'h4000;
defparam \Decoder0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N19
dffeas \registerArray[29][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][0] .is_wysiwyg = "true";
defparam \registerArray[29][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N28
cycloneive_lcell_comb \Decoder0~51 (
// Equation(s):
// \Decoder0~51_combout  = (\WEN~5_combout  & (!\Mux3~1_combout  & (!\Mux1~1_combout  & always1)))

	.dataa(WEN),
	.datab(Mux310),
	.datac(Mux110),
	.datad(always1),
	.cin(gnd),
	.combout(\Decoder0~51_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~51 .lut_mask = 16'h0200;
defparam \Decoder0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N0
cycloneive_lcell_comb \Decoder0~53 (
// Equation(s):
// \Decoder0~53_combout  = (\Mux4~1_combout  & (!\Mux2~1_combout  & (\Mux0~2_combout  & \Decoder0~51_combout )))

	.dataa(Mux410),
	.datab(Mux210),
	.datac(Mux01),
	.datad(\Decoder0~51_combout ),
	.cin(gnd),
	.combout(\Decoder0~53_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~53 .lut_mask = 16'h2000;
defparam \Decoder0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N13
dffeas \registerArray[17][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][0] .is_wysiwyg = "true";
defparam \registerArray[17][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N12
cycloneive_lcell_comb \Mux63~0 (
// Equation(s):
// \Mux63~0_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[21][0]~q )) # (!cuifregT_2 & ((\registerArray[17][0]~q )))))

	.dataa(\registerArray[21][0]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[17][0]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux63~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~0 .lut_mask = 16'hEE30;
defparam \Mux63~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N18
cycloneive_lcell_comb \Mux63~1 (
// Equation(s):
// \Mux63~1_combout  = (cuifregT_3 & ((\Mux63~0_combout  & ((\registerArray[29][0]~q ))) # (!\Mux63~0_combout  & (\registerArray[25][0]~q )))) # (!cuifregT_3 & (((\Mux63~0_combout ))))

	.dataa(\registerArray[25][0]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[29][0]~q ),
	.datad(\Mux63~0_combout ),
	.cin(gnd),
	.combout(\Mux63~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~1 .lut_mask = 16'hF388;
defparam \Mux63~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N8
cycloneive_lcell_comb \registerArray[22][0]~feeder (
// Equation(s):
// \registerArray[22][0]~feeder_combout  = \Mux68~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux68),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[22][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[22][0]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[22][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N22
cycloneive_lcell_comb \Decoder0~62 (
// Equation(s):
// \Decoder0~62_combout  = (\Mux2~1_combout  & (\Decoder0~54_combout  & (\Mux0~2_combout  & !\Mux4~1_combout )))

	.dataa(Mux210),
	.datab(\Decoder0~54_combout ),
	.datac(Mux01),
	.datad(Mux410),
	.cin(gnd),
	.combout(\Decoder0~62_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~62 .lut_mask = 16'h0080;
defparam \Decoder0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N9
dffeas \registerArray[22][0] (
	.clk(clk),
	.d(\registerArray[22][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][0] .is_wysiwyg = "true";
defparam \registerArray[22][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N24
cycloneive_lcell_comb \Decoder0~65 (
// Equation(s):
// \Decoder0~65_combout  = (!\Mux4~1_combout  & (\Mux2~1_combout  & (\Mux3~1_combout  & \Decoder0~50_combout )))

	.dataa(Mux410),
	.datab(Mux210),
	.datac(Mux310),
	.datad(\Decoder0~50_combout ),
	.cin(gnd),
	.combout(\Decoder0~65_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~65 .lut_mask = 16'h4000;
defparam \Decoder0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N15
dffeas \registerArray[30][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][0] .is_wysiwyg = "true";
defparam \registerArray[30][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N18
cycloneive_lcell_comb \Decoder0~64 (
// Equation(s):
// \Decoder0~64_combout  = (!\Mux4~1_combout  & (!\Mux2~1_combout  & (\Mux0~2_combout  & \Decoder0~54_combout )))

	.dataa(Mux410),
	.datab(Mux210),
	.datac(Mux01),
	.datad(\Decoder0~54_combout ),
	.cin(gnd),
	.combout(\Decoder0~64_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~64 .lut_mask = 16'h1000;
defparam \Decoder0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N1
dffeas \registerArray[18][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][0] .is_wysiwyg = "true";
defparam \registerArray[18][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N0
cycloneive_lcell_comb \Mux63~2 (
// Equation(s):
// \Mux63~2_combout  = (cuifregT_3 & ((\registerArray[26][0]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[18][0]~q  & !cuifregT_2))))

	.dataa(\registerArray[26][0]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[18][0]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux63~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~2 .lut_mask = 16'hCCB8;
defparam \Mux63~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N14
cycloneive_lcell_comb \Mux63~3 (
// Equation(s):
// \Mux63~3_combout  = (cuifregT_2 & ((\Mux63~2_combout  & ((\registerArray[30][0]~q ))) # (!\Mux63~2_combout  & (\registerArray[22][0]~q )))) # (!cuifregT_2 & (((\Mux63~2_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[22][0]~q ),
	.datac(\registerArray[30][0]~q ),
	.datad(\Mux63~2_combout ),
	.cin(gnd),
	.combout(\Mux63~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~3 .lut_mask = 16'hF588;
defparam \Mux63~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N8
cycloneive_lcell_comb \Decoder0~67 (
// Equation(s):
// \Decoder0~67_combout  = (\Mux2~1_combout  & (!\Mux3~1_combout  & (\Decoder0~50_combout  & !\Mux4~1_combout )))

	.dataa(Mux210),
	.datab(Mux310),
	.datac(\Decoder0~50_combout ),
	.datad(Mux410),
	.cin(gnd),
	.combout(\Decoder0~67_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~67 .lut_mask = 16'h0020;
defparam \Decoder0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N3
dffeas \registerArray[28][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][0] .is_wysiwyg = "true";
defparam \registerArray[28][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N30
cycloneive_lcell_comb \registerArray[24][0]~feeder (
// Equation(s):
// \registerArray[24][0]~feeder_combout  = \Mux68~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux68),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[24][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[24][0]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[24][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N30
cycloneive_lcell_comb \Decoder0~66 (
// Equation(s):
// \Decoder0~66_combout  = (!\Mux3~1_combout  & (\Decoder0~50_combout  & (!\Mux4~1_combout  & !\Mux2~1_combout )))

	.dataa(Mux310),
	.datab(\Decoder0~50_combout ),
	.datac(Mux410),
	.datad(Mux210),
	.cin(gnd),
	.combout(\Decoder0~66_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~66 .lut_mask = 16'h0004;
defparam \Decoder0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N31
dffeas \registerArray[24][0] (
	.clk(clk),
	.d(\registerArray[24][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][0] .is_wysiwyg = "true";
defparam \registerArray[24][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N12
cycloneive_lcell_comb \Decoder0~56 (
// Equation(s):
// \Decoder0~56_combout  = (\Decoder0~51_combout  & (\Mux0~2_combout  & (!\Mux4~1_combout  & !\Mux2~1_combout )))

	.dataa(\Decoder0~51_combout ),
	.datab(Mux01),
	.datac(Mux410),
	.datad(Mux210),
	.cin(gnd),
	.combout(\Decoder0~56_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~56 .lut_mask = 16'h0008;
defparam \Decoder0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N21
dffeas \registerArray[16][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][0] .is_wysiwyg = "true";
defparam \registerArray[16][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N20
cycloneive_lcell_comb \Mux63~4 (
// Equation(s):
// \Mux63~4_combout  = (cuifregT_3 & ((\registerArray[24][0]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[16][0]~q  & !cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[24][0]~q ),
	.datac(\registerArray[16][0]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux63~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~4 .lut_mask = 16'hAAD8;
defparam \Mux63~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N2
cycloneive_lcell_comb \Mux63~5 (
// Equation(s):
// \Mux63~5_combout  = (cuifregT_2 & ((\Mux63~4_combout  & ((\registerArray[28][0]~q ))) # (!\Mux63~4_combout  & (\registerArray[20][0]~q )))) # (!cuifregT_2 & (((\Mux63~4_combout ))))

	.dataa(\registerArray[20][0]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[28][0]~q ),
	.datad(\Mux63~4_combout ),
	.cin(gnd),
	.combout(\Mux63~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~5 .lut_mask = 16'hF388;
defparam \Mux63~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N12
cycloneive_lcell_comb \Mux63~6 (
// Equation(s):
// \Mux63~6_combout  = (cuifregT_01 & (cuifregT_1)) # (!cuifregT_01 & ((cuifregT_1 & (\Mux63~3_combout )) # (!cuifregT_1 & ((\Mux63~5_combout )))))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\Mux63~3_combout ),
	.datad(\Mux63~5_combout ),
	.cin(gnd),
	.combout(\Mux63~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~6 .lut_mask = 16'hD9C8;
defparam \Mux63~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N2
cycloneive_lcell_comb \Decoder0~57 (
// Equation(s):
// \Decoder0~57_combout  = (\Mux1~1_combout  & (!\Mux0~2_combout  & (\WEN~5_combout  & always1)))

	.dataa(Mux110),
	.datab(Mux01),
	.datac(WEN),
	.datad(always1),
	.cin(gnd),
	.combout(\Decoder0~57_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~57 .lut_mask = 16'h2000;
defparam \Decoder0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N20
cycloneive_lcell_comb \Decoder0~75 (
// Equation(s):
// \Decoder0~75_combout  = (\Mux3~1_combout  & (\Decoder0~57_combout  & (\Mux4~1_combout  & !\Mux2~1_combout )))

	.dataa(Mux310),
	.datab(\Decoder0~57_combout ),
	.datac(Mux410),
	.datad(Mux210),
	.cin(gnd),
	.combout(\Decoder0~75_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~75 .lut_mask = 16'h0080;
defparam \Decoder0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N23
dffeas \registerArray[11][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][0] .is_wysiwyg = "true";
defparam \registerArray[11][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N14
cycloneive_lcell_comb \Decoder0~72 (
// Equation(s):
// \Decoder0~72_combout  = (\Mux4~1_combout  & (!\Mux3~1_combout  & (!\Mux2~1_combout  & \Decoder0~57_combout )))

	.dataa(Mux410),
	.datab(Mux310),
	.datac(Mux210),
	.datad(\Decoder0~57_combout ),
	.cin(gnd),
	.combout(\Decoder0~72_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~72 .lut_mask = 16'h0200;
defparam \Decoder0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N21
dffeas \registerArray[9][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][0] .is_wysiwyg = "true";
defparam \registerArray[9][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N8
cycloneive_lcell_comb \registerArray[10][0]~feeder (
// Equation(s):
// \registerArray[10][0]~feeder_combout  = \Mux68~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux68),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[10][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[10][0]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[10][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N2
cycloneive_lcell_comb \Decoder0~73 (
// Equation(s):
// \Decoder0~73_combout  = (\Mux3~1_combout  & (!\Mux4~1_combout  & (\Decoder0~57_combout  & !\Mux2~1_combout )))

	.dataa(Mux310),
	.datab(Mux410),
	.datac(\Decoder0~57_combout ),
	.datad(Mux210),
	.cin(gnd),
	.combout(\Decoder0~73_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~73 .lut_mask = 16'h0020;
defparam \Decoder0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N9
dffeas \registerArray[10][0] (
	.clk(clk),
	.d(\registerArray[10][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][0] .is_wysiwyg = "true";
defparam \registerArray[10][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N28
cycloneive_lcell_comb \Mux63~10 (
// Equation(s):
// \Mux63~10_combout  = (cuifregT_1 & (((\registerArray[10][0]~q ) # (cuifregT_01)))) # (!cuifregT_1 & (\registerArray[8][0]~q  & ((!cuifregT_01))))

	.dataa(\registerArray[8][0]~q ),
	.datab(\registerArray[10][0]~q ),
	.datac(cuifregT_1),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux63~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~10 .lut_mask = 16'hF0CA;
defparam \Mux63~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N20
cycloneive_lcell_comb \Mux63~11 (
// Equation(s):
// \Mux63~11_combout  = (cuifregT_01 & ((\Mux63~10_combout  & (\registerArray[11][0]~q )) # (!\Mux63~10_combout  & ((\registerArray[9][0]~q ))))) # (!cuifregT_01 & (((\Mux63~10_combout ))))

	.dataa(cuifregT_0),
	.datab(\registerArray[11][0]~q ),
	.datac(\registerArray[9][0]~q ),
	.datad(\Mux63~10_combout ),
	.cin(gnd),
	.combout(\Mux63~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~11 .lut_mask = 16'hDDA0;
defparam \Mux63~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N8
cycloneive_lcell_comb \registerArray[3][0]~feeder (
// Equation(s):
// \registerArray[3][0]~feeder_combout  = \Mux68~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux68),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[3][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[3][0]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[3][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N24
cycloneive_lcell_comb \Decoder0~78 (
// Equation(s):
// \Decoder0~78_combout  = (\Decoder0~54_combout  & (!\Mux0~2_combout  & (\Mux4~1_combout  & !\Mux2~1_combout )))

	.dataa(\Decoder0~54_combout ),
	.datab(Mux01),
	.datac(Mux410),
	.datad(Mux210),
	.cin(gnd),
	.combout(\Decoder0~78_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~78 .lut_mask = 16'h0020;
defparam \Decoder0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N9
dffeas \registerArray[3][0] (
	.clk(clk),
	.d(\registerArray[3][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][0] .is_wysiwyg = "true";
defparam \registerArray[3][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N26
cycloneive_lcell_comb \Decoder0~79 (
// Equation(s):
// \Decoder0~79_combout  = (\Decoder0~51_combout  & (!\Mux0~2_combout  & (\Mux4~1_combout  & !\Mux2~1_combout )))

	.dataa(\Decoder0~51_combout ),
	.datab(Mux01),
	.datac(Mux410),
	.datad(Mux210),
	.cin(gnd),
	.combout(\Decoder0~79_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~79 .lut_mask = 16'h0020;
defparam \Decoder0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N17
dffeas \registerArray[1][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][0] .is_wysiwyg = "true";
defparam \registerArray[1][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N16
cycloneive_lcell_comb \Mux63~14 (
// Equation(s):
// \Mux63~14_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][0]~q )) # (!cuifregT_1 & ((\registerArray[1][0]~q )))))

	.dataa(cuifregT_0),
	.datab(\registerArray[3][0]~q ),
	.datac(\registerArray[1][0]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux63~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~14 .lut_mask = 16'h88A0;
defparam \Mux63~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N22
cycloneive_lcell_comb \Decoder0~80 (
// Equation(s):
// \Decoder0~80_combout  = (!\Mux4~1_combout  & (!\Mux0~2_combout  & (!\Mux2~1_combout  & \Decoder0~54_combout )))

	.dataa(Mux410),
	.datab(Mux01),
	.datac(Mux210),
	.datad(\Decoder0~54_combout ),
	.cin(gnd),
	.combout(\Decoder0~80_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~80 .lut_mask = 16'h0100;
defparam \Decoder0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N27
dffeas \registerArray[2][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][0] .is_wysiwyg = "true";
defparam \registerArray[2][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N26
cycloneive_lcell_comb \Mux63~15 (
// Equation(s):
// \Mux63~15_combout  = (\Mux63~14_combout ) # ((!cuifregT_01 & (\registerArray[2][0]~q  & cuifregT_1)))

	.dataa(cuifregT_0),
	.datab(\Mux63~14_combout ),
	.datac(\registerArray[2][0]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux63~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~15 .lut_mask = 16'hDCCC;
defparam \Mux63~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N8
cycloneive_lcell_comb \Decoder0~77 (
// Equation(s):
// \Decoder0~77_combout  = (\Mux2~1_combout  & (\Decoder0~54_combout  & (!\Mux0~2_combout  & \Mux4~1_combout )))

	.dataa(Mux210),
	.datab(\Decoder0~54_combout ),
	.datac(Mux01),
	.datad(Mux410),
	.cin(gnd),
	.combout(\Decoder0~77_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~77 .lut_mask = 16'h0800;
defparam \Decoder0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N13
dffeas \registerArray[7][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][0] .is_wysiwyg = "true";
defparam \registerArray[7][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N28
cycloneive_lcell_comb \Decoder0~59 (
// Equation(s):
// \Decoder0~59_combout  = (!\Mux4~1_combout  & (!\Mux0~2_combout  & (\Mux2~1_combout  & \Decoder0~51_combout )))

	.dataa(Mux410),
	.datab(Mux01),
	.datac(Mux210),
	.datad(\Decoder0~51_combout ),
	.cin(gnd),
	.combout(\Decoder0~59_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~59 .lut_mask = 16'h1000;
defparam \Decoder0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N27
dffeas \registerArray[4][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][0] .is_wysiwyg = "true";
defparam \registerArray[4][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N26
cycloneive_lcell_comb \Mux63~12 (
// Equation(s):
// \Mux63~12_combout  = (cuifregT_01 & ((\registerArray[5][0]~q ) # ((cuifregT_1)))) # (!cuifregT_01 & (((\registerArray[4][0]~q  & !cuifregT_1))))

	.dataa(\registerArray[5][0]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[4][0]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux63~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~12 .lut_mask = 16'hCCB8;
defparam \Mux63~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N12
cycloneive_lcell_comb \Mux63~13 (
// Equation(s):
// \Mux63~13_combout  = (cuifregT_1 & ((\Mux63~12_combout  & ((\registerArray[7][0]~q ))) # (!\Mux63~12_combout  & (\registerArray[6][0]~q )))) # (!cuifregT_1 & (((\Mux63~12_combout ))))

	.dataa(\registerArray[6][0]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[7][0]~q ),
	.datad(\Mux63~12_combout ),
	.cin(gnd),
	.combout(\Mux63~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~13 .lut_mask = 16'hF388;
defparam \Mux63~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N8
cycloneive_lcell_comb \Mux63~16 (
// Equation(s):
// \Mux63~16_combout  = (cuifregT_3 & (cuifregT_2)) # (!cuifregT_3 & ((cuifregT_2 & ((\Mux63~13_combout ))) # (!cuifregT_2 & (\Mux63~15_combout ))))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\Mux63~15_combout ),
	.datad(\Mux63~13_combout ),
	.cin(gnd),
	.combout(\Mux63~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~16 .lut_mask = 16'hDC98;
defparam \Mux63~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N22
cycloneive_lcell_comb \registerArray[14][0]~feeder (
// Equation(s):
// \registerArray[14][0]~feeder_combout  = \Mux68~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux68),
	.cin(gnd),
	.combout(\registerArray[14][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][0]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[14][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N18
cycloneive_lcell_comb \Decoder0~81 (
// Equation(s):
// \Decoder0~81_combout  = (\Mux3~1_combout  & (\Decoder0~57_combout  & (!\Mux4~1_combout  & \Mux2~1_combout )))

	.dataa(Mux310),
	.datab(\Decoder0~57_combout ),
	.datac(Mux410),
	.datad(Mux210),
	.cin(gnd),
	.combout(\Decoder0~81_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~81 .lut_mask = 16'h0800;
defparam \Decoder0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N23
dffeas \registerArray[14][0] (
	.clk(clk),
	.d(\registerArray[14][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][0] .is_wysiwyg = "true";
defparam \registerArray[14][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N4
cycloneive_lcell_comb \Decoder0~84 (
// Equation(s):
// \Decoder0~84_combout  = (\Mux4~1_combout  & (\Mux2~1_combout  & (\Mux3~1_combout  & \Decoder0~57_combout )))

	.dataa(Mux410),
	.datab(Mux210),
	.datac(Mux310),
	.datad(\Decoder0~57_combout ),
	.cin(gnd),
	.combout(\Decoder0~84_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~84 .lut_mask = 16'h8000;
defparam \Decoder0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y36_N3
dffeas \registerArray[15][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][0] .is_wysiwyg = "true";
defparam \registerArray[15][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N26
cycloneive_lcell_comb \Decoder0~82 (
// Equation(s):
// \Decoder0~82_combout  = (\Mux4~1_combout  & (!\Mux3~1_combout  & (\Mux2~1_combout  & \Decoder0~57_combout )))

	.dataa(Mux410),
	.datab(Mux310),
	.datac(Mux210),
	.datad(\Decoder0~57_combout ),
	.cin(gnd),
	.combout(\Decoder0~82_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~82 .lut_mask = 16'h2000;
defparam \Decoder0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N29
dffeas \registerArray[13][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][0] .is_wysiwyg = "true";
defparam \registerArray[13][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N26
cycloneive_lcell_comb \Decoder0~83 (
// Equation(s):
// \Decoder0~83_combout  = (!\Mux4~1_combout  & (\Mux2~1_combout  & (!\Mux3~1_combout  & \Decoder0~57_combout )))

	.dataa(Mux410),
	.datab(Mux210),
	.datac(Mux310),
	.datad(\Decoder0~57_combout ),
	.cin(gnd),
	.combout(\Decoder0~83_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~83 .lut_mask = 16'h0400;
defparam \Decoder0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y36_N1
dffeas \registerArray[12][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][0] .is_wysiwyg = "true";
defparam \registerArray[12][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N0
cycloneive_lcell_comb \Mux63~17 (
// Equation(s):
// \Mux63~17_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[13][0]~q )) # (!cuifregT_01 & ((\registerArray[12][0]~q )))))

	.dataa(cuifregT_1),
	.datab(\registerArray[13][0]~q ),
	.datac(\registerArray[12][0]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux63~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~17 .lut_mask = 16'hEE50;
defparam \Mux63~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N2
cycloneive_lcell_comb \Mux63~18 (
// Equation(s):
// \Mux63~18_combout  = (cuifregT_1 & ((\Mux63~17_combout  & ((\registerArray[15][0]~q ))) # (!\Mux63~17_combout  & (\registerArray[14][0]~q )))) # (!cuifregT_1 & (((\Mux63~17_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[14][0]~q ),
	.datac(\registerArray[15][0]~q ),
	.datad(\Mux63~17_combout ),
	.cin(gnd),
	.combout(\Mux63~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~18 .lut_mask = 16'hF588;
defparam \Mux63~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N0
cycloneive_lcell_comb \Decoder0~69 (
// Equation(s):
// \Decoder0~69_combout  = (\Mux2~1_combout  & (\Decoder0~54_combout  & (\Mux0~2_combout  & \Mux4~1_combout )))

	.dataa(Mux210),
	.datab(\Decoder0~54_combout ),
	.datac(Mux01),
	.datad(Mux410),
	.cin(gnd),
	.combout(\Decoder0~69_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~69 .lut_mask = 16'h8000;
defparam \Decoder0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N25
dffeas \registerArray[23][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][31] .is_wysiwyg = "true";
defparam \registerArray[23][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N27
dffeas \registerArray[27][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][31] .is_wysiwyg = "true";
defparam \registerArray[27][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N5
dffeas \registerArray[19][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][31] .is_wysiwyg = "true";
defparam \registerArray[19][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N4
cycloneive_lcell_comb \Mux32~7 (
// Equation(s):
// \Mux32~7_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[27][31]~q )) # (!cuifregT_3 & ((\registerArray[19][31]~q )))))

	.dataa(cuifregT_2),
	.datab(\registerArray[27][31]~q ),
	.datac(\registerArray[19][31]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux32~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~7 .lut_mask = 16'hEE50;
defparam \Mux32~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N31
dffeas \registerArray[31][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][31] .is_wysiwyg = "true";
defparam \registerArray[31][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N30
cycloneive_lcell_comb \Mux32~8 (
// Equation(s):
// \Mux32~8_combout  = (\Mux32~7_combout  & (((\registerArray[31][31]~q ) # (!cuifregT_2)))) # (!\Mux32~7_combout  & (\registerArray[23][31]~q  & ((cuifregT_2))))

	.dataa(\registerArray[23][31]~q ),
	.datab(\Mux32~7_combout ),
	.datac(\registerArray[31][31]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux32~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~8 .lut_mask = 16'hE2CC;
defparam \Mux32~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N8
cycloneive_lcell_comb \registerArray[16][31]~feeder (
// Equation(s):
// \registerArray[16][31]~feeder_combout  = \Mux37~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux372),
	.cin(gnd),
	.combout(\registerArray[16][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[16][31]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[16][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N9
dffeas \registerArray[16][31] (
	.clk(clk),
	.d(\registerArray[16][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][31] .is_wysiwyg = "true";
defparam \registerArray[16][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N22
cycloneive_lcell_comb \Decoder0~55 (
// Equation(s):
// \Decoder0~55_combout  = (!\Mux4~1_combout  & (\Mux2~1_combout  & (\Mux0~2_combout  & \Decoder0~51_combout )))

	.dataa(Mux410),
	.datab(Mux210),
	.datac(Mux01),
	.datad(\Decoder0~51_combout ),
	.cin(gnd),
	.combout(\Decoder0~55_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~55 .lut_mask = 16'h4000;
defparam \Decoder0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N27
dffeas \registerArray[20][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][31] .is_wysiwyg = "true";
defparam \registerArray[20][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N28
cycloneive_lcell_comb \Mux32~4 (
// Equation(s):
// \Mux32~4_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & ((\registerArray[20][31]~q ))) # (!cuifregT_2 & (\registerArray[16][31]~q ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[16][31]~q ),
	.datac(\registerArray[20][31]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux32~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~4 .lut_mask = 16'hFA44;
defparam \Mux32~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y34_N19
dffeas \registerArray[28][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][31] .is_wysiwyg = "true";
defparam \registerArray[28][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N18
cycloneive_lcell_comb \Mux32~5 (
// Equation(s):
// \Mux32~5_combout  = (\Mux32~4_combout  & (((\registerArray[28][31]~q ) # (!cuifregT_3)))) # (!\Mux32~4_combout  & (\registerArray[24][31]~q  & ((cuifregT_3))))

	.dataa(\registerArray[24][31]~q ),
	.datab(\Mux32~4_combout ),
	.datac(\registerArray[28][31]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux32~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~5 .lut_mask = 16'hE2CC;
defparam \Mux32~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N7
dffeas \registerArray[30][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][31] .is_wysiwyg = "true";
defparam \registerArray[30][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N13
dffeas \registerArray[18][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][31] .is_wysiwyg = "true";
defparam \registerArray[18][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N12
cycloneive_lcell_comb \Mux32~2 (
// Equation(s):
// \Mux32~2_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[22][31]~q )) # (!cuifregT_2 & ((\registerArray[18][31]~q )))))

	.dataa(\registerArray[22][31]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[18][31]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux32~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~2 .lut_mask = 16'hEE30;
defparam \Mux32~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N6
cycloneive_lcell_comb \Mux32~3 (
// Equation(s):
// \Mux32~3_combout  = (cuifregT_3 & ((\Mux32~2_combout  & ((\registerArray[30][31]~q ))) # (!\Mux32~2_combout  & (\registerArray[26][31]~q )))) # (!cuifregT_3 & (((\Mux32~2_combout ))))

	.dataa(\registerArray[26][31]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[30][31]~q ),
	.datad(\Mux32~2_combout ),
	.cin(gnd),
	.combout(\Mux32~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~3 .lut_mask = 16'hF388;
defparam \Mux32~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N8
cycloneive_lcell_comb \Mux32~6 (
// Equation(s):
// \Mux32~6_combout  = (cuifregT_1 & (((cuifregT_01) # (\Mux32~3_combout )))) # (!cuifregT_1 & (\Mux32~5_combout  & (!cuifregT_01)))

	.dataa(cuifregT_1),
	.datab(\Mux32~5_combout ),
	.datac(cuifregT_0),
	.datad(\Mux32~3_combout ),
	.cin(gnd),
	.combout(\Mux32~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~6 .lut_mask = 16'hAEA4;
defparam \Mux32~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N16
cycloneive_lcell_comb \registerArray[21][31]~feeder (
// Equation(s):
// \registerArray[21][31]~feeder_combout  = \Mux37~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux372),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[21][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[21][31]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[21][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N18
cycloneive_lcell_comb \Decoder0~52 (
// Equation(s):
// \Decoder0~52_combout  = (\Mux4~1_combout  & (\Mux2~1_combout  & (\Mux0~2_combout  & \Decoder0~51_combout )))

	.dataa(Mux410),
	.datab(Mux210),
	.datac(Mux01),
	.datad(\Decoder0~51_combout ),
	.cin(gnd),
	.combout(\Decoder0~52_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~52 .lut_mask = 16'h8000;
defparam \Decoder0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y44_N17
dffeas \registerArray[21][31] (
	.clk(clk),
	.d(\registerArray[21][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][31] .is_wysiwyg = "true";
defparam \registerArray[21][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N18
cycloneive_lcell_comb \registerArray[25][31]~feeder (
// Equation(s):
// \registerArray[25][31]~feeder_combout  = \Mux37~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux372),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[25][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[25][31]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[25][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N19
dffeas \registerArray[25][31] (
	.clk(clk),
	.d(\registerArray[25][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][31] .is_wysiwyg = "true";
defparam \registerArray[25][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N5
dffeas \registerArray[17][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][31] .is_wysiwyg = "true";
defparam \registerArray[17][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N4
cycloneive_lcell_comb \Mux32~0 (
// Equation(s):
// \Mux32~0_combout  = (cuifregT_3 & ((\registerArray[25][31]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[17][31]~q  & !cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[25][31]~q ),
	.datac(\registerArray[17][31]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux32~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~0 .lut_mask = 16'hAAD8;
defparam \Mux32~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N19
dffeas \registerArray[29][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][31] .is_wysiwyg = "true";
defparam \registerArray[29][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N18
cycloneive_lcell_comb \Mux32~1 (
// Equation(s):
// \Mux32~1_combout  = (\Mux32~0_combout  & (((\registerArray[29][31]~q ) # (!cuifregT_2)))) # (!\Mux32~0_combout  & (\registerArray[21][31]~q  & ((cuifregT_2))))

	.dataa(\registerArray[21][31]~q ),
	.datab(\Mux32~0_combout ),
	.datac(\registerArray[29][31]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux32~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~1 .lut_mask = 16'hE2CC;
defparam \Mux32~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N16
cycloneive_lcell_comb \Decoder0~76 (
// Equation(s):
// \Decoder0~76_combout  = (\Decoder0~54_combout  & (!\Mux0~2_combout  & (!\Mux4~1_combout  & \Mux2~1_combout )))

	.dataa(\Decoder0~54_combout ),
	.datab(Mux01),
	.datac(Mux410),
	.datad(Mux210),
	.cin(gnd),
	.combout(\Decoder0~76_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~76 .lut_mask = 16'h0200;
defparam \Decoder0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N5
dffeas \registerArray[6][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][31] .is_wysiwyg = "true";
defparam \registerArray[6][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N4
cycloneive_lcell_comb \Decoder0~58 (
// Equation(s):
// \Decoder0~58_combout  = (\Mux4~1_combout  & (\Mux2~1_combout  & (!\Mux0~2_combout  & \Decoder0~51_combout )))

	.dataa(Mux410),
	.datab(Mux210),
	.datac(Mux01),
	.datad(\Decoder0~51_combout ),
	.cin(gnd),
	.combout(\Decoder0~58_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~58 .lut_mask = 16'h0800;
defparam \Decoder0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N5
dffeas \registerArray[5][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][31] .is_wysiwyg = "true";
defparam \registerArray[5][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N4
cycloneive_lcell_comb \Mux32~10 (
// Equation(s):
// \Mux32~10_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & ((\registerArray[5][31]~q ))) # (!cuifregT_01 & (\registerArray[4][31]~q ))))

	.dataa(\registerArray[4][31]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[5][31]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux32~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~10 .lut_mask = 16'hFC22;
defparam \Mux32~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N3
dffeas \registerArray[7][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][31] .is_wysiwyg = "true";
defparam \registerArray[7][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N2
cycloneive_lcell_comb \Mux32~11 (
// Equation(s):
// \Mux32~11_combout  = (\Mux32~10_combout  & (((\registerArray[7][31]~q ) # (!cuifregT_1)))) # (!\Mux32~10_combout  & (\registerArray[6][31]~q  & ((cuifregT_1))))

	.dataa(\registerArray[6][31]~q ),
	.datab(\Mux32~10_combout ),
	.datac(\registerArray[7][31]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux32~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~11 .lut_mask = 16'hE2CC;
defparam \Mux32~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N3
dffeas \registerArray[14][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][31] .is_wysiwyg = "true";
defparam \registerArray[14][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N19
dffeas \registerArray[15][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][31] .is_wysiwyg = "true";
defparam \registerArray[15][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N1
dffeas \registerArray[13][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][31] .is_wysiwyg = "true";
defparam \registerArray[13][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N17
dffeas \registerArray[12][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][31] .is_wysiwyg = "true";
defparam \registerArray[12][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N16
cycloneive_lcell_comb \Mux32~17 (
// Equation(s):
// \Mux32~17_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[13][31]~q )) # (!cuifregT_01 & ((\registerArray[12][31]~q )))))

	.dataa(cuifregT_1),
	.datab(\registerArray[13][31]~q ),
	.datac(\registerArray[12][31]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux32~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~17 .lut_mask = 16'hEE50;
defparam \Mux32~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N18
cycloneive_lcell_comb \Mux32~18 (
// Equation(s):
// \Mux32~18_combout  = (cuifregT_1 & ((\Mux32~17_combout  & ((\registerArray[15][31]~q ))) # (!\Mux32~17_combout  & (\registerArray[14][31]~q )))) # (!cuifregT_1 & (((\Mux32~17_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[14][31]~q ),
	.datac(\registerArray[15][31]~q ),
	.datad(\Mux32~17_combout ),
	.cin(gnd),
	.combout(\Mux32~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~18 .lut_mask = 16'hF588;
defparam \Mux32~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N26
cycloneive_lcell_comb \Decoder0~74 (
// Equation(s):
// \Decoder0~74_combout  = (!\Mux3~1_combout  & (\Decoder0~57_combout  & (!\Mux4~1_combout  & !\Mux2~1_combout )))

	.dataa(Mux310),
	.datab(\Decoder0~57_combout ),
	.datac(Mux410),
	.datad(Mux210),
	.cin(gnd),
	.combout(\Decoder0~74_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~74 .lut_mask = 16'h0004;
defparam \Decoder0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N9
dffeas \registerArray[8][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][31] .is_wysiwyg = "true";
defparam \registerArray[8][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N8
cycloneive_lcell_comb \Mux32~12 (
// Equation(s):
// \Mux32~12_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & (\registerArray[10][31]~q )) # (!cuifregT_1 & ((\registerArray[8][31]~q )))))

	.dataa(\registerArray[10][31]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[8][31]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux32~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~12 .lut_mask = 16'hEE30;
defparam \Mux32~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N15
dffeas \registerArray[11][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][31] .is_wysiwyg = "true";
defparam \registerArray[11][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N14
cycloneive_lcell_comb \Mux32~13 (
// Equation(s):
// \Mux32~13_combout  = (\Mux32~12_combout  & (((\registerArray[11][31]~q ) # (!cuifregT_01)))) # (!\Mux32~12_combout  & (\registerArray[9][31]~q  & ((cuifregT_01))))

	.dataa(\registerArray[9][31]~q ),
	.datab(\Mux32~12_combout ),
	.datac(\registerArray[11][31]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux32~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~13 .lut_mask = 16'hE2CC;
defparam \Mux32~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N13
dffeas \registerArray[2][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][31] .is_wysiwyg = "true";
defparam \registerArray[2][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N0
cycloneive_lcell_comb \registerArray[3][31]~feeder (
// Equation(s):
// \registerArray[3][31]~feeder_combout  = \Mux37~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux372),
	.cin(gnd),
	.combout(\registerArray[3][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[3][31]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[3][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y43_N1
dffeas \registerArray[3][31] (
	.clk(clk),
	.d(\registerArray[3][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][31] .is_wysiwyg = "true";
defparam \registerArray[3][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N24
cycloneive_lcell_comb \Mux32~14 (
// Equation(s):
// \Mux32~14_combout  = (cuifregT_01 & ((cuifregT_1 & ((\registerArray[3][31]~q ))) # (!cuifregT_1 & (\registerArray[1][31]~q ))))

	.dataa(\registerArray[1][31]~q ),
	.datab(\registerArray[3][31]~q ),
	.datac(cuifregT_1),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux32~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~14 .lut_mask = 16'hCA00;
defparam \Mux32~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N12
cycloneive_lcell_comb \Mux32~15 (
// Equation(s):
// \Mux32~15_combout  = (\Mux32~14_combout ) # ((cuifregT_1 & (!cuifregT_01 & \registerArray[2][31]~q )))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\registerArray[2][31]~q ),
	.datad(\Mux32~14_combout ),
	.cin(gnd),
	.combout(\Mux32~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~15 .lut_mask = 16'hFF20;
defparam \Mux32~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y34_N16
cycloneive_lcell_comb \Mux32~16 (
// Equation(s):
// \Mux32~16_combout  = (cuifregT_3 & ((\Mux32~13_combout ) # ((cuifregT_2)))) # (!cuifregT_3 & (((!cuifregT_2 & \Mux32~15_combout ))))

	.dataa(cuifregT_3),
	.datab(\Mux32~13_combout ),
	.datac(cuifregT_2),
	.datad(\Mux32~15_combout ),
	.cin(gnd),
	.combout(\Mux32~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~16 .lut_mask = 16'hADA8;
defparam \Mux32~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N3
dffeas \registerArray[7][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][30] .is_wysiwyg = "true";
defparam \registerArray[7][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N9
dffeas \registerArray[4][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][30] .is_wysiwyg = "true";
defparam \registerArray[4][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N24
cycloneive_lcell_comb \Mux33~2 (
// Equation(s):
// \Mux33~2_combout  = (cuifregT_01 & ((\registerArray[5][30]~q ) # ((cuifregT_1)))) # (!cuifregT_01 & (((\registerArray[4][30]~q  & !cuifregT_1))))

	.dataa(\registerArray[5][30]~q ),
	.datab(\registerArray[4][30]~q ),
	.datac(cuifregT_0),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux33~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~2 .lut_mask = 16'hF0AC;
defparam \Mux33~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N2
cycloneive_lcell_comb \Mux33~3 (
// Equation(s):
// \Mux33~3_combout  = (cuifregT_1 & ((\Mux33~2_combout  & ((\registerArray[7][30]~q ))) # (!\Mux33~2_combout  & (\registerArray[6][30]~q )))) # (!cuifregT_1 & (((\Mux33~2_combout ))))

	.dataa(\registerArray[6][30]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[7][30]~q ),
	.datad(\Mux33~2_combout ),
	.cin(gnd),
	.combout(\Mux33~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~3 .lut_mask = 16'hF388;
defparam \Mux33~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N11
dffeas \registerArray[2][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][30] .is_wysiwyg = "true";
defparam \registerArray[2][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N13
dffeas \registerArray[1][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][30] .is_wysiwyg = "true";
defparam \registerArray[1][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N12
cycloneive_lcell_comb \Mux33~4 (
// Equation(s):
// \Mux33~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][30]~q )) # (!cuifregT_1 & ((\registerArray[1][30]~q )))))

	.dataa(\registerArray[3][30]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[1][30]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux33~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~4 .lut_mask = 16'hB800;
defparam \Mux33~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N10
cycloneive_lcell_comb \Mux33~5 (
// Equation(s):
// \Mux33~5_combout  = (\Mux33~4_combout ) # ((!cuifregT_01 & (cuifregT_1 & \registerArray[2][30]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[2][30]~q ),
	.datad(\Mux33~4_combout ),
	.cin(gnd),
	.combout(\Mux33~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~5 .lut_mask = 16'hFF40;
defparam \Mux33~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N4
cycloneive_lcell_comb \Mux33~6 (
// Equation(s):
// \Mux33~6_combout  = (cuifregT_3 & (cuifregT_2)) # (!cuifregT_3 & ((cuifregT_2 & (\Mux33~3_combout )) # (!cuifregT_2 & ((\Mux33~5_combout )))))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\Mux33~3_combout ),
	.datad(\Mux33~5_combout ),
	.cin(gnd),
	.combout(\Mux33~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~6 .lut_mask = 16'hD9C8;
defparam \Mux33~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N13
dffeas \registerArray[9][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][30] .is_wysiwyg = "true";
defparam \registerArray[9][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N27
dffeas \registerArray[11][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][30] .is_wysiwyg = "true";
defparam \registerArray[11][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N13
dffeas \registerArray[8][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][30] .is_wysiwyg = "true";
defparam \registerArray[8][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N12
cycloneive_lcell_comb \Mux33~0 (
// Equation(s):
// \Mux33~0_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & (\registerArray[10][30]~q )) # (!cuifregT_1 & ((\registerArray[8][30]~q )))))

	.dataa(\registerArray[10][30]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[8][30]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux33~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~0 .lut_mask = 16'hEE30;
defparam \Mux33~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N26
cycloneive_lcell_comb \Mux33~1 (
// Equation(s):
// \Mux33~1_combout  = (cuifregT_01 & ((\Mux33~0_combout  & ((\registerArray[11][30]~q ))) # (!\Mux33~0_combout  & (\registerArray[9][30]~q )))) # (!cuifregT_01 & (((\Mux33~0_combout ))))

	.dataa(\registerArray[9][30]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[11][30]~q ),
	.datad(\Mux33~0_combout ),
	.cin(gnd),
	.combout(\Mux33~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~1 .lut_mask = 16'hF388;
defparam \Mux33~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N19
dffeas \registerArray[14][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][30] .is_wysiwyg = "true";
defparam \registerArray[14][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N7
dffeas \registerArray[15][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][30] .is_wysiwyg = "true";
defparam \registerArray[15][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N13
dffeas \registerArray[12][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][30] .is_wysiwyg = "true";
defparam \registerArray[12][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N12
cycloneive_lcell_comb \Mux33~7 (
// Equation(s):
// \Mux33~7_combout  = (cuifregT_01 & ((\registerArray[13][30]~q ) # ((cuifregT_1)))) # (!cuifregT_01 & (((\registerArray[12][30]~q  & !cuifregT_1))))

	.dataa(\registerArray[13][30]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[12][30]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux33~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~7 .lut_mask = 16'hCCB8;
defparam \Mux33~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N6
cycloneive_lcell_comb \Mux33~8 (
// Equation(s):
// \Mux33~8_combout  = (cuifregT_1 & ((\Mux33~7_combout  & ((\registerArray[15][30]~q ))) # (!\Mux33~7_combout  & (\registerArray[14][30]~q )))) # (!cuifregT_1 & (((\Mux33~7_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[14][30]~q ),
	.datac(\registerArray[15][30]~q ),
	.datad(\Mux33~7_combout ),
	.cin(gnd),
	.combout(\Mux33~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~8 .lut_mask = 16'hF588;
defparam \Mux33~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N17
dffeas \registerArray[27][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][30] .is_wysiwyg = "true";
defparam \registerArray[27][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N23
dffeas \registerArray[31][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][30] .is_wysiwyg = "true";
defparam \registerArray[31][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N13
dffeas \registerArray[19][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][30] .is_wysiwyg = "true";
defparam \registerArray[19][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N12
cycloneive_lcell_comb \Mux33~17 (
// Equation(s):
// \Mux33~17_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[23][30]~q )) # (!cuifregT_2 & ((\registerArray[19][30]~q )))))

	.dataa(\registerArray[23][30]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[19][30]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux33~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~17 .lut_mask = 16'hEE30;
defparam \Mux33~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N22
cycloneive_lcell_comb \Mux33~18 (
// Equation(s):
// \Mux33~18_combout  = (cuifregT_3 & ((\Mux33~17_combout  & ((\registerArray[31][30]~q ))) # (!\Mux33~17_combout  & (\registerArray[27][30]~q )))) # (!cuifregT_3 & (((\Mux33~17_combout ))))

	.dataa(\registerArray[27][30]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[31][30]~q ),
	.datad(\Mux33~17_combout ),
	.cin(gnd),
	.combout(\Mux33~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~18 .lut_mask = 16'hF388;
defparam \Mux33~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y41_N5
dffeas \registerArray[25][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][30] .is_wysiwyg = "true";
defparam \registerArray[25][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N15
dffeas \registerArray[29][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][30] .is_wysiwyg = "true";
defparam \registerArray[29][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y42_N1
dffeas \registerArray[21][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][30] .is_wysiwyg = "true";
defparam \registerArray[21][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N25
dffeas \registerArray[17][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][30] .is_wysiwyg = "true";
defparam \registerArray[17][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N24
cycloneive_lcell_comb \Mux33~10 (
// Equation(s):
// \Mux33~10_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[21][30]~q )) # (!cuifregT_2 & ((\registerArray[17][30]~q )))))

	.dataa(cuifregT_3),
	.datab(\registerArray[21][30]~q ),
	.datac(\registerArray[17][30]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux33~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~10 .lut_mask = 16'hEE50;
defparam \Mux33~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N14
cycloneive_lcell_comb \Mux33~11 (
// Equation(s):
// \Mux33~11_combout  = (cuifregT_3 & ((\Mux33~10_combout  & ((\registerArray[29][30]~q ))) # (!\Mux33~10_combout  & (\registerArray[25][30]~q )))) # (!cuifregT_3 & (((\Mux33~10_combout ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[25][30]~q ),
	.datac(\registerArray[29][30]~q ),
	.datad(\Mux33~10_combout ),
	.cin(gnd),
	.combout(\Mux33~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~11 .lut_mask = 16'hF588;
defparam \Mux33~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N19
dffeas \registerArray[22][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][30] .is_wysiwyg = "true";
defparam \registerArray[22][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N11
dffeas \registerArray[30][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][30] .is_wysiwyg = "true";
defparam \registerArray[30][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N17
dffeas \registerArray[18][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][30] .is_wysiwyg = "true";
defparam \registerArray[18][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N16
cycloneive_lcell_comb \Mux33~12 (
// Equation(s):
// \Mux33~12_combout  = (cuifregT_3 & ((\registerArray[26][30]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[18][30]~q  & !cuifregT_2))))

	.dataa(\registerArray[26][30]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[18][30]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux33~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~12 .lut_mask = 16'hCCB8;
defparam \Mux33~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N10
cycloneive_lcell_comb \Mux33~13 (
// Equation(s):
// \Mux33~13_combout  = (cuifregT_2 & ((\Mux33~12_combout  & ((\registerArray[30][30]~q ))) # (!\Mux33~12_combout  & (\registerArray[22][30]~q )))) # (!cuifregT_2 & (((\Mux33~12_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[22][30]~q ),
	.datac(\registerArray[30][30]~q ),
	.datad(\Mux33~12_combout ),
	.cin(gnd),
	.combout(\Mux33~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~13 .lut_mask = 16'hF588;
defparam \Mux33~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N8
cycloneive_lcell_comb \registerArray[20][30]~feeder (
// Equation(s):
// \registerArray[20][30]~feeder_combout  = \Mux38~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux382),
	.cin(gnd),
	.combout(\registerArray[20][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[20][30]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[20][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y44_N9
dffeas \registerArray[20][30] (
	.clk(clk),
	.d(\registerArray[20][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][30] .is_wysiwyg = "true";
defparam \registerArray[20][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N4
cycloneive_lcell_comb \registerArray[16][30]~feeder (
// Equation(s):
// \registerArray[16][30]~feeder_combout  = \Mux38~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux382),
	.cin(gnd),
	.combout(\registerArray[16][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[16][30]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[16][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N5
dffeas \registerArray[16][30] (
	.clk(clk),
	.d(\registerArray[16][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][30] .is_wysiwyg = "true";
defparam \registerArray[16][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N22
cycloneive_lcell_comb \Mux33~14 (
// Equation(s):
// \Mux33~14_combout  = (cuifregT_3 & ((\registerArray[24][30]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[16][30]~q  & !cuifregT_2))))

	.dataa(\registerArray[24][30]~q ),
	.datab(\registerArray[16][30]~q ),
	.datac(cuifregT_3),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux33~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~14 .lut_mask = 16'hF0AC;
defparam \Mux33~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N16
cycloneive_lcell_comb \Mux33~15 (
// Equation(s):
// \Mux33~15_combout  = (cuifregT_2 & ((\Mux33~14_combout  & (\registerArray[28][30]~q )) # (!\Mux33~14_combout  & ((\registerArray[20][30]~q ))))) # (!cuifregT_2 & (((\Mux33~14_combout ))))

	.dataa(\registerArray[28][30]~q ),
	.datab(\registerArray[20][30]~q ),
	.datac(cuifregT_2),
	.datad(\Mux33~14_combout ),
	.cin(gnd),
	.combout(\Mux33~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~15 .lut_mask = 16'hAFC0;
defparam \Mux33~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N20
cycloneive_lcell_comb \Mux33~16 (
// Equation(s):
// \Mux33~16_combout  = (cuifregT_1 & ((cuifregT_01) # ((\Mux33~13_combout )))) # (!cuifregT_1 & (!cuifregT_01 & ((\Mux33~15_combout ))))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\Mux33~13_combout ),
	.datad(\Mux33~15_combout ),
	.cin(gnd),
	.combout(\Mux33~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~16 .lut_mask = 16'hB9A8;
defparam \Mux33~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N5
dffeas \registerArray[23][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][29] .is_wysiwyg = "true";
defparam \registerArray[23][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N19
dffeas \registerArray[27][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][29] .is_wysiwyg = "true";
defparam \registerArray[27][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N9
dffeas \registerArray[19][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][29] .is_wysiwyg = "true";
defparam \registerArray[19][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N8
cycloneive_lcell_comb \Mux34~7 (
// Equation(s):
// \Mux34~7_combout  = (cuifregT_3 & ((\registerArray[27][29]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[19][29]~q  & !cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[27][29]~q ),
	.datac(\registerArray[19][29]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux34~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~7 .lut_mask = 16'hAAD8;
defparam \Mux34~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y30_N11
dffeas \registerArray[31][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][29] .is_wysiwyg = "true";
defparam \registerArray[31][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N10
cycloneive_lcell_comb \Mux34~8 (
// Equation(s):
// \Mux34~8_combout  = (\Mux34~7_combout  & (((\registerArray[31][29]~q ) # (!cuifregT_2)))) # (!\Mux34~7_combout  & (\registerArray[23][29]~q  & ((cuifregT_2))))

	.dataa(\registerArray[23][29]~q ),
	.datab(\Mux34~7_combout ),
	.datac(\registerArray[31][29]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux34~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~8 .lut_mask = 16'hE2CC;
defparam \Mux34~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y30_N5
dffeas \registerArray[21][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][29] .is_wysiwyg = "true";
defparam \registerArray[21][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N4
cycloneive_lcell_comb \registerArray[25][29]~feeder (
// Equation(s):
// \registerArray[25][29]~feeder_combout  = \Mux39~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux392),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[25][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[25][29]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[25][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N5
dffeas \registerArray[25][29] (
	.clk(clk),
	.d(\registerArray[25][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][29] .is_wysiwyg = "true";
defparam \registerArray[25][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N9
dffeas \registerArray[17][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][29] .is_wysiwyg = "true";
defparam \registerArray[17][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N8
cycloneive_lcell_comb \Mux34~0 (
// Equation(s):
// \Mux34~0_combout  = (cuifregT_3 & ((\registerArray[25][29]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[17][29]~q  & !cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[25][29]~q ),
	.datac(\registerArray[17][29]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux34~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~0 .lut_mask = 16'hAAD8;
defparam \Mux34~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N3
dffeas \registerArray[29][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][29] .is_wysiwyg = "true";
defparam \registerArray[29][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N2
cycloneive_lcell_comb \Mux34~1 (
// Equation(s):
// \Mux34~1_combout  = (\Mux34~0_combout  & (((\registerArray[29][29]~q ) # (!cuifregT_2)))) # (!\Mux34~0_combout  & (\registerArray[21][29]~q  & ((cuifregT_2))))

	.dataa(\registerArray[21][29]~q ),
	.datab(\Mux34~0_combout ),
	.datac(\registerArray[29][29]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux34~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~1 .lut_mask = 16'hE2CC;
defparam \Mux34~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y32_N31
dffeas \registerArray[28][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][29] .is_wysiwyg = "true";
defparam \registerArray[28][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N17
dffeas \registerArray[16][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][29] .is_wysiwyg = "true";
defparam \registerArray[16][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N16
cycloneive_lcell_comb \Mux34~4 (
// Equation(s):
// \Mux34~4_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[20][29]~q )) # (!cuifregT_2 & ((\registerArray[16][29]~q )))))

	.dataa(\registerArray[20][29]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[16][29]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux34~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~4 .lut_mask = 16'hEE30;
defparam \Mux34~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N30
cycloneive_lcell_comb \Mux34~5 (
// Equation(s):
// \Mux34~5_combout  = (cuifregT_3 & ((\Mux34~4_combout  & ((\registerArray[28][29]~q ))) # (!\Mux34~4_combout  & (\registerArray[24][29]~q )))) # (!cuifregT_3 & (((\Mux34~4_combout ))))

	.dataa(\registerArray[24][29]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[28][29]~q ),
	.datad(\Mux34~4_combout ),
	.cin(gnd),
	.combout(\Mux34~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~5 .lut_mask = 16'hF388;
defparam \Mux34~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N31
dffeas \registerArray[30][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][29] .is_wysiwyg = "true";
defparam \registerArray[30][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N28
cycloneive_lcell_comb \registerArray[22][29]~feeder (
// Equation(s):
// \registerArray[22][29]~feeder_combout  = \Mux39~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux392),
	.cin(gnd),
	.combout(\registerArray[22][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[22][29]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[22][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N29
dffeas \registerArray[22][29] (
	.clk(clk),
	.d(\registerArray[22][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][29] .is_wysiwyg = "true";
defparam \registerArray[22][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N29
dffeas \registerArray[18][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][29] .is_wysiwyg = "true";
defparam \registerArray[18][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N28
cycloneive_lcell_comb \Mux34~2 (
// Equation(s):
// \Mux34~2_combout  = (cuifregT_2 & ((\registerArray[22][29]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[18][29]~q  & !cuifregT_3))))

	.dataa(cuifregT_2),
	.datab(\registerArray[22][29]~q ),
	.datac(\registerArray[18][29]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux34~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~2 .lut_mask = 16'hAAD8;
defparam \Mux34~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N30
cycloneive_lcell_comb \Mux34~3 (
// Equation(s):
// \Mux34~3_combout  = (cuifregT_3 & ((\Mux34~2_combout  & ((\registerArray[30][29]~q ))) # (!\Mux34~2_combout  & (\registerArray[26][29]~q )))) # (!cuifregT_3 & (((\Mux34~2_combout ))))

	.dataa(\registerArray[26][29]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[30][29]~q ),
	.datad(\Mux34~2_combout ),
	.cin(gnd),
	.combout(\Mux34~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~3 .lut_mask = 16'hF388;
defparam \Mux34~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N24
cycloneive_lcell_comb \Mux34~6 (
// Equation(s):
// \Mux34~6_combout  = (cuifregT_1 & (((\Mux34~3_combout ) # (cuifregT_01)))) # (!cuifregT_1 & (\Mux34~5_combout  & ((!cuifregT_01))))

	.dataa(\Mux34~5_combout ),
	.datab(cuifregT_1),
	.datac(\Mux34~3_combout ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux34~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~6 .lut_mask = 16'hCCE2;
defparam \Mux34~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N1
dffeas \registerArray[6][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][29] .is_wysiwyg = "true";
defparam \registerArray[6][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N5
dffeas \registerArray[4][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][29] .is_wysiwyg = "true";
defparam \registerArray[4][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N4
cycloneive_lcell_comb \Mux34~10 (
// Equation(s):
// \Mux34~10_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[5][29]~q )) # (!cuifregT_01 & ((\registerArray[4][29]~q )))))

	.dataa(\registerArray[5][29]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[4][29]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux34~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~10 .lut_mask = 16'hEE30;
defparam \Mux34~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N31
dffeas \registerArray[7][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][29] .is_wysiwyg = "true";
defparam \registerArray[7][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N30
cycloneive_lcell_comb \Mux34~11 (
// Equation(s):
// \Mux34~11_combout  = (\Mux34~10_combout  & (((\registerArray[7][29]~q ) # (!cuifregT_1)))) # (!\Mux34~10_combout  & (\registerArray[6][29]~q  & ((cuifregT_1))))

	.dataa(\registerArray[6][29]~q ),
	.datab(\Mux34~10_combout ),
	.datac(\registerArray[7][29]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux34~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~11 .lut_mask = 16'hE2CC;
defparam \Mux34~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N15
dffeas \registerArray[14][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][29] .is_wysiwyg = "true";
defparam \registerArray[14][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N15
dffeas \registerArray[15][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][29] .is_wysiwyg = "true";
defparam \registerArray[15][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N13
dffeas \registerArray[13][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][29] .is_wysiwyg = "true";
defparam \registerArray[13][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N25
dffeas \registerArray[12][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][29] .is_wysiwyg = "true";
defparam \registerArray[12][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N24
cycloneive_lcell_comb \Mux34~17 (
// Equation(s):
// \Mux34~17_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[13][29]~q )) # (!cuifregT_01 & ((\registerArray[12][29]~q )))))

	.dataa(cuifregT_1),
	.datab(\registerArray[13][29]~q ),
	.datac(\registerArray[12][29]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux34~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~17 .lut_mask = 16'hEE50;
defparam \Mux34~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N14
cycloneive_lcell_comb \Mux34~18 (
// Equation(s):
// \Mux34~18_combout  = (cuifregT_1 & ((\Mux34~17_combout  & ((\registerArray[15][29]~q ))) # (!\Mux34~17_combout  & (\registerArray[14][29]~q )))) # (!cuifregT_1 & (((\Mux34~17_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[14][29]~q ),
	.datac(\registerArray[15][29]~q ),
	.datad(\Mux34~17_combout ),
	.cin(gnd),
	.combout(\Mux34~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~18 .lut_mask = 16'hF588;
defparam \Mux34~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N19
dffeas \registerArray[11][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][29] .is_wysiwyg = "true";
defparam \registerArray[11][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N25
dffeas \registerArray[8][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][29] .is_wysiwyg = "true";
defparam \registerArray[8][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N24
cycloneive_lcell_comb \Mux34~12 (
// Equation(s):
// \Mux34~12_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & (\registerArray[10][29]~q )) # (!cuifregT_1 & ((\registerArray[8][29]~q )))))

	.dataa(\registerArray[10][29]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[8][29]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux34~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~12 .lut_mask = 16'hEE30;
defparam \Mux34~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N18
cycloneive_lcell_comb \Mux34~13 (
// Equation(s):
// \Mux34~13_combout  = (cuifregT_01 & ((\Mux34~12_combout  & ((\registerArray[11][29]~q ))) # (!\Mux34~12_combout  & (\registerArray[9][29]~q )))) # (!cuifregT_01 & (((\Mux34~12_combout ))))

	.dataa(\registerArray[9][29]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[11][29]~q ),
	.datad(\Mux34~12_combout ),
	.cin(gnd),
	.combout(\Mux34~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~13 .lut_mask = 16'hF388;
defparam \Mux34~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N31
dffeas \registerArray[2][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][29] .is_wysiwyg = "true";
defparam \registerArray[2][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N4
cycloneive_lcell_comb \registerArray[3][29]~feeder (
// Equation(s):
// \registerArray[3][29]~feeder_combout  = \Mux39~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux392),
	.cin(gnd),
	.combout(\registerArray[3][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[3][29]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[3][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N5
dffeas \registerArray[3][29] (
	.clk(clk),
	.d(\registerArray[3][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][29] .is_wysiwyg = "true";
defparam \registerArray[3][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N25
dffeas \registerArray[1][29] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux392),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][29] .is_wysiwyg = "true";
defparam \registerArray[1][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N24
cycloneive_lcell_comb \Mux34~14 (
// Equation(s):
// \Mux34~14_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][29]~q )) # (!cuifregT_1 & ((\registerArray[1][29]~q )))))

	.dataa(cuifregT_0),
	.datab(\registerArray[3][29]~q ),
	.datac(\registerArray[1][29]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux34~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~14 .lut_mask = 16'h88A0;
defparam \Mux34~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N30
cycloneive_lcell_comb \Mux34~15 (
// Equation(s):
// \Mux34~15_combout  = (\Mux34~14_combout ) # ((!cuifregT_01 & (cuifregT_1 & \registerArray[2][29]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[2][29]~q ),
	.datad(\Mux34~14_combout ),
	.cin(gnd),
	.combout(\Mux34~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~15 .lut_mask = 16'hFF40;
defparam \Mux34~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N24
cycloneive_lcell_comb \Mux34~16 (
// Equation(s):
// \Mux34~16_combout  = (cuifregT_3 & ((cuifregT_2) # ((\Mux34~13_combout )))) # (!cuifregT_3 & (!cuifregT_2 & ((\Mux34~15_combout ))))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\Mux34~13_combout ),
	.datad(\Mux34~15_combout ),
	.cin(gnd),
	.combout(\Mux34~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~16 .lut_mask = 16'hB9A8;
defparam \Mux34~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y43_N13
dffeas \registerArray[9][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][28] .is_wysiwyg = "true";
defparam \registerArray[9][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y43_N3
dffeas \registerArray[10][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][28] .is_wysiwyg = "true";
defparam \registerArray[10][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N5
dffeas \registerArray[8][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][28] .is_wysiwyg = "true";
defparam \registerArray[8][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N4
cycloneive_lcell_comb \Mux35~0 (
// Equation(s):
// \Mux35~0_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & (\registerArray[10][28]~q )) # (!cuifregT_1 & ((\registerArray[8][28]~q )))))

	.dataa(cuifregT_0),
	.datab(\registerArray[10][28]~q ),
	.datac(\registerArray[8][28]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux35~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~0 .lut_mask = 16'hEE50;
defparam \Mux35~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N23
dffeas \registerArray[11][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][28] .is_wysiwyg = "true";
defparam \registerArray[11][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N22
cycloneive_lcell_comb \Mux35~1 (
// Equation(s):
// \Mux35~1_combout  = (\Mux35~0_combout  & (((\registerArray[11][28]~q ) # (!cuifregT_01)))) # (!\Mux35~0_combout  & (\registerArray[9][28]~q  & ((cuifregT_01))))

	.dataa(\registerArray[9][28]~q ),
	.datab(\Mux35~0_combout ),
	.datac(\registerArray[11][28]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux35~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~1 .lut_mask = 16'hE2CC;
defparam \Mux35~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N11
dffeas \registerArray[14][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][28] .is_wysiwyg = "true";
defparam \registerArray[14][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N11
dffeas \registerArray[15][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][28] .is_wysiwyg = "true";
defparam \registerArray[15][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N21
dffeas \registerArray[13][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][28] .is_wysiwyg = "true";
defparam \registerArray[13][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N29
dffeas \registerArray[12][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][28] .is_wysiwyg = "true";
defparam \registerArray[12][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N28
cycloneive_lcell_comb \Mux35~7 (
// Equation(s):
// \Mux35~7_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[13][28]~q )) # (!cuifregT_01 & ((\registerArray[12][28]~q )))))

	.dataa(cuifregT_1),
	.datab(\registerArray[13][28]~q ),
	.datac(\registerArray[12][28]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux35~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~7 .lut_mask = 16'hEE50;
defparam \Mux35~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N10
cycloneive_lcell_comb \Mux35~8 (
// Equation(s):
// \Mux35~8_combout  = (cuifregT_1 & ((\Mux35~7_combout  & ((\registerArray[15][28]~q ))) # (!\Mux35~7_combout  & (\registerArray[14][28]~q )))) # (!cuifregT_1 & (((\Mux35~7_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[14][28]~q ),
	.datac(\registerArray[15][28]~q ),
	.datad(\Mux35~7_combout ),
	.cin(gnd),
	.combout(\Mux35~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~8 .lut_mask = 16'hF588;
defparam \Mux35~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N7
dffeas \registerArray[7][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][28] .is_wysiwyg = "true";
defparam \registerArray[7][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N1
dffeas \registerArray[4][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][28] .is_wysiwyg = "true";
defparam \registerArray[4][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N0
cycloneive_lcell_comb \Mux35~2 (
// Equation(s):
// \Mux35~2_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[5][28]~q )) # (!cuifregT_01 & ((\registerArray[4][28]~q )))))

	.dataa(\registerArray[5][28]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[4][28]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux35~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~2 .lut_mask = 16'hEE30;
defparam \Mux35~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N6
cycloneive_lcell_comb \Mux35~3 (
// Equation(s):
// \Mux35~3_combout  = (cuifregT_1 & ((\Mux35~2_combout  & ((\registerArray[7][28]~q ))) # (!\Mux35~2_combout  & (\registerArray[6][28]~q )))) # (!cuifregT_1 & (((\Mux35~2_combout ))))

	.dataa(\registerArray[6][28]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[7][28]~q ),
	.datad(\Mux35~2_combout ),
	.cin(gnd),
	.combout(\Mux35~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~3 .lut_mask = 16'hF388;
defparam \Mux35~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N15
dffeas \registerArray[2][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][28] .is_wysiwyg = "true";
defparam \registerArray[2][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N18
cycloneive_lcell_comb \registerArray[3][28]~feeder (
// Equation(s):
// \registerArray[3][28]~feeder_combout  = \Mux40~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux402),
	.cin(gnd),
	.combout(\registerArray[3][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[3][28]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[3][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y38_N19
dffeas \registerArray[3][28] (
	.clk(clk),
	.d(\registerArray[3][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][28] .is_wysiwyg = "true";
defparam \registerArray[3][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N25
dffeas \registerArray[1][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][28] .is_wysiwyg = "true";
defparam \registerArray[1][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N24
cycloneive_lcell_comb \Mux35~4 (
// Equation(s):
// \Mux35~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][28]~q )) # (!cuifregT_1 & ((\registerArray[1][28]~q )))))

	.dataa(cuifregT_1),
	.datab(\registerArray[3][28]~q ),
	.datac(\registerArray[1][28]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux35~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~4 .lut_mask = 16'hD800;
defparam \Mux35~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N14
cycloneive_lcell_comb \Mux35~5 (
// Equation(s):
// \Mux35~5_combout  = (\Mux35~4_combout ) # ((cuifregT_1 & (!cuifregT_01 & \registerArray[2][28]~q )))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\registerArray[2][28]~q ),
	.datad(\Mux35~4_combout ),
	.cin(gnd),
	.combout(\Mux35~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~5 .lut_mask = 16'hFF20;
defparam \Mux35~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N6
cycloneive_lcell_comb \Mux35~6 (
// Equation(s):
// \Mux35~6_combout  = (cuifregT_2 & ((cuifregT_3) # ((\Mux35~3_combout )))) # (!cuifregT_2 & (!cuifregT_3 & ((\Mux35~5_combout ))))

	.dataa(cuifregT_2),
	.datab(cuifregT_3),
	.datac(\Mux35~3_combout ),
	.datad(\Mux35~5_combout ),
	.cin(gnd),
	.combout(\Mux35~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~6 .lut_mask = 16'hB9A8;
defparam \Mux35~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N24
cycloneive_lcell_comb \registerArray[23][28]~feeder (
// Equation(s):
// \registerArray[23][28]~feeder_combout  = \Mux40~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux402),
	.cin(gnd),
	.combout(\registerArray[23][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[23][28]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[23][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N25
dffeas \registerArray[23][28] (
	.clk(clk),
	.d(\registerArray[23][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][28] .is_wysiwyg = "true";
defparam \registerArray[23][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N29
dffeas \registerArray[19][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][28] .is_wysiwyg = "true";
defparam \registerArray[19][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N28
cycloneive_lcell_comb \Mux35~17 (
// Equation(s):
// \Mux35~17_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[23][28]~q )) # (!cuifregT_2 & ((\registerArray[19][28]~q )))))

	.dataa(cuifregT_3),
	.datab(\registerArray[23][28]~q ),
	.datac(\registerArray[19][28]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux35~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~17 .lut_mask = 16'hEE50;
defparam \Mux35~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y32_N3
dffeas \registerArray[31][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][28] .is_wysiwyg = "true";
defparam \registerArray[31][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y38_N28
cycloneive_lcell_comb \registerArray[27][28]~feeder (
// Equation(s):
// \registerArray[27][28]~feeder_combout  = \Mux40~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux402),
	.cin(gnd),
	.combout(\registerArray[27][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[27][28]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[27][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y38_N29
dffeas \registerArray[27][28] (
	.clk(clk),
	.d(\registerArray[27][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][28] .is_wysiwyg = "true";
defparam \registerArray[27][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N2
cycloneive_lcell_comb \Mux35~18 (
// Equation(s):
// \Mux35~18_combout  = (cuifregT_3 & ((\Mux35~17_combout  & (\registerArray[31][28]~q )) # (!\Mux35~17_combout  & ((\registerArray[27][28]~q ))))) # (!cuifregT_3 & (\Mux35~17_combout ))

	.dataa(cuifregT_3),
	.datab(\Mux35~17_combout ),
	.datac(\registerArray[31][28]~q ),
	.datad(\registerArray[27][28]~q ),
	.cin(gnd),
	.combout(\Mux35~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~18 .lut_mask = 16'hE6C4;
defparam \Mux35~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N21
dffeas \registerArray[20][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][28] .is_wysiwyg = "true";
defparam \registerArray[20][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y34_N15
dffeas \registerArray[28][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][28] .is_wysiwyg = "true";
defparam \registerArray[28][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N14
cycloneive_lcell_comb \Mux35~15 (
// Equation(s):
// \Mux35~15_combout  = (\Mux35~14_combout  & (((\registerArray[28][28]~q ) # (!cuifregT_2)))) # (!\Mux35~14_combout  & (\registerArray[20][28]~q  & ((cuifregT_2))))

	.dataa(\Mux35~14_combout ),
	.datab(\registerArray[20][28]~q ),
	.datac(\registerArray[28][28]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux35~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~15 .lut_mask = 16'hE4AA;
defparam \Mux35~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N0
cycloneive_lcell_comb \Decoder0~63 (
// Equation(s):
// \Decoder0~63_combout  = (\Mux3~1_combout  & (!\Mux2~1_combout  & (!\Mux4~1_combout  & \Decoder0~50_combout )))

	.dataa(Mux310),
	.datab(Mux210),
	.datac(Mux410),
	.datad(\Decoder0~50_combout ),
	.cin(gnd),
	.combout(\Decoder0~63_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~63 .lut_mask = 16'h0200;
defparam \Decoder0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N23
dffeas \registerArray[26][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][28] .is_wysiwyg = "true";
defparam \registerArray[26][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N9
dffeas \registerArray[18][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][28] .is_wysiwyg = "true";
defparam \registerArray[18][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N8
cycloneive_lcell_comb \Mux35~12 (
// Equation(s):
// \Mux35~12_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[26][28]~q )) # (!cuifregT_3 & ((\registerArray[18][28]~q )))))

	.dataa(cuifregT_2),
	.datab(\registerArray[26][28]~q ),
	.datac(\registerArray[18][28]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux35~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~12 .lut_mask = 16'hEE50;
defparam \Mux35~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N27
dffeas \registerArray[30][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][28] .is_wysiwyg = "true";
defparam \registerArray[30][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N26
cycloneive_lcell_comb \Mux35~13 (
// Equation(s):
// \Mux35~13_combout  = (\Mux35~12_combout  & (((\registerArray[30][28]~q ) # (!cuifregT_2)))) # (!\Mux35~12_combout  & (\registerArray[22][28]~q  & ((cuifregT_2))))

	.dataa(\registerArray[22][28]~q ),
	.datab(\Mux35~12_combout ),
	.datac(\registerArray[30][28]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux35~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~13 .lut_mask = 16'hE2CC;
defparam \Mux35~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N14
cycloneive_lcell_comb \Mux35~16 (
// Equation(s):
// \Mux35~16_combout  = (cuifregT_1 & (((\Mux35~13_combout ) # (cuifregT_01)))) # (!cuifregT_1 & (\Mux35~15_combout  & ((!cuifregT_01))))

	.dataa(\Mux35~15_combout ),
	.datab(cuifregT_1),
	.datac(\Mux35~13_combout ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux35~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~16 .lut_mask = 16'hCCE2;
defparam \Mux35~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N12
cycloneive_lcell_comb \registerArray[29][28]~feeder (
// Equation(s):
// \registerArray[29][28]~feeder_combout  = \Mux40~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux402),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[29][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[29][28]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[29][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N13
dffeas \registerArray[29][28] (
	.clk(clk),
	.d(\registerArray[29][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][28] .is_wysiwyg = "true";
defparam \registerArray[29][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N20
cycloneive_lcell_comb \registerArray[25][28]~feeder (
// Equation(s):
// \registerArray[25][28]~feeder_combout  = \Mux40~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux402),
	.cin(gnd),
	.combout(\registerArray[25][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[25][28]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[25][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N21
dffeas \registerArray[25][28] (
	.clk(clk),
	.d(\registerArray[25][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][28] .is_wysiwyg = "true";
defparam \registerArray[25][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N28
cycloneive_lcell_comb \registerArray[21][28]~feeder (
// Equation(s):
// \registerArray[21][28]~feeder_combout  = \Mux40~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux402),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[21][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[21][28]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[21][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N29
dffeas \registerArray[21][28] (
	.clk(clk),
	.d(\registerArray[21][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][28] .is_wysiwyg = "true";
defparam \registerArray[21][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N2
cycloneive_lcell_comb \Mux35~10 (
// Equation(s):
// \Mux35~10_combout  = (cuifregT_2 & (((\registerArray[21][28]~q ) # (cuifregT_3)))) # (!cuifregT_2 & (\registerArray[17][28]~q  & ((!cuifregT_3))))

	.dataa(\registerArray[17][28]~q ),
	.datab(\registerArray[21][28]~q ),
	.datac(cuifregT_2),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux35~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~10 .lut_mask = 16'hF0CA;
defparam \Mux35~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N26
cycloneive_lcell_comb \Mux35~11 (
// Equation(s):
// \Mux35~11_combout  = (cuifregT_3 & ((\Mux35~10_combout  & (\registerArray[29][28]~q )) # (!\Mux35~10_combout  & ((\registerArray[25][28]~q ))))) # (!cuifregT_3 & (((\Mux35~10_combout ))))

	.dataa(\registerArray[29][28]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[25][28]~q ),
	.datad(\Mux35~10_combout ),
	.cin(gnd),
	.combout(\Mux35~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~11 .lut_mask = 16'hBBC0;
defparam \Mux35~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N7
dffeas \registerArray[5][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][27] .is_wysiwyg = "true";
defparam \registerArray[5][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N1
dffeas \registerArray[4][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][27] .is_wysiwyg = "true";
defparam \registerArray[4][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N0
cycloneive_lcell_comb \Mux36~0 (
// Equation(s):
// \Mux36~0_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[5][27]~q )) # (!cuifregT_01 & ((\registerArray[4][27]~q )))))

	.dataa(cuifregT_1),
	.datab(\registerArray[5][27]~q ),
	.datac(\registerArray[4][27]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux36~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~0 .lut_mask = 16'hEE50;
defparam \Mux36~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N25
dffeas \registerArray[7][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][27] .is_wysiwyg = "true";
defparam \registerArray[7][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N11
dffeas \registerArray[6][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][27] .is_wysiwyg = "true";
defparam \registerArray[6][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N24
cycloneive_lcell_comb \Mux36~1 (
// Equation(s):
// \Mux36~1_combout  = (cuifregT_1 & ((\Mux36~0_combout  & (\registerArray[7][27]~q )) # (!\Mux36~0_combout  & ((\registerArray[6][27]~q ))))) # (!cuifregT_1 & (\Mux36~0_combout ))

	.dataa(cuifregT_1),
	.datab(\Mux36~0_combout ),
	.datac(\registerArray[7][27]~q ),
	.datad(\registerArray[6][27]~q ),
	.cin(gnd),
	.combout(\Mux36~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~1 .lut_mask = 16'hE6C4;
defparam \Mux36~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N31
dffeas \registerArray[14][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][27] .is_wysiwyg = "true";
defparam \registerArray[14][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N25
dffeas \registerArray[13][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][27] .is_wysiwyg = "true";
defparam \registerArray[13][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N5
dffeas \registerArray[12][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][27] .is_wysiwyg = "true";
defparam \registerArray[12][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N4
cycloneive_lcell_comb \Mux36~7 (
// Equation(s):
// \Mux36~7_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[13][27]~q )) # (!cuifregT_01 & ((\registerArray[12][27]~q )))))

	.dataa(cuifregT_1),
	.datab(\registerArray[13][27]~q ),
	.datac(\registerArray[12][27]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux36~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~7 .lut_mask = 16'hEE50;
defparam \Mux36~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y36_N27
dffeas \registerArray[15][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][27] .is_wysiwyg = "true";
defparam \registerArray[15][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N26
cycloneive_lcell_comb \Mux36~8 (
// Equation(s):
// \Mux36~8_combout  = (\Mux36~7_combout  & (((\registerArray[15][27]~q ) # (!cuifregT_1)))) # (!\Mux36~7_combout  & (\registerArray[14][27]~q  & ((cuifregT_1))))

	.dataa(\registerArray[14][27]~q ),
	.datab(\Mux36~7_combout ),
	.datac(\registerArray[15][27]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux36~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~8 .lut_mask = 16'hE2CC;
defparam \Mux36~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N27
dffeas \registerArray[2][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][27] .is_wysiwyg = "true";
defparam \registerArray[2][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N23
dffeas \registerArray[3][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][27] .is_wysiwyg = "true";
defparam \registerArray[3][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N17
dffeas \registerArray[1][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][27] .is_wysiwyg = "true";
defparam \registerArray[1][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N16
cycloneive_lcell_comb \Mux36~4 (
// Equation(s):
// \Mux36~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][27]~q )) # (!cuifregT_1 & ((\registerArray[1][27]~q )))))

	.dataa(cuifregT_0),
	.datab(\registerArray[3][27]~q ),
	.datac(\registerArray[1][27]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux36~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~4 .lut_mask = 16'h88A0;
defparam \Mux36~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N26
cycloneive_lcell_comb \Mux36~5 (
// Equation(s):
// \Mux36~5_combout  = (\Mux36~4_combout ) # ((!cuifregT_01 & (cuifregT_1 & \registerArray[2][27]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[2][27]~q ),
	.datad(\Mux36~4_combout ),
	.cin(gnd),
	.combout(\Mux36~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~5 .lut_mask = 16'hFF40;
defparam \Mux36~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N25
dffeas \registerArray[9][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][27] .is_wysiwyg = "true";
defparam \registerArray[9][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N3
dffeas \registerArray[11][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][27] .is_wysiwyg = "true";
defparam \registerArray[11][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N17
dffeas \registerArray[8][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][27] .is_wysiwyg = "true";
defparam \registerArray[8][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N16
cycloneive_lcell_comb \Mux36~2 (
// Equation(s):
// \Mux36~2_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & (\registerArray[10][27]~q )) # (!cuifregT_1 & ((\registerArray[8][27]~q )))))

	.dataa(\registerArray[10][27]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[8][27]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux36~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~2 .lut_mask = 16'hEE30;
defparam \Mux36~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N2
cycloneive_lcell_comb \Mux36~3 (
// Equation(s):
// \Mux36~3_combout  = (cuifregT_01 & ((\Mux36~2_combout  & ((\registerArray[11][27]~q ))) # (!\Mux36~2_combout  & (\registerArray[9][27]~q )))) # (!cuifregT_01 & (((\Mux36~2_combout ))))

	.dataa(cuifregT_0),
	.datab(\registerArray[9][27]~q ),
	.datac(\registerArray[11][27]~q ),
	.datad(\Mux36~2_combout ),
	.cin(gnd),
	.combout(\Mux36~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~3 .lut_mask = 16'hF588;
defparam \Mux36~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N10
cycloneive_lcell_comb \Mux36~6 (
// Equation(s):
// \Mux36~6_combout  = (cuifregT_2 & (cuifregT_3)) # (!cuifregT_2 & ((cuifregT_3 & ((\Mux36~3_combout ))) # (!cuifregT_3 & (\Mux36~5_combout ))))

	.dataa(cuifregT_2),
	.datab(cuifregT_3),
	.datac(\Mux36~5_combout ),
	.datad(\Mux36~3_combout ),
	.cin(gnd),
	.combout(\Mux36~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~6 .lut_mask = 16'hDC98;
defparam \Mux36~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N12
cycloneive_lcell_comb \registerArray[21][27]~feeder (
// Equation(s):
// \registerArray[21][27]~feeder_combout  = \Mux41~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux412),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[21][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[21][27]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[21][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N13
dffeas \registerArray[21][27] (
	.clk(clk),
	.d(\registerArray[21][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][27] .is_wysiwyg = "true";
defparam \registerArray[21][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N19
dffeas \registerArray[29][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][27] .is_wysiwyg = "true";
defparam \registerArray[29][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N26
cycloneive_lcell_comb \registerArray[25][27]~feeder (
// Equation(s):
// \registerArray[25][27]~feeder_combout  = \Mux41~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux412),
	.cin(gnd),
	.combout(\registerArray[25][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[25][27]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[25][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N27
dffeas \registerArray[25][27] (
	.clk(clk),
	.d(\registerArray[25][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][27] .is_wysiwyg = "true";
defparam \registerArray[25][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N24
cycloneive_lcell_comb \registerArray[17][27]~feeder (
// Equation(s):
// \registerArray[17][27]~feeder_combout  = \Mux41~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux412),
	.cin(gnd),
	.combout(\registerArray[17][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[17][27]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[17][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N25
dffeas \registerArray[17][27] (
	.clk(clk),
	.d(\registerArray[17][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][27] .is_wysiwyg = "true";
defparam \registerArray[17][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N16
cycloneive_lcell_comb \Mux36~10 (
// Equation(s):
// \Mux36~10_combout  = (cuifregT_3 & ((\registerArray[25][27]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((!cuifregT_2 & \registerArray[17][27]~q ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[25][27]~q ),
	.datac(cuifregT_2),
	.datad(\registerArray[17][27]~q ),
	.cin(gnd),
	.combout(\Mux36~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~10 .lut_mask = 16'hADA8;
defparam \Mux36~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N18
cycloneive_lcell_comb \Mux36~11 (
// Equation(s):
// \Mux36~11_combout  = (cuifregT_2 & ((\Mux36~10_combout  & ((\registerArray[29][27]~q ))) # (!\Mux36~10_combout  & (\registerArray[21][27]~q )))) # (!cuifregT_2 & (((\Mux36~10_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[21][27]~q ),
	.datac(\registerArray[29][27]~q ),
	.datad(\Mux36~10_combout ),
	.cin(gnd),
	.combout(\Mux36~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~11 .lut_mask = 16'hF588;
defparam \Mux36~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N5
dffeas \registerArray[18][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][27] .is_wysiwyg = "true";
defparam \registerArray[18][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N4
cycloneive_lcell_comb \Mux36~12 (
// Equation(s):
// \Mux36~12_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[22][27]~q )) # (!cuifregT_2 & ((\registerArray[18][27]~q )))))

	.dataa(\registerArray[22][27]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[18][27]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux36~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~12 .lut_mask = 16'hEE30;
defparam \Mux36~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N23
dffeas \registerArray[30][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][27] .is_wysiwyg = "true";
defparam \registerArray[30][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N22
cycloneive_lcell_comb \Mux36~13 (
// Equation(s):
// \Mux36~13_combout  = (\Mux36~12_combout  & (((\registerArray[30][27]~q ) # (!cuifregT_3)))) # (!\Mux36~12_combout  & (\registerArray[26][27]~q  & ((cuifregT_3))))

	.dataa(\registerArray[26][27]~q ),
	.datab(\Mux36~12_combout ),
	.datac(\registerArray[30][27]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux36~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~13 .lut_mask = 16'hE2CC;
defparam \Mux36~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N21
dffeas \registerArray[24][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][27] .is_wysiwyg = "true";
defparam \registerArray[24][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y34_N17
dffeas \registerArray[28][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][27] .is_wysiwyg = "true";
defparam \registerArray[28][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N16
cycloneive_lcell_comb \Mux36~15 (
// Equation(s):
// \Mux36~15_combout  = (\Mux36~14_combout  & (((\registerArray[28][27]~q ) # (!cuifregT_3)))) # (!\Mux36~14_combout  & (\registerArray[24][27]~q  & ((cuifregT_3))))

	.dataa(\Mux36~14_combout ),
	.datab(\registerArray[24][27]~q ),
	.datac(\registerArray[28][27]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux36~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~15 .lut_mask = 16'hE4AA;
defparam \Mux36~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N14
cycloneive_lcell_comb \Mux36~16 (
// Equation(s):
// \Mux36~16_combout  = (cuifregT_1 & ((cuifregT_01) # ((\Mux36~13_combout )))) # (!cuifregT_1 & (!cuifregT_01 & ((\Mux36~15_combout ))))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\Mux36~13_combout ),
	.datad(\Mux36~15_combout ),
	.cin(gnd),
	.combout(\Mux36~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~16 .lut_mask = 16'hB9A8;
defparam \Mux36~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N17
dffeas \registerArray[27][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][27] .is_wysiwyg = "true";
defparam \registerArray[27][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N23
dffeas \registerArray[19][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][27] .is_wysiwyg = "true";
defparam \registerArray[19][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N22
cycloneive_lcell_comb \Mux36~17 (
// Equation(s):
// \Mux36~17_combout  = (cuifregT_3 & ((\registerArray[27][27]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[19][27]~q  & !cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[27][27]~q ),
	.datac(\registerArray[19][27]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux36~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~17 .lut_mask = 16'hAAD8;
defparam \Mux36~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N22
cycloneive_lcell_comb \registerArray[23][27]~feeder (
// Equation(s):
// \registerArray[23][27]~feeder_combout  = \Mux41~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux412),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[23][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[23][27]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[23][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N23
dffeas \registerArray[23][27] (
	.clk(clk),
	.d(\registerArray[23][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][27] .is_wysiwyg = "true";
defparam \registerArray[23][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N17
dffeas \registerArray[31][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][27] .is_wysiwyg = "true";
defparam \registerArray[31][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N16
cycloneive_lcell_comb \Mux36~18 (
// Equation(s):
// \Mux36~18_combout  = (\Mux36~17_combout  & (((\registerArray[31][27]~q ) # (!cuifregT_2)))) # (!\Mux36~17_combout  & (\registerArray[23][27]~q  & ((cuifregT_2))))

	.dataa(\Mux36~17_combout ),
	.datab(\registerArray[23][27]~q ),
	.datac(\registerArray[31][27]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux36~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~18 .lut_mask = 16'hE4AA;
defparam \Mux36~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N26
cycloneive_lcell_comb \registerArray[14][26]~feeder (
// Equation(s):
// \registerArray[14][26]~feeder_combout  = \Mux42~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux422),
	.cin(gnd),
	.combout(\registerArray[14][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][26]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[14][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N27
dffeas \registerArray[14][26] (
	.clk(clk),
	.d(\registerArray[14][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][26] .is_wysiwyg = "true";
defparam \registerArray[14][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N23
dffeas \registerArray[15][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][26] .is_wysiwyg = "true";
defparam \registerArray[15][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N8
cycloneive_lcell_comb \registerArray[13][26]~feeder (
// Equation(s):
// \registerArray[13][26]~feeder_combout  = \Mux42~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux422),
	.cin(gnd),
	.combout(\registerArray[13][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[13][26]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[13][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N9
dffeas \registerArray[13][26] (
	.clk(clk),
	.d(\registerArray[13][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][26] .is_wysiwyg = "true";
defparam \registerArray[13][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N21
dffeas \registerArray[12][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][26] .is_wysiwyg = "true";
defparam \registerArray[12][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N20
cycloneive_lcell_comb \Mux37~7 (
// Equation(s):
// \Mux37~7_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[13][26]~q )) # (!cuifregT_01 & ((\registerArray[12][26]~q )))))

	.dataa(cuifregT_1),
	.datab(\registerArray[13][26]~q ),
	.datac(\registerArray[12][26]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux37~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~7 .lut_mask = 16'hEE50;
defparam \Mux37~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N22
cycloneive_lcell_comb \Mux37~8 (
// Equation(s):
// \Mux37~8_combout  = (cuifregT_1 & ((\Mux37~7_combout  & ((\registerArray[15][26]~q ))) # (!\Mux37~7_combout  & (\registerArray[14][26]~q )))) # (!cuifregT_1 & (((\Mux37~7_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[14][26]~q ),
	.datac(\registerArray[15][26]~q ),
	.datad(\Mux37~7_combout ),
	.cin(gnd),
	.combout(\Mux37~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~8 .lut_mask = 16'hF588;
defparam \Mux37~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N15
dffeas \registerArray[6][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][26] .is_wysiwyg = "true";
defparam \registerArray[6][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N19
dffeas \registerArray[7][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][26] .is_wysiwyg = "true";
defparam \registerArray[7][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N26
cycloneive_lcell_comb \registerArray[5][26]~feeder (
// Equation(s):
// \registerArray[5][26]~feeder_combout  = \Mux42~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux422),
	.cin(gnd),
	.combout(\registerArray[5][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[5][26]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[5][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y31_N27
dffeas \registerArray[5][26] (
	.clk(clk),
	.d(\registerArray[5][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][26] .is_wysiwyg = "true";
defparam \registerArray[5][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N29
dffeas \registerArray[4][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][26] .is_wysiwyg = "true";
defparam \registerArray[4][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N28
cycloneive_lcell_comb \Mux37~2 (
// Equation(s):
// \Mux37~2_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[5][26]~q )) # (!cuifregT_01 & ((\registerArray[4][26]~q )))))

	.dataa(cuifregT_1),
	.datab(\registerArray[5][26]~q ),
	.datac(\registerArray[4][26]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux37~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~2 .lut_mask = 16'hEE50;
defparam \Mux37~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N18
cycloneive_lcell_comb \Mux37~3 (
// Equation(s):
// \Mux37~3_combout  = (cuifregT_1 & ((\Mux37~2_combout  & ((\registerArray[7][26]~q ))) # (!\Mux37~2_combout  & (\registerArray[6][26]~q )))) # (!cuifregT_1 & (((\Mux37~2_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[6][26]~q ),
	.datac(\registerArray[7][26]~q ),
	.datad(\Mux37~2_combout ),
	.cin(gnd),
	.combout(\Mux37~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~3 .lut_mask = 16'hF588;
defparam \Mux37~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y38_N3
dffeas \registerArray[2][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][26] .is_wysiwyg = "true";
defparam \registerArray[2][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y38_N29
dffeas \registerArray[1][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][26] .is_wysiwyg = "true";
defparam \registerArray[1][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N28
cycloneive_lcell_comb \Mux37~4 (
// Equation(s):
// \Mux37~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][26]~q )) # (!cuifregT_1 & ((\registerArray[1][26]~q )))))

	.dataa(\registerArray[3][26]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[1][26]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux37~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~4 .lut_mask = 16'h88C0;
defparam \Mux37~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N2
cycloneive_lcell_comb \Mux37~5 (
// Equation(s):
// \Mux37~5_combout  = (\Mux37~4_combout ) # ((cuifregT_1 & (!cuifregT_01 & \registerArray[2][26]~q )))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\registerArray[2][26]~q ),
	.datad(\Mux37~4_combout ),
	.cin(gnd),
	.combout(\Mux37~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~5 .lut_mask = 16'hFF20;
defparam \Mux37~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y34_N4
cycloneive_lcell_comb \Mux37~6 (
// Equation(s):
// \Mux37~6_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\Mux37~3_combout )) # (!cuifregT_2 & ((\Mux37~5_combout )))))

	.dataa(cuifregT_3),
	.datab(\Mux37~3_combout ),
	.datac(cuifregT_2),
	.datad(\Mux37~5_combout ),
	.cin(gnd),
	.combout(\Mux37~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~6 .lut_mask = 16'hE5E0;
defparam \Mux37~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N21
dffeas \registerArray[11][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][26] .is_wysiwyg = "true";
defparam \registerArray[11][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N31
dffeas \registerArray[9][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][26] .is_wysiwyg = "true";
defparam \registerArray[9][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N17
dffeas \registerArray[8][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][26] .is_wysiwyg = "true";
defparam \registerArray[8][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N15
dffeas \registerArray[10][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][26] .is_wysiwyg = "true";
defparam \registerArray[10][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N14
cycloneive_lcell_comb \Mux37~0 (
// Equation(s):
// \Mux37~0_combout  = (cuifregT_1 & (((\registerArray[10][26]~q ) # (cuifregT_01)))) # (!cuifregT_1 & (\registerArray[8][26]~q  & ((!cuifregT_01))))

	.dataa(cuifregT_1),
	.datab(\registerArray[8][26]~q ),
	.datac(\registerArray[10][26]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~0 .lut_mask = 16'hAAE4;
defparam \Mux37~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N30
cycloneive_lcell_comb \Mux37~1 (
// Equation(s):
// \Mux37~1_combout  = (cuifregT_01 & ((\Mux37~0_combout  & (\registerArray[11][26]~q )) # (!\Mux37~0_combout  & ((\registerArray[9][26]~q ))))) # (!cuifregT_01 & (((\Mux37~0_combout ))))

	.dataa(cuifregT_0),
	.datab(\registerArray[11][26]~q ),
	.datac(\registerArray[9][26]~q ),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\Mux37~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~1 .lut_mask = 16'hDDA0;
defparam \Mux37~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y41_N21
dffeas \registerArray[25][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][26] .is_wysiwyg = "true";
defparam \registerArray[25][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N23
dffeas \registerArray[29][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][26] .is_wysiwyg = "true";
defparam \registerArray[29][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y41_N19
dffeas \registerArray[21][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][26] .is_wysiwyg = "true";
defparam \registerArray[21][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N13
dffeas \registerArray[17][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][26] .is_wysiwyg = "true";
defparam \registerArray[17][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N12
cycloneive_lcell_comb \Mux37~10 (
// Equation(s):
// \Mux37~10_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[21][26]~q )) # (!cuifregT_2 & ((\registerArray[17][26]~q )))))

	.dataa(cuifregT_3),
	.datab(\registerArray[21][26]~q ),
	.datac(\registerArray[17][26]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux37~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~10 .lut_mask = 16'hEE50;
defparam \Mux37~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N22
cycloneive_lcell_comb \Mux37~11 (
// Equation(s):
// \Mux37~11_combout  = (cuifregT_3 & ((\Mux37~10_combout  & ((\registerArray[29][26]~q ))) # (!\Mux37~10_combout  & (\registerArray[25][26]~q )))) # (!cuifregT_3 & (((\Mux37~10_combout ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[25][26]~q ),
	.datac(\registerArray[29][26]~q ),
	.datad(\Mux37~10_combout ),
	.cin(gnd),
	.combout(\Mux37~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~11 .lut_mask = 16'hF588;
defparam \Mux37~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y31_N5
dffeas \registerArray[19][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][26] .is_wysiwyg = "true";
defparam \registerArray[19][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N18
cycloneive_lcell_comb \Mux37~17 (
// Equation(s):
// \Mux37~17_combout  = (cuifregT_2 & ((\registerArray[23][26]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[19][26]~q  & !cuifregT_3))))

	.dataa(\registerArray[23][26]~q ),
	.datab(\registerArray[19][26]~q ),
	.datac(cuifregT_2),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux37~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~17 .lut_mask = 16'hF0AC;
defparam \Mux37~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N3
dffeas \registerArray[31][26] (
	.clk(clk),
	.d(Mux422),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][26] .is_wysiwyg = "true";
defparam \registerArray[31][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N17
dffeas \registerArray[27][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][26] .is_wysiwyg = "true";
defparam \registerArray[27][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N16
cycloneive_lcell_comb \Mux37~18 (
// Equation(s):
// \Mux37~18_combout  = (\Mux37~17_combout  & ((\registerArray[31][26]~q ) # ((!cuifregT_3)))) # (!\Mux37~17_combout  & (((\registerArray[27][26]~q  & cuifregT_3))))

	.dataa(\Mux37~17_combout ),
	.datab(\registerArray[31][26]~q ),
	.datac(\registerArray[27][26]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux37~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~18 .lut_mask = 16'hD8AA;
defparam \Mux37~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y35_N23
dffeas \registerArray[28][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][26] .is_wysiwyg = "true";
defparam \registerArray[28][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N8
cycloneive_lcell_comb \registerArray[24][26]~feeder (
// Equation(s):
// \registerArray[24][26]~feeder_combout  = \Mux42~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux422),
	.cin(gnd),
	.combout(\registerArray[24][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[24][26]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[24][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N9
dffeas \registerArray[24][26] (
	.clk(clk),
	.d(\registerArray[24][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][26] .is_wysiwyg = "true";
defparam \registerArray[24][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y35_N1
dffeas \registerArray[16][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][26] .is_wysiwyg = "true";
defparam \registerArray[16][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N0
cycloneive_lcell_comb \Mux37~14 (
// Equation(s):
// \Mux37~14_combout  = (cuifregT_3 & ((\registerArray[24][26]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[16][26]~q  & !cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[24][26]~q ),
	.datac(\registerArray[16][26]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux37~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~14 .lut_mask = 16'hAAD8;
defparam \Mux37~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N22
cycloneive_lcell_comb \Mux37~15 (
// Equation(s):
// \Mux37~15_combout  = (cuifregT_2 & ((\Mux37~14_combout  & ((\registerArray[28][26]~q ))) # (!\Mux37~14_combout  & (\registerArray[20][26]~q )))) # (!cuifregT_2 & (((\Mux37~14_combout ))))

	.dataa(\registerArray[20][26]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[28][26]~q ),
	.datad(\Mux37~14_combout ),
	.cin(gnd),
	.combout(\Mux37~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~15 .lut_mask = 16'hF388;
defparam \Mux37~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N17
dffeas \registerArray[22][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][26] .is_wysiwyg = "true";
defparam \registerArray[22][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N3
dffeas \registerArray[30][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][26] .is_wysiwyg = "true";
defparam \registerArray[30][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N7
dffeas \registerArray[26][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][26] .is_wysiwyg = "true";
defparam \registerArray[26][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N21
dffeas \registerArray[18][26] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux422),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][26] .is_wysiwyg = "true";
defparam \registerArray[18][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N20
cycloneive_lcell_comb \Mux37~12 (
// Equation(s):
// \Mux37~12_combout  = (cuifregT_3 & ((\registerArray[26][26]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[18][26]~q  & !cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[26][26]~q ),
	.datac(\registerArray[18][26]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux37~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~12 .lut_mask = 16'hAAD8;
defparam \Mux37~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N2
cycloneive_lcell_comb \Mux37~13 (
// Equation(s):
// \Mux37~13_combout  = (cuifregT_2 & ((\Mux37~12_combout  & ((\registerArray[30][26]~q ))) # (!\Mux37~12_combout  & (\registerArray[22][26]~q )))) # (!cuifregT_2 & (((\Mux37~12_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[22][26]~q ),
	.datac(\registerArray[30][26]~q ),
	.datad(\Mux37~12_combout ),
	.cin(gnd),
	.combout(\Mux37~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~13 .lut_mask = 16'hF588;
defparam \Mux37~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y35_N28
cycloneive_lcell_comb \Mux37~16 (
// Equation(s):
// \Mux37~16_combout  = (cuifregT_01 & (cuifregT_1)) # (!cuifregT_01 & ((cuifregT_1 & ((\Mux37~13_combout ))) # (!cuifregT_1 & (\Mux37~15_combout ))))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\Mux37~15_combout ),
	.datad(\Mux37~13_combout ),
	.cin(gnd),
	.combout(\Mux37~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~16 .lut_mask = 16'hDC98;
defparam \Mux37~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N23
dffeas \registerArray[14][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][25] .is_wysiwyg = "true";
defparam \registerArray[14][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N29
dffeas \registerArray[12][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][25] .is_wysiwyg = "true";
defparam \registerArray[12][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N3
dffeas \registerArray[13][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][25] .is_wysiwyg = "true";
defparam \registerArray[13][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N28
cycloneive_lcell_comb \Mux38~7 (
// Equation(s):
// \Mux38~7_combout  = (cuifregT_01 & ((cuifregT_1) # ((\registerArray[13][25]~q )))) # (!cuifregT_01 & (!cuifregT_1 & (\registerArray[12][25]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[12][25]~q ),
	.datad(\registerArray[13][25]~q ),
	.cin(gnd),
	.combout(\Mux38~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~7 .lut_mask = 16'hBA98;
defparam \Mux38~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y38_N3
dffeas \registerArray[15][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][25] .is_wysiwyg = "true";
defparam \registerArray[15][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N2
cycloneive_lcell_comb \Mux38~8 (
// Equation(s):
// \Mux38~8_combout  = (\Mux38~7_combout  & (((\registerArray[15][25]~q ) # (!cuifregT_1)))) # (!\Mux38~7_combout  & (\registerArray[14][25]~q  & ((cuifregT_1))))

	.dataa(\registerArray[14][25]~q ),
	.datab(\Mux38~7_combout ),
	.datac(\registerArray[15][25]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux38~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~8 .lut_mask = 16'hE2CC;
defparam \Mux38~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N1
dffeas \registerArray[6][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][25] .is_wysiwyg = "true";
defparam \registerArray[6][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N15
dffeas \registerArray[7][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][25] .is_wysiwyg = "true";
defparam \registerArray[7][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N26
cycloneive_lcell_comb \registerArray[5][25]~feeder (
// Equation(s):
// \registerArray[5][25]~feeder_combout  = \Mux43~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux432),
	.cin(gnd),
	.combout(\registerArray[5][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[5][25]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[5][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N27
dffeas \registerArray[5][25] (
	.clk(clk),
	.d(\registerArray[5][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][25] .is_wysiwyg = "true";
defparam \registerArray[5][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y32_N17
dffeas \registerArray[4][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][25] .is_wysiwyg = "true";
defparam \registerArray[4][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N16
cycloneive_lcell_comb \Mux38~0 (
// Equation(s):
// \Mux38~0_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[5][25]~q )) # (!cuifregT_01 & ((\registerArray[4][25]~q )))))

	.dataa(cuifregT_1),
	.datab(\registerArray[5][25]~q ),
	.datac(\registerArray[4][25]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux38~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~0 .lut_mask = 16'hEE50;
defparam \Mux38~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N14
cycloneive_lcell_comb \Mux38~1 (
// Equation(s):
// \Mux38~1_combout  = (cuifregT_1 & ((\Mux38~0_combout  & ((\registerArray[7][25]~q ))) # (!\Mux38~0_combout  & (\registerArray[6][25]~q )))) # (!cuifregT_1 & (((\Mux38~0_combout ))))

	.dataa(\registerArray[6][25]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[7][25]~q ),
	.datad(\Mux38~0_combout ),
	.cin(gnd),
	.combout(\Mux38~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~1 .lut_mask = 16'hF388;
defparam \Mux38~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N7
dffeas \registerArray[11][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][25] .is_wysiwyg = "true";
defparam \registerArray[11][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N21
dffeas \registerArray[8][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][25] .is_wysiwyg = "true";
defparam \registerArray[8][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N20
cycloneive_lcell_comb \Mux38~2 (
// Equation(s):
// \Mux38~2_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & (\registerArray[10][25]~q )) # (!cuifregT_1 & ((\registerArray[8][25]~q )))))

	.dataa(\registerArray[10][25]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[8][25]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux38~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~2 .lut_mask = 16'hEE30;
defparam \Mux38~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N6
cycloneive_lcell_comb \Mux38~3 (
// Equation(s):
// \Mux38~3_combout  = (cuifregT_01 & ((\Mux38~2_combout  & ((\registerArray[11][25]~q ))) # (!\Mux38~2_combout  & (\registerArray[9][25]~q )))) # (!cuifregT_01 & (((\Mux38~2_combout ))))

	.dataa(\registerArray[9][25]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[11][25]~q ),
	.datad(\Mux38~2_combout ),
	.cin(gnd),
	.combout(\Mux38~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~3 .lut_mask = 16'hF388;
defparam \Mux38~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y41_N7
dffeas \registerArray[2][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][25] .is_wysiwyg = "true";
defparam \registerArray[2][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N25
dffeas \registerArray[3][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][25] .is_wysiwyg = "true";
defparam \registerArray[3][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y41_N25
dffeas \registerArray[1][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][25] .is_wysiwyg = "true";
defparam \registerArray[1][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N24
cycloneive_lcell_comb \Mux38~4 (
// Equation(s):
// \Mux38~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][25]~q )) # (!cuifregT_1 & ((\registerArray[1][25]~q )))))

	.dataa(cuifregT_0),
	.datab(\registerArray[3][25]~q ),
	.datac(\registerArray[1][25]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux38~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~4 .lut_mask = 16'h88A0;
defparam \Mux38~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N6
cycloneive_lcell_comb \Mux38~5 (
// Equation(s):
// \Mux38~5_combout  = (\Mux38~4_combout ) # ((!cuifregT_01 & (cuifregT_1 & \registerArray[2][25]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[2][25]~q ),
	.datad(\Mux38~4_combout ),
	.cin(gnd),
	.combout(\Mux38~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~5 .lut_mask = 16'hFF40;
defparam \Mux38~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N20
cycloneive_lcell_comb \Mux38~6 (
// Equation(s):
// \Mux38~6_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\Mux38~3_combout )) # (!cuifregT_3 & ((\Mux38~5_combout )))))

	.dataa(\Mux38~3_combout ),
	.datab(cuifregT_2),
	.datac(cuifregT_3),
	.datad(\Mux38~5_combout ),
	.cin(gnd),
	.combout(\Mux38~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~6 .lut_mask = 16'hE3E0;
defparam \Mux38~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N27
dffeas \registerArray[30][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][25] .is_wysiwyg = "true";
defparam \registerArray[30][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N5
dffeas \registerArray[18][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][25] .is_wysiwyg = "true";
defparam \registerArray[18][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N4
cycloneive_lcell_comb \Mux38~12 (
// Equation(s):
// \Mux38~12_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[22][25]~q )) # (!cuifregT_2 & ((\registerArray[18][25]~q )))))

	.dataa(\registerArray[22][25]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[18][25]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux38~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~12 .lut_mask = 16'hEE30;
defparam \Mux38~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N26
cycloneive_lcell_comb \Mux38~13 (
// Equation(s):
// \Mux38~13_combout  = (cuifregT_3 & ((\Mux38~12_combout  & ((\registerArray[30][25]~q ))) # (!\Mux38~12_combout  & (\registerArray[26][25]~q )))) # (!cuifregT_3 & (((\Mux38~12_combout ))))

	.dataa(\registerArray[26][25]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[30][25]~q ),
	.datad(\Mux38~12_combout ),
	.cin(gnd),
	.combout(\Mux38~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~13 .lut_mask = 16'hF388;
defparam \Mux38~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y30_N7
dffeas \registerArray[28][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][25] .is_wysiwyg = "true";
defparam \registerArray[28][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N15
dffeas \registerArray[20][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][25] .is_wysiwyg = "true";
defparam \registerArray[20][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N25
dffeas \registerArray[16][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][25] .is_wysiwyg = "true";
defparam \registerArray[16][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N24
cycloneive_lcell_comb \Mux38~14 (
// Equation(s):
// \Mux38~14_combout  = (cuifregT_2 & ((\registerArray[20][25]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[16][25]~q  & !cuifregT_3))))

	.dataa(cuifregT_2),
	.datab(\registerArray[20][25]~q ),
	.datac(\registerArray[16][25]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux38~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~14 .lut_mask = 16'hAAD8;
defparam \Mux38~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N6
cycloneive_lcell_comb \Mux38~15 (
// Equation(s):
// \Mux38~15_combout  = (cuifregT_3 & ((\Mux38~14_combout  & ((\registerArray[28][25]~q ))) # (!\Mux38~14_combout  & (\registerArray[24][25]~q )))) # (!cuifregT_3 & (((\Mux38~14_combout ))))

	.dataa(\registerArray[24][25]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[28][25]~q ),
	.datad(\Mux38~14_combout ),
	.cin(gnd),
	.combout(\Mux38~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~15 .lut_mask = 16'hF388;
defparam \Mux38~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N0
cycloneive_lcell_comb \Mux38~16 (
// Equation(s):
// \Mux38~16_combout  = (cuifregT_1 & ((cuifregT_01) # ((\Mux38~13_combout )))) # (!cuifregT_1 & (!cuifregT_01 & ((\Mux38~15_combout ))))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\Mux38~13_combout ),
	.datad(\Mux38~15_combout ),
	.cin(gnd),
	.combout(\Mux38~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~16 .lut_mask = 16'hB9A8;
defparam \Mux38~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y41_N25
dffeas \registerArray[23][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][25] .is_wysiwyg = "true";
defparam \registerArray[23][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y41_N25
dffeas \registerArray[31][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][25] .is_wysiwyg = "true";
defparam \registerArray[31][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N7
dffeas \registerArray[19][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][25] .is_wysiwyg = "true";
defparam \registerArray[19][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N6
cycloneive_lcell_comb \Mux38~17 (
// Equation(s):
// \Mux38~17_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[27][25]~q )) # (!cuifregT_3 & ((\registerArray[19][25]~q )))))

	.dataa(\registerArray[27][25]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[19][25]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux38~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~17 .lut_mask = 16'hEE30;
defparam \Mux38~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N24
cycloneive_lcell_comb \Mux38~18 (
// Equation(s):
// \Mux38~18_combout  = (cuifregT_2 & ((\Mux38~17_combout  & ((\registerArray[31][25]~q ))) # (!\Mux38~17_combout  & (\registerArray[23][25]~q )))) # (!cuifregT_2 & (((\Mux38~17_combout ))))

	.dataa(\registerArray[23][25]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[31][25]~q ),
	.datad(\Mux38~17_combout ),
	.cin(gnd),
	.combout(\Mux38~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~18 .lut_mask = 16'hF388;
defparam \Mux38~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y30_N23
dffeas \registerArray[21][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][25] .is_wysiwyg = "true";
defparam \registerArray[21][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N7
dffeas \registerArray[29][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][25] .is_wysiwyg = "true";
defparam \registerArray[29][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N25
dffeas \registerArray[25][25] (
	.clk(clk),
	.d(Mux432),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][25] .is_wysiwyg = "true";
defparam \registerArray[25][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N17
dffeas \registerArray[17][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][25] .is_wysiwyg = "true";
defparam \registerArray[17][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N16
cycloneive_lcell_comb \Mux38~10 (
// Equation(s):
// \Mux38~10_combout  = (cuifregT_3 & ((\registerArray[25][25]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[17][25]~q  & !cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[25][25]~q ),
	.datac(\registerArray[17][25]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux38~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~10 .lut_mask = 16'hAAD8;
defparam \Mux38~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N6
cycloneive_lcell_comb \Mux38~11 (
// Equation(s):
// \Mux38~11_combout  = (cuifregT_2 & ((\Mux38~10_combout  & ((\registerArray[29][25]~q ))) # (!\Mux38~10_combout  & (\registerArray[21][25]~q )))) # (!cuifregT_2 & (((\Mux38~10_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[21][25]~q ),
	.datac(\registerArray[29][25]~q ),
	.datad(\Mux38~10_combout ),
	.cin(gnd),
	.combout(\Mux38~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~11 .lut_mask = 16'hF588;
defparam \Mux38~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N0
cycloneive_lcell_comb \registerArray[29][24]~feeder (
// Equation(s):
// \registerArray[29][24]~feeder_combout  = \Mux44~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux442),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[29][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[29][24]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[29][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N1
dffeas \registerArray[29][24] (
	.clk(clk),
	.d(\registerArray[29][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][24] .is_wysiwyg = "true";
defparam \registerArray[29][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N4
cycloneive_lcell_comb \registerArray[25][24]~feeder (
// Equation(s):
// \registerArray[25][24]~feeder_combout  = \Mux44~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux442),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[25][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[25][24]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[25][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N5
dffeas \registerArray[25][24] (
	.clk(clk),
	.d(\registerArray[25][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][24] .is_wysiwyg = "true";
defparam \registerArray[25][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N4
cycloneive_lcell_comb \registerArray[17][24]~feeder (
// Equation(s):
// \registerArray[17][24]~feeder_combout  = \Mux44~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux442),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[17][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[17][24]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[17][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N5
dffeas \registerArray[17][24] (
	.clk(clk),
	.d(\registerArray[17][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][24] .is_wysiwyg = "true";
defparam \registerArray[17][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N16
cycloneive_lcell_comb \registerArray[21][24]~feeder (
// Equation(s):
// \registerArray[21][24]~feeder_combout  = \Mux44~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux442),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[21][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[21][24]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[21][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N17
dffeas \registerArray[21][24] (
	.clk(clk),
	.d(\registerArray[21][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][24] .is_wysiwyg = "true";
defparam \registerArray[21][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N6
cycloneive_lcell_comb \Mux39~0 (
// Equation(s):
// \Mux39~0_combout  = (cuifregT_2 & (((cuifregT_3) # (\registerArray[21][24]~q )))) # (!cuifregT_2 & (\registerArray[17][24]~q  & (!cuifregT_3)))

	.dataa(cuifregT_2),
	.datab(\registerArray[17][24]~q ),
	.datac(cuifregT_3),
	.datad(\registerArray[21][24]~q ),
	.cin(gnd),
	.combout(\Mux39~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~0 .lut_mask = 16'hAEA4;
defparam \Mux39~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N22
cycloneive_lcell_comb \Mux39~1 (
// Equation(s):
// \Mux39~1_combout  = (cuifregT_3 & ((\Mux39~0_combout  & (\registerArray[29][24]~q )) # (!\Mux39~0_combout  & ((\registerArray[25][24]~q ))))) # (!cuifregT_3 & (((\Mux39~0_combout ))))

	.dataa(\registerArray[29][24]~q ),
	.datab(\registerArray[25][24]~q ),
	.datac(cuifregT_3),
	.datad(\Mux39~0_combout ),
	.cin(gnd),
	.combout(\Mux39~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~1 .lut_mask = 16'hAFC0;
defparam \Mux39~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N13
dffeas \registerArray[27][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][24] .is_wysiwyg = "true";
defparam \registerArray[27][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N7
dffeas \registerArray[31][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][24] .is_wysiwyg = "true";
defparam \registerArray[31][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N23
dffeas \registerArray[19][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][24] .is_wysiwyg = "true";
defparam \registerArray[19][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N22
cycloneive_lcell_comb \Mux39~7 (
// Equation(s):
// \Mux39~7_combout  = (cuifregT_2 & ((\registerArray[23][24]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[19][24]~q  & !cuifregT_3))))

	.dataa(\registerArray[23][24]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[19][24]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux39~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~7 .lut_mask = 16'hCCB8;
defparam \Mux39~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N6
cycloneive_lcell_comb \Mux39~8 (
// Equation(s):
// \Mux39~8_combout  = (cuifregT_3 & ((\Mux39~7_combout  & ((\registerArray[31][24]~q ))) # (!\Mux39~7_combout  & (\registerArray[27][24]~q )))) # (!cuifregT_3 & (((\Mux39~7_combout ))))

	.dataa(\registerArray[27][24]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[31][24]~q ),
	.datad(\Mux39~7_combout ),
	.cin(gnd),
	.combout(\Mux39~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~8 .lut_mask = 16'hF388;
defparam \Mux39~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N30
cycloneive_lcell_comb \registerArray[28][24]~feeder (
// Equation(s):
// \registerArray[28][24]~feeder_combout  = \Mux44~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux442),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[28][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[28][24]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[28][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N31
dffeas \registerArray[28][24] (
	.clk(clk),
	.d(\registerArray[28][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][24] .is_wysiwyg = "true";
defparam \registerArray[28][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N30
cycloneive_lcell_comb \registerArray[24][24]~feeder (
// Equation(s):
// \registerArray[24][24]~feeder_combout  = \Mux44~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux442),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[24][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[24][24]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[24][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N31
dffeas \registerArray[24][24] (
	.clk(clk),
	.d(\registerArray[24][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][24] .is_wysiwyg = "true";
defparam \registerArray[24][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N0
cycloneive_lcell_comb \Mux39~4 (
// Equation(s):
// \Mux39~4_combout  = (cuifregT_3 & (((cuifregT_2) # (\registerArray[24][24]~q )))) # (!cuifregT_3 & (\registerArray[16][24]~q  & (!cuifregT_2)))

	.dataa(\registerArray[16][24]~q ),
	.datab(cuifregT_3),
	.datac(cuifregT_2),
	.datad(\registerArray[24][24]~q ),
	.cin(gnd),
	.combout(\Mux39~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~4 .lut_mask = 16'hCEC2;
defparam \Mux39~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N12
cycloneive_lcell_comb \Mux39~5 (
// Equation(s):
// \Mux39~5_combout  = (cuifregT_2 & ((\Mux39~4_combout  & ((\registerArray[28][24]~q ))) # (!\Mux39~4_combout  & (\registerArray[20][24]~q )))) # (!cuifregT_2 & (((\Mux39~4_combout ))))

	.dataa(\registerArray[20][24]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[28][24]~q ),
	.datad(\Mux39~4_combout ),
	.cin(gnd),
	.combout(\Mux39~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~5 .lut_mask = 16'hF388;
defparam \Mux39~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N9
dffeas \registerArray[22][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][24] .is_wysiwyg = "true";
defparam \registerArray[22][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N7
dffeas \registerArray[30][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][24] .is_wysiwyg = "true";
defparam \registerArray[30][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N25
dffeas \registerArray[18][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][24] .is_wysiwyg = "true";
defparam \registerArray[18][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N24
cycloneive_lcell_comb \Mux39~2 (
// Equation(s):
// \Mux39~2_combout  = (cuifregT_3 & ((\registerArray[26][24]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[18][24]~q  & !cuifregT_2))))

	.dataa(\registerArray[26][24]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[18][24]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux39~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~2 .lut_mask = 16'hCCB8;
defparam \Mux39~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N6
cycloneive_lcell_comb \Mux39~3 (
// Equation(s):
// \Mux39~3_combout  = (cuifregT_2 & ((\Mux39~2_combout  & ((\registerArray[30][24]~q ))) # (!\Mux39~2_combout  & (\registerArray[22][24]~q )))) # (!cuifregT_2 & (((\Mux39~2_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[22][24]~q ),
	.datac(\registerArray[30][24]~q ),
	.datad(\Mux39~2_combout ),
	.cin(gnd),
	.combout(\Mux39~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~3 .lut_mask = 16'hF588;
defparam \Mux39~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N6
cycloneive_lcell_comb \Mux39~6 (
// Equation(s):
// \Mux39~6_combout  = (cuifregT_1 & (((cuifregT_01) # (\Mux39~3_combout )))) # (!cuifregT_1 & (\Mux39~5_combout  & (!cuifregT_01)))

	.dataa(\Mux39~5_combout ),
	.datab(cuifregT_1),
	.datac(cuifregT_0),
	.datad(\Mux39~3_combout ),
	.cin(gnd),
	.combout(\Mux39~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~6 .lut_mask = 16'hCEC2;
defparam \Mux39~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N30
cycloneive_lcell_comb \registerArray[14][24]~feeder (
// Equation(s):
// \registerArray[14][24]~feeder_combout  = \Mux44~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux442),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[14][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][24]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[14][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N31
dffeas \registerArray[14][24] (
	.clk(clk),
	.d(\registerArray[14][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][24] .is_wysiwyg = "true";
defparam \registerArray[14][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N31
dffeas \registerArray[15][24] (
	.clk(clk),
	.d(Mux442),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][24] .is_wysiwyg = "true";
defparam \registerArray[15][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N25
dffeas \registerArray[13][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][24] .is_wysiwyg = "true";
defparam \registerArray[13][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N28
cycloneive_lcell_comb \Mux39~17 (
// Equation(s):
// \Mux39~17_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & ((\registerArray[13][24]~q ))) # (!cuifregT_01 & (\registerArray[12][24]~q ))))

	.dataa(\registerArray[12][24]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[13][24]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux39~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~17 .lut_mask = 16'hFC22;
defparam \Mux39~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N18
cycloneive_lcell_comb \Mux39~18 (
// Equation(s):
// \Mux39~18_combout  = (cuifregT_1 & ((\Mux39~17_combout  & ((\registerArray[15][24]~q ))) # (!\Mux39~17_combout  & (\registerArray[14][24]~q )))) # (!cuifregT_1 & (((\Mux39~17_combout ))))

	.dataa(\registerArray[14][24]~q ),
	.datab(\registerArray[15][24]~q ),
	.datac(cuifregT_1),
	.datad(\Mux39~17_combout ),
	.cin(gnd),
	.combout(\Mux39~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~18 .lut_mask = 16'hCFA0;
defparam \Mux39~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y43_N25
dffeas \registerArray[9][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][24] .is_wysiwyg = "true";
defparam \registerArray[9][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N31
dffeas \registerArray[11][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][24] .is_wysiwyg = "true";
defparam \registerArray[11][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N1
dffeas \registerArray[8][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][24] .is_wysiwyg = "true";
defparam \registerArray[8][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N0
cycloneive_lcell_comb \Mux39~10 (
// Equation(s):
// \Mux39~10_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & (\registerArray[10][24]~q )) # (!cuifregT_1 & ((\registerArray[8][24]~q )))))

	.dataa(\registerArray[10][24]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[8][24]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux39~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~10 .lut_mask = 16'hEE30;
defparam \Mux39~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N30
cycloneive_lcell_comb \Mux39~11 (
// Equation(s):
// \Mux39~11_combout  = (cuifregT_01 & ((\Mux39~10_combout  & ((\registerArray[11][24]~q ))) # (!\Mux39~10_combout  & (\registerArray[9][24]~q )))) # (!cuifregT_01 & (((\Mux39~10_combout ))))

	.dataa(\registerArray[9][24]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[11][24]~q ),
	.datad(\Mux39~10_combout ),
	.cin(gnd),
	.combout(\Mux39~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~11 .lut_mask = 16'hF388;
defparam \Mux39~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y42_N21
dffeas \registerArray[6][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][24] .is_wysiwyg = "true";
defparam \registerArray[6][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N23
dffeas \registerArray[4][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][24] .is_wysiwyg = "true";
defparam \registerArray[4][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N22
cycloneive_lcell_comb \Mux39~12 (
// Equation(s):
// \Mux39~12_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[5][24]~q )) # (!cuifregT_01 & ((\registerArray[4][24]~q )))))

	.dataa(\registerArray[5][24]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[4][24]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux39~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~12 .lut_mask = 16'hEE30;
defparam \Mux39~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N6
cycloneive_lcell_comb \Mux39~13 (
// Equation(s):
// \Mux39~13_combout  = (cuifregT_1 & ((\Mux39~12_combout  & (\registerArray[7][24]~q )) # (!\Mux39~12_combout  & ((\registerArray[6][24]~q ))))) # (!cuifregT_1 & (((\Mux39~12_combout ))))

	.dataa(\registerArray[7][24]~q ),
	.datab(\registerArray[6][24]~q ),
	.datac(cuifregT_1),
	.datad(\Mux39~12_combout ),
	.cin(gnd),
	.combout(\Mux39~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~13 .lut_mask = 16'hAFC0;
defparam \Mux39~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N15
dffeas \registerArray[2][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][24] .is_wysiwyg = "true";
defparam \registerArray[2][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y37_N25
dffeas \registerArray[1][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][24] .is_wysiwyg = "true";
defparam \registerArray[1][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N24
cycloneive_lcell_comb \Mux39~14 (
// Equation(s):
// \Mux39~14_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][24]~q )) # (!cuifregT_1 & ((\registerArray[1][24]~q )))))

	.dataa(\registerArray[3][24]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[1][24]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux39~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~14 .lut_mask = 16'h88C0;
defparam \Mux39~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N14
cycloneive_lcell_comb \Mux39~15 (
// Equation(s):
// \Mux39~15_combout  = (\Mux39~14_combout ) # ((cuifregT_1 & (!cuifregT_01 & \registerArray[2][24]~q )))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\registerArray[2][24]~q ),
	.datad(\Mux39~14_combout ),
	.cin(gnd),
	.combout(\Mux39~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~15 .lut_mask = 16'hFF20;
defparam \Mux39~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N24
cycloneive_lcell_comb \Mux39~16 (
// Equation(s):
// \Mux39~16_combout  = (cuifregT_2 & ((\Mux39~13_combout ) # ((cuifregT_3)))) # (!cuifregT_2 & (((!cuifregT_3 & \Mux39~15_combout ))))

	.dataa(\Mux39~13_combout ),
	.datab(cuifregT_2),
	.datac(cuifregT_3),
	.datad(\Mux39~15_combout ),
	.cin(gnd),
	.combout(\Mux39~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~16 .lut_mask = 16'hCBC8;
defparam \Mux39~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N28
cycloneive_lcell_comb \registerArray[14][23]~feeder (
// Equation(s):
// \registerArray[14][23]~feeder_combout  = \Mux45~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux452),
	.cin(gnd),
	.combout(\registerArray[14][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][23]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[14][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N29
dffeas \registerArray[14][23] (
	.clk(clk),
	.d(\registerArray[14][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][23] .is_wysiwyg = "true";
defparam \registerArray[14][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N19
dffeas \registerArray[15][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][23] .is_wysiwyg = "true";
defparam \registerArray[15][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N1
dffeas \registerArray[12][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][23] .is_wysiwyg = "true";
defparam \registerArray[12][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N30
cycloneive_lcell_comb \registerArray[13][23]~feeder (
// Equation(s):
// \registerArray[13][23]~feeder_combout  = \Mux45~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux452),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[13][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[13][23]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[13][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N31
dffeas \registerArray[13][23] (
	.clk(clk),
	.d(\registerArray[13][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][23] .is_wysiwyg = "true";
defparam \registerArray[13][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N0
cycloneive_lcell_comb \Mux40~7 (
// Equation(s):
// \Mux40~7_combout  = (cuifregT_01 & ((cuifregT_1) # ((\registerArray[13][23]~q )))) # (!cuifregT_01 & (!cuifregT_1 & (\registerArray[12][23]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[12][23]~q ),
	.datad(\registerArray[13][23]~q ),
	.cin(gnd),
	.combout(\Mux40~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~7 .lut_mask = 16'hBA98;
defparam \Mux40~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N18
cycloneive_lcell_comb \Mux40~8 (
// Equation(s):
// \Mux40~8_combout  = (cuifregT_1 & ((\Mux40~7_combout  & ((\registerArray[15][23]~q ))) # (!\Mux40~7_combout  & (\registerArray[14][23]~q )))) # (!cuifregT_1 & (((\Mux40~7_combout ))))

	.dataa(\registerArray[14][23]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[15][23]~q ),
	.datad(\Mux40~7_combout ),
	.cin(gnd),
	.combout(\Mux40~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~8 .lut_mask = 16'hF388;
defparam \Mux40~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N11
dffeas \registerArray[6][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][23] .is_wysiwyg = "true";
defparam \registerArray[6][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N17
dffeas \registerArray[7][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][23] .is_wysiwyg = "true";
defparam \registerArray[7][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N31
dffeas \registerArray[4][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][23] .is_wysiwyg = "true";
defparam \registerArray[4][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N30
cycloneive_lcell_comb \Mux40~0 (
// Equation(s):
// \Mux40~0_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[5][23]~q )) # (!cuifregT_01 & ((\registerArray[4][23]~q )))))

	.dataa(\registerArray[5][23]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[4][23]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux40~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~0 .lut_mask = 16'hEE30;
defparam \Mux40~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N16
cycloneive_lcell_comb \Mux40~1 (
// Equation(s):
// \Mux40~1_combout  = (cuifregT_1 & ((\Mux40~0_combout  & ((\registerArray[7][23]~q ))) # (!\Mux40~0_combout  & (\registerArray[6][23]~q )))) # (!cuifregT_1 & (((\Mux40~0_combout ))))

	.dataa(\registerArray[6][23]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[7][23]~q ),
	.datad(\Mux40~0_combout ),
	.cin(gnd),
	.combout(\Mux40~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~1 .lut_mask = 16'hF388;
defparam \Mux40~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y41_N23
dffeas \registerArray[2][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][23] .is_wysiwyg = "true";
defparam \registerArray[2][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N25
dffeas \registerArray[1][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][23] .is_wysiwyg = "true";
defparam \registerArray[1][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N24
cycloneive_lcell_comb \Mux40~4 (
// Equation(s):
// \Mux40~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][23]~q )) # (!cuifregT_1 & ((\registerArray[1][23]~q )))))

	.dataa(\registerArray[3][23]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[1][23]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux40~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~4 .lut_mask = 16'h88C0;
defparam \Mux40~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N22
cycloneive_lcell_comb \Mux40~5 (
// Equation(s):
// \Mux40~5_combout  = (\Mux40~4_combout ) # ((cuifregT_1 & (!cuifregT_01 & \registerArray[2][23]~q )))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\registerArray[2][23]~q ),
	.datad(\Mux40~4_combout ),
	.cin(gnd),
	.combout(\Mux40~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~5 .lut_mask = 16'hFF20;
defparam \Mux40~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y43_N29
dffeas \registerArray[9][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][23] .is_wysiwyg = "true";
defparam \registerArray[9][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N7
dffeas \registerArray[11][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][23] .is_wysiwyg = "true";
defparam \registerArray[11][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N29
dffeas \registerArray[8][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][23] .is_wysiwyg = "true";
defparam \registerArray[8][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N28
cycloneive_lcell_comb \Mux40~2 (
// Equation(s):
// \Mux40~2_combout  = (cuifregT_1 & ((\registerArray[10][23]~q ) # ((cuifregT_01)))) # (!cuifregT_1 & (((\registerArray[8][23]~q  & !cuifregT_01))))

	.dataa(\registerArray[10][23]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[8][23]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux40~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~2 .lut_mask = 16'hCCB8;
defparam \Mux40~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N6
cycloneive_lcell_comb \Mux40~3 (
// Equation(s):
// \Mux40~3_combout  = (cuifregT_01 & ((\Mux40~2_combout  & ((\registerArray[11][23]~q ))) # (!\Mux40~2_combout  & (\registerArray[9][23]~q )))) # (!cuifregT_01 & (((\Mux40~2_combout ))))

	.dataa(cuifregT_0),
	.datab(\registerArray[9][23]~q ),
	.datac(\registerArray[11][23]~q ),
	.datad(\Mux40~2_combout ),
	.cin(gnd),
	.combout(\Mux40~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~3 .lut_mask = 16'hF588;
defparam \Mux40~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N0
cycloneive_lcell_comb \Mux40~6 (
// Equation(s):
// \Mux40~6_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & ((\Mux40~3_combout ))) # (!cuifregT_3 & (\Mux40~5_combout ))))

	.dataa(\Mux40~5_combout ),
	.datab(cuifregT_2),
	.datac(cuifregT_3),
	.datad(\Mux40~3_combout ),
	.cin(gnd),
	.combout(\Mux40~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~6 .lut_mask = 16'hF2C2;
defparam \Mux40~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N11
dffeas \registerArray[22][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][23] .is_wysiwyg = "true";
defparam \registerArray[22][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N9
dffeas \registerArray[18][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][23] .is_wysiwyg = "true";
defparam \registerArray[18][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N8
cycloneive_lcell_comb \Mux40~12 (
// Equation(s):
// \Mux40~12_combout  = (cuifregT_2 & ((\registerArray[22][23]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[18][23]~q  & !cuifregT_3))))

	.dataa(cuifregT_2),
	.datab(\registerArray[22][23]~q ),
	.datac(\registerArray[18][23]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux40~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~12 .lut_mask = 16'hAAD8;
defparam \Mux40~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N15
dffeas \registerArray[30][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][23] .is_wysiwyg = "true";
defparam \registerArray[30][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N14
cycloneive_lcell_comb \Mux40~13 (
// Equation(s):
// \Mux40~13_combout  = (\Mux40~12_combout  & (((\registerArray[30][23]~q ) # (!cuifregT_3)))) # (!\Mux40~12_combout  & (\registerArray[26][23]~q  & ((cuifregT_3))))

	.dataa(\registerArray[26][23]~q ),
	.datab(\Mux40~12_combout ),
	.datac(\registerArray[30][23]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux40~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~13 .lut_mask = 16'hE2CC;
defparam \Mux40~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N3
dffeas \registerArray[28][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][23] .is_wysiwyg = "true";
defparam \registerArray[28][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y34_N17
dffeas \registerArray[16][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][23] .is_wysiwyg = "true";
defparam \registerArray[16][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N16
cycloneive_lcell_comb \Mux40~14 (
// Equation(s):
// \Mux40~14_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[20][23]~q )) # (!cuifregT_2 & ((\registerArray[16][23]~q )))))

	.dataa(\registerArray[20][23]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[16][23]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux40~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~14 .lut_mask = 16'hEE30;
defparam \Mux40~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N2
cycloneive_lcell_comb \Mux40~15 (
// Equation(s):
// \Mux40~15_combout  = (cuifregT_3 & ((\Mux40~14_combout  & ((\registerArray[28][23]~q ))) # (!\Mux40~14_combout  & (\registerArray[24][23]~q )))) # (!cuifregT_3 & (((\Mux40~14_combout ))))

	.dataa(\registerArray[24][23]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[28][23]~q ),
	.datad(\Mux40~14_combout ),
	.cin(gnd),
	.combout(\Mux40~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~15 .lut_mask = 16'hF388;
defparam \Mux40~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N4
cycloneive_lcell_comb \Mux40~16 (
// Equation(s):
// \Mux40~16_combout  = (cuifregT_1 & ((\Mux40~13_combout ) # ((cuifregT_01)))) # (!cuifregT_1 & (((!cuifregT_01 & \Mux40~15_combout ))))

	.dataa(\Mux40~13_combout ),
	.datab(cuifregT_1),
	.datac(cuifregT_0),
	.datad(\Mux40~15_combout ),
	.cin(gnd),
	.combout(\Mux40~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~16 .lut_mask = 16'hCBC8;
defparam \Mux40~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y41_N29
dffeas \registerArray[21][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][23] .is_wysiwyg = "true";
defparam \registerArray[21][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N9
dffeas \registerArray[29][23] (
	.clk(clk),
	.d(Mux452),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][23] .is_wysiwyg = "true";
defparam \registerArray[29][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N23
dffeas \registerArray[17][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][23] .is_wysiwyg = "true";
defparam \registerArray[17][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y41_N15
dffeas \registerArray[25][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][23] .is_wysiwyg = "true";
defparam \registerArray[25][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N22
cycloneive_lcell_comb \Mux40~10 (
// Equation(s):
// \Mux40~10_combout  = (cuifregT_2 & (cuifregT_3)) # (!cuifregT_2 & ((cuifregT_3 & ((\registerArray[25][23]~q ))) # (!cuifregT_3 & (\registerArray[17][23]~q ))))

	.dataa(cuifregT_2),
	.datab(cuifregT_3),
	.datac(\registerArray[17][23]~q ),
	.datad(\registerArray[25][23]~q ),
	.cin(gnd),
	.combout(\Mux40~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~10 .lut_mask = 16'hDC98;
defparam \Mux40~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N14
cycloneive_lcell_comb \Mux40~11 (
// Equation(s):
// \Mux40~11_combout  = (\Mux40~10_combout  & (((\registerArray[29][23]~q ) # (!cuifregT_2)))) # (!\Mux40~10_combout  & (\registerArray[21][23]~q  & ((cuifregT_2))))

	.dataa(\registerArray[21][23]~q ),
	.datab(\registerArray[29][23]~q ),
	.datac(\Mux40~10_combout ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux40~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~11 .lut_mask = 16'hCAF0;
defparam \Mux40~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N26
cycloneive_lcell_comb \registerArray[19][23]~feeder (
// Equation(s):
// \registerArray[19][23]~feeder_combout  = \Mux45~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux452),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[19][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[19][23]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[19][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y41_N27
dffeas \registerArray[19][23] (
	.clk(clk),
	.d(\registerArray[19][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][23] .is_wysiwyg = "true";
defparam \registerArray[19][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N12
cycloneive_lcell_comb \Mux40~17 (
// Equation(s):
// \Mux40~17_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[27][23]~q )) # (!cuifregT_3 & ((\registerArray[19][23]~q )))))

	.dataa(\registerArray[27][23]~q ),
	.datab(\registerArray[19][23]~q ),
	.datac(cuifregT_2),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux40~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~17 .lut_mask = 16'hFA0C;
defparam \Mux40~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N3
dffeas \registerArray[31][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][23] .is_wysiwyg = "true";
defparam \registerArray[31][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N28
cycloneive_lcell_comb \registerArray[23][23]~feeder (
// Equation(s):
// \registerArray[23][23]~feeder_combout  = \Mux45~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux452),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[23][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[23][23]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[23][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y41_N29
dffeas \registerArray[23][23] (
	.clk(clk),
	.d(\registerArray[23][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][23] .is_wysiwyg = "true";
defparam \registerArray[23][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N2
cycloneive_lcell_comb \Mux40~18 (
// Equation(s):
// \Mux40~18_combout  = (\Mux40~17_combout  & (((\registerArray[31][23]~q )) # (!cuifregT_2))) # (!\Mux40~17_combout  & (cuifregT_2 & ((\registerArray[23][23]~q ))))

	.dataa(\Mux40~17_combout ),
	.datab(cuifregT_2),
	.datac(\registerArray[31][23]~q ),
	.datad(\registerArray[23][23]~q ),
	.cin(gnd),
	.combout(\Mux40~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~18 .lut_mask = 16'hE6A2;
defparam \Mux40~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N15
dffeas \registerArray[14][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][22] .is_wysiwyg = "true";
defparam \registerArray[14][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N23
dffeas \registerArray[15][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][22] .is_wysiwyg = "true";
defparam \registerArray[15][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N25
dffeas \registerArray[12][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][22] .is_wysiwyg = "true";
defparam \registerArray[12][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N20
cycloneive_lcell_comb \registerArray[13][22]~feeder (
// Equation(s):
// \registerArray[13][22]~feeder_combout  = \Mux46~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux462),
	.cin(gnd),
	.combout(\registerArray[13][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[13][22]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[13][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N21
dffeas \registerArray[13][22] (
	.clk(clk),
	.d(\registerArray[13][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][22] .is_wysiwyg = "true";
defparam \registerArray[13][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N24
cycloneive_lcell_comb \Mux41~7 (
// Equation(s):
// \Mux41~7_combout  = (cuifregT_01 & ((cuifregT_1) # ((\registerArray[13][22]~q )))) # (!cuifregT_01 & (!cuifregT_1 & (\registerArray[12][22]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[12][22]~q ),
	.datad(\registerArray[13][22]~q ),
	.cin(gnd),
	.combout(\Mux41~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~7 .lut_mask = 16'hBA98;
defparam \Mux41~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N22
cycloneive_lcell_comb \Mux41~8 (
// Equation(s):
// \Mux41~8_combout  = (cuifregT_1 & ((\Mux41~7_combout  & ((\registerArray[15][22]~q ))) # (!\Mux41~7_combout  & (\registerArray[14][22]~q )))) # (!cuifregT_1 & (((\Mux41~7_combout ))))

	.dataa(\registerArray[14][22]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[15][22]~q ),
	.datad(\Mux41~7_combout ),
	.cin(gnd),
	.combout(\Mux41~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~8 .lut_mask = 16'hF388;
defparam \Mux41~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N16
cycloneive_lcell_comb \registerArray[9][22]~feeder (
// Equation(s):
// \registerArray[9][22]~feeder_combout  = \Mux46~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux462),
	.cin(gnd),
	.combout(\registerArray[9][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[9][22]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[9][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y43_N17
dffeas \registerArray[9][22] (
	.clk(clk),
	.d(\registerArray[9][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][22] .is_wysiwyg = "true";
defparam \registerArray[9][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N23
dffeas \registerArray[11][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][22] .is_wysiwyg = "true";
defparam \registerArray[11][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N13
dffeas \registerArray[8][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][22] .is_wysiwyg = "true";
defparam \registerArray[8][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N12
cycloneive_lcell_comb \Mux41~0 (
// Equation(s):
// \Mux41~0_combout  = (cuifregT_1 & ((\registerArray[10][22]~q ) # ((cuifregT_01)))) # (!cuifregT_1 & (((\registerArray[8][22]~q  & !cuifregT_01))))

	.dataa(\registerArray[10][22]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[8][22]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux41~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~0 .lut_mask = 16'hCCB8;
defparam \Mux41~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N22
cycloneive_lcell_comb \Mux41~1 (
// Equation(s):
// \Mux41~1_combout  = (cuifregT_01 & ((\Mux41~0_combout  & ((\registerArray[11][22]~q ))) # (!\Mux41~0_combout  & (\registerArray[9][22]~q )))) # (!cuifregT_01 & (((\Mux41~0_combout ))))

	.dataa(\registerArray[9][22]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[11][22]~q ),
	.datad(\Mux41~0_combout ),
	.cin(gnd),
	.combout(\Mux41~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~1 .lut_mask = 16'hF388;
defparam \Mux41~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y41_N11
dffeas \registerArray[2][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][22] .is_wysiwyg = "true";
defparam \registerArray[2][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y41_N13
dffeas \registerArray[1][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][22] .is_wysiwyg = "true";
defparam \registerArray[1][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N12
cycloneive_lcell_comb \Mux41~4 (
// Equation(s):
// \Mux41~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][22]~q )) # (!cuifregT_1 & ((\registerArray[1][22]~q )))))

	.dataa(\registerArray[3][22]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[1][22]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux41~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~4 .lut_mask = 16'h88C0;
defparam \Mux41~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N10
cycloneive_lcell_comb \Mux41~5 (
// Equation(s):
// \Mux41~5_combout  = (\Mux41~4_combout ) # ((cuifregT_1 & (!cuifregT_01 & \registerArray[2][22]~q )))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\registerArray[2][22]~q ),
	.datad(\Mux41~4_combout ),
	.cin(gnd),
	.combout(\Mux41~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~5 .lut_mask = 16'hFF20;
defparam \Mux41~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N9
dffeas \registerArray[7][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][22] .is_wysiwyg = "true";
defparam \registerArray[7][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N11
dffeas \registerArray[4][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][22] .is_wysiwyg = "true";
defparam \registerArray[4][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N9
dffeas \registerArray[5][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][22] .is_wysiwyg = "true";
defparam \registerArray[5][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N10
cycloneive_lcell_comb \Mux41~2 (
// Equation(s):
// \Mux41~2_combout  = (cuifregT_01 & ((cuifregT_1) # ((\registerArray[5][22]~q )))) # (!cuifregT_01 & (!cuifregT_1 & (\registerArray[4][22]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[4][22]~q ),
	.datad(\registerArray[5][22]~q ),
	.cin(gnd),
	.combout(\Mux41~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~2 .lut_mask = 16'hBA98;
defparam \Mux41~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N8
cycloneive_lcell_comb \Mux41~3 (
// Equation(s):
// \Mux41~3_combout  = (cuifregT_1 & ((\Mux41~2_combout  & ((\registerArray[7][22]~q ))) # (!\Mux41~2_combout  & (\registerArray[6][22]~q )))) # (!cuifregT_1 & (((\Mux41~2_combout ))))

	.dataa(\registerArray[6][22]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[7][22]~q ),
	.datad(\Mux41~2_combout ),
	.cin(gnd),
	.combout(\Mux41~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~3 .lut_mask = 16'hF388;
defparam \Mux41~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N28
cycloneive_lcell_comb \Mux41~6 (
// Equation(s):
// \Mux41~6_combout  = (cuifregT_3 & (cuifregT_2)) # (!cuifregT_3 & ((cuifregT_2 & ((\Mux41~3_combout ))) # (!cuifregT_2 & (\Mux41~5_combout ))))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\Mux41~5_combout ),
	.datad(\Mux41~3_combout ),
	.cin(gnd),
	.combout(\Mux41~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~6 .lut_mask = 16'hDC98;
defparam \Mux41~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N26
cycloneive_lcell_comb \registerArray[31][22]~feeder (
// Equation(s):
// \registerArray[31][22]~feeder_combout  = \Mux46~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux462),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[31][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[31][22]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[31][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N27
dffeas \registerArray[31][22] (
	.clk(clk),
	.d(\registerArray[31][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][22] .is_wysiwyg = "true";
defparam \registerArray[31][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N5
dffeas \registerArray[27][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][22] .is_wysiwyg = "true";
defparam \registerArray[27][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N11
dffeas \registerArray[19][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][22] .is_wysiwyg = "true";
defparam \registerArray[19][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N10
cycloneive_lcell_comb \Mux41~17 (
// Equation(s):
// \Mux41~17_combout  = (cuifregT_2 & ((\registerArray[23][22]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[19][22]~q  & !cuifregT_3))))

	.dataa(\registerArray[23][22]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[19][22]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux41~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~17 .lut_mask = 16'hCCB8;
defparam \Mux41~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N12
cycloneive_lcell_comb \Mux41~18 (
// Equation(s):
// \Mux41~18_combout  = (cuifregT_3 & ((\Mux41~17_combout  & (\registerArray[31][22]~q )) # (!\Mux41~17_combout  & ((\registerArray[27][22]~q ))))) # (!cuifregT_3 & (((\Mux41~17_combout ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[31][22]~q ),
	.datac(\registerArray[27][22]~q ),
	.datad(\Mux41~17_combout ),
	.cin(gnd),
	.combout(\Mux41~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~18 .lut_mask = 16'hDDA0;
defparam \Mux41~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y41_N9
dffeas \registerArray[25][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][22] .is_wysiwyg = "true";
defparam \registerArray[25][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N7
dffeas \registerArray[29][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][22] .is_wysiwyg = "true";
defparam \registerArray[29][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N29
dffeas \registerArray[17][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][22] .is_wysiwyg = "true";
defparam \registerArray[17][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y41_N23
dffeas \registerArray[21][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][22] .is_wysiwyg = "true";
defparam \registerArray[21][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N28
cycloneive_lcell_comb \Mux41~10 (
// Equation(s):
// \Mux41~10_combout  = (cuifregT_2 & ((cuifregT_3) # ((\registerArray[21][22]~q )))) # (!cuifregT_2 & (!cuifregT_3 & (\registerArray[17][22]~q )))

	.dataa(cuifregT_2),
	.datab(cuifregT_3),
	.datac(\registerArray[17][22]~q ),
	.datad(\registerArray[21][22]~q ),
	.cin(gnd),
	.combout(\Mux41~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~10 .lut_mask = 16'hBA98;
defparam \Mux41~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N6
cycloneive_lcell_comb \Mux41~11 (
// Equation(s):
// \Mux41~11_combout  = (cuifregT_3 & ((\Mux41~10_combout  & ((\registerArray[29][22]~q ))) # (!\Mux41~10_combout  & (\registerArray[25][22]~q )))) # (!cuifregT_3 & (((\Mux41~10_combout ))))

	.dataa(\registerArray[25][22]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[29][22]~q ),
	.datad(\Mux41~10_combout ),
	.cin(gnd),
	.combout(\Mux41~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~11 .lut_mask = 16'hF388;
defparam \Mux41~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N29
dffeas \registerArray[22][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][22] .is_wysiwyg = "true";
defparam \registerArray[22][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N23
dffeas \registerArray[30][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][22] .is_wysiwyg = "true";
defparam \registerArray[30][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N31
dffeas \registerArray[26][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][22] .is_wysiwyg = "true";
defparam \registerArray[26][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N17
dffeas \registerArray[18][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][22] .is_wysiwyg = "true";
defparam \registerArray[18][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N16
cycloneive_lcell_comb \Mux41~12 (
// Equation(s):
// \Mux41~12_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[26][22]~q )) # (!cuifregT_3 & ((\registerArray[18][22]~q )))))

	.dataa(cuifregT_2),
	.datab(\registerArray[26][22]~q ),
	.datac(\registerArray[18][22]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux41~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~12 .lut_mask = 16'hEE50;
defparam \Mux41~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N22
cycloneive_lcell_comb \Mux41~13 (
// Equation(s):
// \Mux41~13_combout  = (cuifregT_2 & ((\Mux41~12_combout  & ((\registerArray[30][22]~q ))) # (!\Mux41~12_combout  & (\registerArray[22][22]~q )))) # (!cuifregT_2 & (((\Mux41~12_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[22][22]~q ),
	.datac(\registerArray[30][22]~q ),
	.datad(\Mux41~12_combout ),
	.cin(gnd),
	.combout(\Mux41~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~13 .lut_mask = 16'hF588;
defparam \Mux41~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N21
dffeas \registerArray[16][22] (
	.clk(clk),
	.d(Mux462),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][22] .is_wysiwyg = "true";
defparam \registerArray[16][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y35_N9
dffeas \registerArray[24][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][22] .is_wysiwyg = "true";
defparam \registerArray[24][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N8
cycloneive_lcell_comb \Mux41~14 (
// Equation(s):
// \Mux41~14_combout  = (cuifregT_3 & (((\registerArray[24][22]~q ) # (cuifregT_2)))) # (!cuifregT_3 & (\registerArray[16][22]~q  & ((!cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[16][22]~q ),
	.datac(\registerArray[24][22]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux41~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~14 .lut_mask = 16'hAAE4;
defparam \Mux41~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N14
cycloneive_lcell_comb \registerArray[28][22]~feeder (
// Equation(s):
// \registerArray[28][22]~feeder_combout  = \Mux46~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux462),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[28][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[28][22]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[28][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y35_N15
dffeas \registerArray[28][22] (
	.clk(clk),
	.d(\registerArray[28][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][22] .is_wysiwyg = "true";
defparam \registerArray[28][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N4
cycloneive_lcell_comb \Mux41~15 (
// Equation(s):
// \Mux41~15_combout  = (\Mux41~14_combout  & (((\registerArray[28][22]~q ) # (!cuifregT_2)))) # (!\Mux41~14_combout  & (\registerArray[20][22]~q  & ((cuifregT_2))))

	.dataa(\registerArray[20][22]~q ),
	.datab(\Mux41~14_combout ),
	.datac(\registerArray[28][22]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux41~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~15 .lut_mask = 16'hE2CC;
defparam \Mux41~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y35_N2
cycloneive_lcell_comb \Mux41~16 (
// Equation(s):
// \Mux41~16_combout  = (cuifregT_1 & ((cuifregT_01) # ((\Mux41~13_combout )))) # (!cuifregT_1 & (!cuifregT_01 & ((\Mux41~15_combout ))))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\Mux41~13_combout ),
	.datad(\Mux41~15_combout ),
	.cin(gnd),
	.combout(\Mux41~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~16 .lut_mask = 16'hB9A8;
defparam \Mux41~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y44_N13
dffeas \registerArray[14][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][21] .is_wysiwyg = "true";
defparam \registerArray[14][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N15
dffeas \registerArray[15][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][21] .is_wysiwyg = "true";
defparam \registerArray[15][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N21
dffeas \registerArray[12][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][21] .is_wysiwyg = "true";
defparam \registerArray[12][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y44_N7
dffeas \registerArray[13][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][21] .is_wysiwyg = "true";
defparam \registerArray[13][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N20
cycloneive_lcell_comb \Mux42~7 (
// Equation(s):
// \Mux42~7_combout  = (cuifregT_01 & ((cuifregT_1) # ((\registerArray[13][21]~q )))) # (!cuifregT_01 & (!cuifregT_1 & (\registerArray[12][21]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[12][21]~q ),
	.datad(\registerArray[13][21]~q ),
	.cin(gnd),
	.combout(\Mux42~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~7 .lut_mask = 16'hBA98;
defparam \Mux42~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N14
cycloneive_lcell_comb \Mux42~8 (
// Equation(s):
// \Mux42~8_combout  = (cuifregT_1 & ((\Mux42~7_combout  & ((\registerArray[15][21]~q ))) # (!\Mux42~7_combout  & (\registerArray[14][21]~q )))) # (!cuifregT_1 & (((\Mux42~7_combout ))))

	.dataa(\registerArray[14][21]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[15][21]~q ),
	.datad(\Mux42~7_combout ),
	.cin(gnd),
	.combout(\Mux42~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~8 .lut_mask = 16'hF388;
defparam \Mux42~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y42_N27
dffeas \registerArray[2][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][21] .is_wysiwyg = "true";
defparam \registerArray[2][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N30
cycloneive_lcell_comb \registerArray[1][21]~feeder (
// Equation(s):
// \registerArray[1][21]~feeder_combout  = \Mux47~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux472),
	.cin(gnd),
	.combout(\registerArray[1][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[1][21]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[1][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y42_N31
dffeas \registerArray[1][21] (
	.clk(clk),
	.d(\registerArray[1][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][21] .is_wysiwyg = "true";
defparam \registerArray[1][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N16
cycloneive_lcell_comb \Mux42~4 (
// Equation(s):
// \Mux42~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][21]~q )) # (!cuifregT_1 & ((\registerArray[1][21]~q )))))

	.dataa(\registerArray[3][21]~q ),
	.datab(\registerArray[1][21]~q ),
	.datac(cuifregT_1),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux42~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~4 .lut_mask = 16'hAC00;
defparam \Mux42~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N26
cycloneive_lcell_comb \Mux42~5 (
// Equation(s):
// \Mux42~5_combout  = (\Mux42~4_combout ) # ((!cuifregT_01 & (cuifregT_1 & \registerArray[2][21]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[2][21]~q ),
	.datad(\Mux42~4_combout ),
	.cin(gnd),
	.combout(\Mux42~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~5 .lut_mask = 16'hFF40;
defparam \Mux42~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y43_N1
dffeas \registerArray[9][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][21] .is_wysiwyg = "true";
defparam \registerArray[9][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N5
dffeas \registerArray[8][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][21] .is_wysiwyg = "true";
defparam \registerArray[8][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N4
cycloneive_lcell_comb \Mux42~2 (
// Equation(s):
// \Mux42~2_combout  = (cuifregT_1 & ((\registerArray[10][21]~q ) # ((cuifregT_01)))) # (!cuifregT_1 & (((\registerArray[8][21]~q  & !cuifregT_01))))

	.dataa(\registerArray[10][21]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[8][21]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux42~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~2 .lut_mask = 16'hCCB8;
defparam \Mux42~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N24
cycloneive_lcell_comb \Mux42~3 (
// Equation(s):
// \Mux42~3_combout  = (cuifregT_01 & ((\Mux42~2_combout  & (\registerArray[11][21]~q )) # (!\Mux42~2_combout  & ((\registerArray[9][21]~q ))))) # (!cuifregT_01 & (((\Mux42~2_combout ))))

	.dataa(\registerArray[11][21]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[9][21]~q ),
	.datad(\Mux42~2_combout ),
	.cin(gnd),
	.combout(\Mux42~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~3 .lut_mask = 16'hBBC0;
defparam \Mux42~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N26
cycloneive_lcell_comb \Mux42~6 (
// Equation(s):
// \Mux42~6_combout  = (cuifregT_2 & (cuifregT_3)) # (!cuifregT_2 & ((cuifregT_3 & ((\Mux42~3_combout ))) # (!cuifregT_3 & (\Mux42~5_combout ))))

	.dataa(cuifregT_2),
	.datab(cuifregT_3),
	.datac(\Mux42~5_combout ),
	.datad(\Mux42~3_combout ),
	.cin(gnd),
	.combout(\Mux42~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~6 .lut_mask = 16'hDC98;
defparam \Mux42~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N20
cycloneive_lcell_comb \registerArray[6][21]~feeder (
// Equation(s):
// \registerArray[6][21]~feeder_combout  = \Mux47~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux472),
	.cin(gnd),
	.combout(\registerArray[6][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[6][21]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[6][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y44_N21
dffeas \registerArray[6][21] (
	.clk(clk),
	.d(\registerArray[6][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][21] .is_wysiwyg = "true";
defparam \registerArray[6][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N15
dffeas \registerArray[7][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][21] .is_wysiwyg = "true";
defparam \registerArray[7][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N19
dffeas \registerArray[4][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][21] .is_wysiwyg = "true";
defparam \registerArray[4][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N18
cycloneive_lcell_comb \Mux42~0 (
// Equation(s):
// \Mux42~0_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[5][21]~q )) # (!cuifregT_01 & ((\registerArray[4][21]~q )))))

	.dataa(\registerArray[5][21]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[4][21]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux42~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~0 .lut_mask = 16'hEE30;
defparam \Mux42~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N14
cycloneive_lcell_comb \Mux42~1 (
// Equation(s):
// \Mux42~1_combout  = (cuifregT_1 & ((\Mux42~0_combout  & ((\registerArray[7][21]~q ))) # (!\Mux42~0_combout  & (\registerArray[6][21]~q )))) # (!cuifregT_1 & (((\Mux42~0_combout ))))

	.dataa(\registerArray[6][21]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[7][21]~q ),
	.datad(\Mux42~0_combout ),
	.cin(gnd),
	.combout(\Mux42~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~1 .lut_mask = 16'hF388;
defparam \Mux42~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N26
cycloneive_lcell_comb \registerArray[21][21]~feeder (
// Equation(s):
// \registerArray[21][21]~feeder_combout  = \Mux47~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux472),
	.cin(gnd),
	.combout(\registerArray[21][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[21][21]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[21][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y44_N27
dffeas \registerArray[21][21] (
	.clk(clk),
	.d(\registerArray[21][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][21] .is_wysiwyg = "true";
defparam \registerArray[21][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N13
dffeas \registerArray[29][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][21] .is_wysiwyg = "true";
defparam \registerArray[29][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N4
cycloneive_lcell_comb \registerArray[17][21]~feeder (
// Equation(s):
// \registerArray[17][21]~feeder_combout  = \Mux47~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux472),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[17][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[17][21]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[17][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N5
dffeas \registerArray[17][21] (
	.clk(clk),
	.d(\registerArray[17][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][21] .is_wysiwyg = "true";
defparam \registerArray[17][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N24
cycloneive_lcell_comb \registerArray[25][21]~feeder (
// Equation(s):
// \registerArray[25][21]~feeder_combout  = \Mux47~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux472),
	.cin(gnd),
	.combout(\registerArray[25][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[25][21]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[25][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y44_N25
dffeas \registerArray[25][21] (
	.clk(clk),
	.d(\registerArray[25][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][21] .is_wysiwyg = "true";
defparam \registerArray[25][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N10
cycloneive_lcell_comb \Mux42~10 (
// Equation(s):
// \Mux42~10_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & ((\registerArray[25][21]~q ))) # (!cuifregT_3 & (\registerArray[17][21]~q ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[17][21]~q ),
	.datac(cuifregT_3),
	.datad(\registerArray[25][21]~q ),
	.cin(gnd),
	.combout(\Mux42~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~10 .lut_mask = 16'hF4A4;
defparam \Mux42~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N12
cycloneive_lcell_comb \Mux42~11 (
// Equation(s):
// \Mux42~11_combout  = (cuifregT_2 & ((\Mux42~10_combout  & ((\registerArray[29][21]~q ))) # (!\Mux42~10_combout  & (\registerArray[21][21]~q )))) # (!cuifregT_2 & (((\Mux42~10_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[21][21]~q ),
	.datac(\registerArray[29][21]~q ),
	.datad(\Mux42~10_combout ),
	.cin(gnd),
	.combout(\Mux42~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~11 .lut_mask = 16'hF588;
defparam \Mux42~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N26
cycloneive_lcell_comb \registerArray[31][21]~feeder (
// Equation(s):
// \registerArray[31][21]~feeder_combout  = \Mux47~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux472),
	.cin(gnd),
	.combout(\registerArray[31][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[31][21]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[31][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N27
dffeas \registerArray[31][21] (
	.clk(clk),
	.d(\registerArray[31][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][21] .is_wysiwyg = "true";
defparam \registerArray[31][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N17
dffeas \registerArray[23][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][21] .is_wysiwyg = "true";
defparam \registerArray[23][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N19
dffeas \registerArray[19][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][21] .is_wysiwyg = "true";
defparam \registerArray[19][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N18
cycloneive_lcell_comb \Mux42~17 (
// Equation(s):
// \Mux42~17_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[27][21]~q )) # (!cuifregT_3 & ((\registerArray[19][21]~q )))))

	.dataa(\registerArray[27][21]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[19][21]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux42~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~17 .lut_mask = 16'hEE30;
defparam \Mux42~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N8
cycloneive_lcell_comb \Mux42~18 (
// Equation(s):
// \Mux42~18_combout  = (cuifregT_2 & ((\Mux42~17_combout  & (\registerArray[31][21]~q )) # (!\Mux42~17_combout  & ((\registerArray[23][21]~q ))))) # (!cuifregT_2 & (((\Mux42~17_combout ))))

	.dataa(\registerArray[31][21]~q ),
	.datab(\registerArray[23][21]~q ),
	.datac(cuifregT_2),
	.datad(\Mux42~17_combout ),
	.cin(gnd),
	.combout(\Mux42~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~18 .lut_mask = 16'hAFC0;
defparam \Mux42~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y31_N31
dffeas \registerArray[28][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][21] .is_wysiwyg = "true";
defparam \registerArray[28][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y40_N11
dffeas \registerArray[20][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][21] .is_wysiwyg = "true";
defparam \registerArray[20][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N28
cycloneive_lcell_comb \Mux42~14 (
// Equation(s):
// \Mux42~14_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & ((\registerArray[20][21]~q ))) # (!cuifregT_2 & (\registerArray[16][21]~q ))))

	.dataa(\registerArray[16][21]~q ),
	.datab(\registerArray[20][21]~q ),
	.datac(cuifregT_3),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux42~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~14 .lut_mask = 16'hFC0A;
defparam \Mux42~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N30
cycloneive_lcell_comb \Mux42~15 (
// Equation(s):
// \Mux42~15_combout  = (cuifregT_3 & ((\Mux42~14_combout  & ((\registerArray[28][21]~q ))) # (!\Mux42~14_combout  & (\registerArray[24][21]~q )))) # (!cuifregT_3 & (((\Mux42~14_combout ))))

	.dataa(\registerArray[24][21]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[28][21]~q ),
	.datad(\Mux42~14_combout ),
	.cin(gnd),
	.combout(\Mux42~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~15 .lut_mask = 16'hF388;
defparam \Mux42~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N3
dffeas \registerArray[30][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][21] .is_wysiwyg = "true";
defparam \registerArray[30][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N1
dffeas \registerArray[18][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][21] .is_wysiwyg = "true";
defparam \registerArray[18][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N0
cycloneive_lcell_comb \Mux42~12 (
// Equation(s):
// \Mux42~12_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[22][21]~q )) # (!cuifregT_2 & ((\registerArray[18][21]~q )))))

	.dataa(\registerArray[22][21]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[18][21]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux42~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~12 .lut_mask = 16'hEE30;
defparam \Mux42~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N2
cycloneive_lcell_comb \Mux42~13 (
// Equation(s):
// \Mux42~13_combout  = (cuifregT_3 & ((\Mux42~12_combout  & ((\registerArray[30][21]~q ))) # (!\Mux42~12_combout  & (\registerArray[26][21]~q )))) # (!cuifregT_3 & (((\Mux42~12_combout ))))

	.dataa(\registerArray[26][21]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[30][21]~q ),
	.datad(\Mux42~12_combout ),
	.cin(gnd),
	.combout(\Mux42~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~13 .lut_mask = 16'hF388;
defparam \Mux42~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N16
cycloneive_lcell_comb \Mux42~16 (
// Equation(s):
// \Mux42~16_combout  = (cuifregT_1 & ((cuifregT_01) # ((\Mux42~13_combout )))) # (!cuifregT_1 & (!cuifregT_01 & (\Mux42~15_combout )))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\Mux42~15_combout ),
	.datad(\Mux42~13_combout ),
	.cin(gnd),
	.combout(\Mux42~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~16 .lut_mask = 16'hBA98;
defparam \Mux42~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N31
dffeas \registerArray[14][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][20] .is_wysiwyg = "true";
defparam \registerArray[14][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N11
dffeas \registerArray[15][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][20] .is_wysiwyg = "true";
defparam \registerArray[15][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N13
dffeas \registerArray[12][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][20] .is_wysiwyg = "true";
defparam \registerArray[12][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N31
dffeas \registerArray[13][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][20] .is_wysiwyg = "true";
defparam \registerArray[13][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N12
cycloneive_lcell_comb \Mux43~7 (
// Equation(s):
// \Mux43~7_combout  = (cuifregT_01 & ((cuifregT_1) # ((\registerArray[13][20]~q )))) # (!cuifregT_01 & (!cuifregT_1 & (\registerArray[12][20]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[12][20]~q ),
	.datad(\registerArray[13][20]~q ),
	.cin(gnd),
	.combout(\Mux43~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~7 .lut_mask = 16'hBA98;
defparam \Mux43~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N10
cycloneive_lcell_comb \Mux43~8 (
// Equation(s):
// \Mux43~8_combout  = (cuifregT_1 & ((\Mux43~7_combout  & ((\registerArray[15][20]~q ))) # (!\Mux43~7_combout  & (\registerArray[14][20]~q )))) # (!cuifregT_1 & (((\Mux43~7_combout ))))

	.dataa(\registerArray[14][20]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[15][20]~q ),
	.datad(\Mux43~7_combout ),
	.cin(gnd),
	.combout(\Mux43~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~8 .lut_mask = 16'hF388;
defparam \Mux43~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N24
cycloneive_lcell_comb \registerArray[11][20]~feeder (
// Equation(s):
// \registerArray[11][20]~feeder_combout  = \Mux48~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux482),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[11][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[11][20]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[11][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y42_N25
dffeas \registerArray[11][20] (
	.clk(clk),
	.d(\registerArray[11][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][20] .is_wysiwyg = "true";
defparam \registerArray[11][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N14
cycloneive_lcell_comb \registerArray[9][20]~feeder (
// Equation(s):
// \registerArray[9][20]~feeder_combout  = \Mux48~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux482),
	.cin(gnd),
	.combout(\registerArray[9][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[9][20]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[9][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N15
dffeas \registerArray[9][20] (
	.clk(clk),
	.d(\registerArray[9][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][20] .is_wysiwyg = "true";
defparam \registerArray[9][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N27
dffeas \registerArray[8][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][20] .is_wysiwyg = "true";
defparam \registerArray[8][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N26
cycloneive_lcell_comb \Mux43~0 (
// Equation(s):
// \Mux43~0_combout  = (cuifregT_1 & ((\registerArray[10][20]~q ) # ((cuifregT_01)))) # (!cuifregT_1 & (((\registerArray[8][20]~q  & !cuifregT_01))))

	.dataa(\registerArray[10][20]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[8][20]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux43~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~0 .lut_mask = 16'hCCB8;
defparam \Mux43~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N0
cycloneive_lcell_comb \Mux43~1 (
// Equation(s):
// \Mux43~1_combout  = (cuifregT_01 & ((\Mux43~0_combout  & (\registerArray[11][20]~q )) # (!\Mux43~0_combout  & ((\registerArray[9][20]~q ))))) # (!cuifregT_01 & (((\Mux43~0_combout ))))

	.dataa(cuifregT_0),
	.datab(\registerArray[11][20]~q ),
	.datac(\registerArray[9][20]~q ),
	.datad(\Mux43~0_combout ),
	.cin(gnd),
	.combout(\Mux43~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~1 .lut_mask = 16'hDDA0;
defparam \Mux43~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N19
dffeas \registerArray[7][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][20] .is_wysiwyg = "true";
defparam \registerArray[7][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N3
dffeas \registerArray[4][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][20] .is_wysiwyg = "true";
defparam \registerArray[4][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N2
cycloneive_lcell_comb \Mux43~2 (
// Equation(s):
// \Mux43~2_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[5][20]~q )) # (!cuifregT_01 & ((\registerArray[4][20]~q )))))

	.dataa(\registerArray[5][20]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[4][20]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux43~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~2 .lut_mask = 16'hEE30;
defparam \Mux43~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N18
cycloneive_lcell_comb \Mux43~3 (
// Equation(s):
// \Mux43~3_combout  = (cuifregT_1 & ((\Mux43~2_combout  & ((\registerArray[7][20]~q ))) # (!\Mux43~2_combout  & (\registerArray[6][20]~q )))) # (!cuifregT_1 & (((\Mux43~2_combout ))))

	.dataa(\registerArray[6][20]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[7][20]~q ),
	.datad(\Mux43~2_combout ),
	.cin(gnd),
	.combout(\Mux43~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~3 .lut_mask = 16'hF388;
defparam \Mux43~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y42_N19
dffeas \registerArray[2][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][20] .is_wysiwyg = "true";
defparam \registerArray[2][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y42_N29
dffeas \registerArray[1][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][20] .is_wysiwyg = "true";
defparam \registerArray[1][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N28
cycloneive_lcell_comb \Mux43~4 (
// Equation(s):
// \Mux43~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][20]~q )) # (!cuifregT_1 & ((\registerArray[1][20]~q )))))

	.dataa(\registerArray[3][20]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[1][20]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux43~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~4 .lut_mask = 16'hB800;
defparam \Mux43~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N18
cycloneive_lcell_comb \Mux43~5 (
// Equation(s):
// \Mux43~5_combout  = (\Mux43~4_combout ) # ((!cuifregT_01 & (cuifregT_1 & \registerArray[2][20]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[2][20]~q ),
	.datad(\Mux43~4_combout ),
	.cin(gnd),
	.combout(\Mux43~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~5 .lut_mask = 16'hFF40;
defparam \Mux43~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N24
cycloneive_lcell_comb \Mux43~6 (
// Equation(s):
// \Mux43~6_combout  = (cuifregT_2 & ((cuifregT_3) # ((\Mux43~3_combout )))) # (!cuifregT_2 & (!cuifregT_3 & ((\Mux43~5_combout ))))

	.dataa(cuifregT_2),
	.datab(cuifregT_3),
	.datac(\Mux43~3_combout ),
	.datad(\Mux43~5_combout ),
	.cin(gnd),
	.combout(\Mux43~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~6 .lut_mask = 16'hB9A8;
defparam \Mux43~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N0
cycloneive_lcell_comb \registerArray[16][20]~feeder (
// Equation(s):
// \registerArray[16][20]~feeder_combout  = \Mux48~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux482),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[16][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[16][20]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[16][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N1
dffeas \registerArray[16][20] (
	.clk(clk),
	.d(\registerArray[16][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][20] .is_wysiwyg = "true";
defparam \registerArray[16][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y38_N15
dffeas \registerArray[24][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][20] .is_wysiwyg = "true";
defparam \registerArray[24][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N14
cycloneive_lcell_comb \Mux43~14 (
// Equation(s):
// \Mux43~14_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & ((\registerArray[24][20]~q ))) # (!cuifregT_3 & (\registerArray[16][20]~q ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[16][20]~q ),
	.datac(\registerArray[24][20]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux43~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~14 .lut_mask = 16'hFA44;
defparam \Mux43~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y38_N9
dffeas \registerArray[28][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][20] .is_wysiwyg = "true";
defparam \registerArray[28][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N8
cycloneive_lcell_comb \Mux43~15 (
// Equation(s):
// \Mux43~15_combout  = (\Mux43~14_combout  & (((\registerArray[28][20]~q ) # (!cuifregT_2)))) # (!\Mux43~14_combout  & (\registerArray[20][20]~q  & ((cuifregT_2))))

	.dataa(\registerArray[20][20]~q ),
	.datab(\Mux43~14_combout ),
	.datac(\registerArray[28][20]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux43~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~15 .lut_mask = 16'hE2CC;
defparam \Mux43~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N25
dffeas \registerArray[22][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][20] .is_wysiwyg = "true";
defparam \registerArray[22][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N19
dffeas \registerArray[30][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][20] .is_wysiwyg = "true";
defparam \registerArray[30][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N28
cycloneive_lcell_comb \registerArray[26][20]~feeder (
// Equation(s):
// \registerArray[26][20]~feeder_combout  = \Mux48~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux482),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[26][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[26][20]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[26][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y44_N29
dffeas \registerArray[26][20] (
	.clk(clk),
	.d(\registerArray[26][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][20] .is_wysiwyg = "true";
defparam \registerArray[26][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N13
dffeas \registerArray[18][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][20] .is_wysiwyg = "true";
defparam \registerArray[18][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N12
cycloneive_lcell_comb \Mux43~12 (
// Equation(s):
// \Mux43~12_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[26][20]~q )) # (!cuifregT_3 & ((\registerArray[18][20]~q )))))

	.dataa(cuifregT_2),
	.datab(\registerArray[26][20]~q ),
	.datac(\registerArray[18][20]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux43~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~12 .lut_mask = 16'hEE50;
defparam \Mux43~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N18
cycloneive_lcell_comb \Mux43~13 (
// Equation(s):
// \Mux43~13_combout  = (cuifregT_2 & ((\Mux43~12_combout  & ((\registerArray[30][20]~q ))) # (!\Mux43~12_combout  & (\registerArray[22][20]~q )))) # (!cuifregT_2 & (((\Mux43~12_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[22][20]~q ),
	.datac(\registerArray[30][20]~q ),
	.datad(\Mux43~12_combout ),
	.cin(gnd),
	.combout(\Mux43~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~13 .lut_mask = 16'hF588;
defparam \Mux43~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y38_N22
cycloneive_lcell_comb \Mux43~16 (
// Equation(s):
// \Mux43~16_combout  = (cuifregT_1 & ((cuifregT_01) # ((\Mux43~13_combout )))) # (!cuifregT_1 & (!cuifregT_01 & (\Mux43~15_combout )))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\Mux43~15_combout ),
	.datad(\Mux43~13_combout ),
	.cin(gnd),
	.combout(\Mux43~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~16 .lut_mask = 16'hBA98;
defparam \Mux43~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y41_N17
dffeas \registerArray[25][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][20] .is_wysiwyg = "true";
defparam \registerArray[25][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N21
dffeas \registerArray[29][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][20] .is_wysiwyg = "true";
defparam \registerArray[29][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N7
dffeas \registerArray[17][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][20] .is_wysiwyg = "true";
defparam \registerArray[17][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N6
cycloneive_lcell_comb \Mux43~10 (
// Equation(s):
// \Mux43~10_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[21][20]~q )) # (!cuifregT_2 & ((\registerArray[17][20]~q )))))

	.dataa(\registerArray[21][20]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[17][20]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux43~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~10 .lut_mask = 16'hEE30;
defparam \Mux43~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N20
cycloneive_lcell_comb \Mux43~11 (
// Equation(s):
// \Mux43~11_combout  = (cuifregT_3 & ((\Mux43~10_combout  & ((\registerArray[29][20]~q ))) # (!\Mux43~10_combout  & (\registerArray[25][20]~q )))) # (!cuifregT_3 & (((\Mux43~10_combout ))))

	.dataa(\registerArray[25][20]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[29][20]~q ),
	.datad(\Mux43~10_combout ),
	.cin(gnd),
	.combout(\Mux43~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~11 .lut_mask = 16'hF388;
defparam \Mux43~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N21
dffeas \registerArray[27][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][20] .is_wysiwyg = "true";
defparam \registerArray[27][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y41_N29
dffeas \registerArray[31][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][20] .is_wysiwyg = "true";
defparam \registerArray[31][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N0
cycloneive_lcell_comb \registerArray[19][20]~feeder (
// Equation(s):
// \registerArray[19][20]~feeder_combout  = \Mux48~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux482),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[19][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[19][20]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[19][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y41_N1
dffeas \registerArray[19][20] (
	.clk(clk),
	.d(\registerArray[19][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][20] .is_wysiwyg = "true";
defparam \registerArray[19][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N10
cycloneive_lcell_comb \Mux43~17 (
// Equation(s):
// \Mux43~17_combout  = (cuifregT_2 & ((\registerArray[23][20]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[19][20]~q  & !cuifregT_3))))

	.dataa(\registerArray[23][20]~q ),
	.datab(\registerArray[19][20]~q ),
	.datac(cuifregT_2),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux43~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~17 .lut_mask = 16'hF0AC;
defparam \Mux43~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N28
cycloneive_lcell_comb \Mux43~18 (
// Equation(s):
// \Mux43~18_combout  = (cuifregT_3 & ((\Mux43~17_combout  & ((\registerArray[31][20]~q ))) # (!\Mux43~17_combout  & (\registerArray[27][20]~q )))) # (!cuifregT_3 & (((\Mux43~17_combout ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[27][20]~q ),
	.datac(\registerArray[31][20]~q ),
	.datad(\Mux43~17_combout ),
	.cin(gnd),
	.combout(\Mux43~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~18 .lut_mask = 16'hF588;
defparam \Mux43~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N28
cycloneive_lcell_comb \registerArray[14][5]~feeder (
// Equation(s):
// \registerArray[14][5]~feeder_combout  = \Mux63~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux632),
	.cin(gnd),
	.combout(\registerArray[14][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][5]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[14][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y32_N29
dffeas \registerArray[14][5] (
	.clk(clk),
	.d(\registerArray[14][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][5] .is_wysiwyg = "true";
defparam \registerArray[14][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N31
dffeas \registerArray[15][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][5] .is_wysiwyg = "true";
defparam \registerArray[15][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N13
dffeas \registerArray[12][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][5] .is_wysiwyg = "true";
defparam \registerArray[12][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N12
cycloneive_lcell_comb \Mux58~7 (
// Equation(s):
// \Mux58~7_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[13][5]~q )) # (!cuifregT_01 & ((\registerArray[12][5]~q )))))

	.dataa(\registerArray[13][5]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[12][5]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux58~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~7 .lut_mask = 16'hEE30;
defparam \Mux58~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N30
cycloneive_lcell_comb \Mux58~8 (
// Equation(s):
// \Mux58~8_combout  = (cuifregT_1 & ((\Mux58~7_combout  & ((\registerArray[15][5]~q ))) # (!\Mux58~7_combout  & (\registerArray[14][5]~q )))) # (!cuifregT_1 & (((\Mux58~7_combout ))))

	.dataa(\registerArray[14][5]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[15][5]~q ),
	.datad(\Mux58~7_combout ),
	.cin(gnd),
	.combout(\Mux58~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~8 .lut_mask = 16'hF388;
defparam \Mux58~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N28
cycloneive_lcell_comb \registerArray[6][5]~feeder (
// Equation(s):
// \registerArray[6][5]~feeder_combout  = \Mux63~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux632),
	.cin(gnd),
	.combout(\registerArray[6][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[6][5]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[6][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y30_N29
dffeas \registerArray[6][5] (
	.clk(clk),
	.d(\registerArray[6][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][5] .is_wysiwyg = "true";
defparam \registerArray[6][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N17
dffeas \registerArray[7][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][5] .is_wysiwyg = "true";
defparam \registerArray[7][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N28
cycloneive_lcell_comb \registerArray[4][5]~feeder (
// Equation(s):
// \registerArray[4][5]~feeder_combout  = \Mux63~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux632),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[4][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[4][5]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[4][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y31_N29
dffeas \registerArray[4][5] (
	.clk(clk),
	.d(\registerArray[4][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][5] .is_wysiwyg = "true";
defparam \registerArray[4][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N6
cycloneive_lcell_comb \Mux58~0 (
// Equation(s):
// \Mux58~0_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[5][5]~q )) # (!cuifregT_01 & ((\registerArray[4][5]~q )))))

	.dataa(\registerArray[5][5]~q ),
	.datab(\registerArray[4][5]~q ),
	.datac(cuifregT_1),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux58~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~0 .lut_mask = 16'hFA0C;
defparam \Mux58~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N16
cycloneive_lcell_comb \Mux58~1 (
// Equation(s):
// \Mux58~1_combout  = (cuifregT_1 & ((\Mux58~0_combout  & ((\registerArray[7][5]~q ))) # (!\Mux58~0_combout  & (\registerArray[6][5]~q )))) # (!cuifregT_1 & (((\Mux58~0_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[6][5]~q ),
	.datac(\registerArray[7][5]~q ),
	.datad(\Mux58~0_combout ),
	.cin(gnd),
	.combout(\Mux58~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~1 .lut_mask = 16'hF588;
defparam \Mux58~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y43_N9
dffeas \registerArray[3][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][5] .is_wysiwyg = "true";
defparam \registerArray[3][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N6
cycloneive_lcell_comb \Mux58~4 (
// Equation(s):
// \Mux58~4_combout  = (cuifregT_01 & ((cuifregT_1 & ((\registerArray[3][5]~q ))) # (!cuifregT_1 & (\registerArray[1][5]~q ))))

	.dataa(\registerArray[1][5]~q ),
	.datab(\registerArray[3][5]~q ),
	.datac(cuifregT_1),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux58~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~4 .lut_mask = 16'hCA00;
defparam \Mux58~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N22
cycloneive_lcell_comb \Mux58~5 (
// Equation(s):
// \Mux58~5_combout  = (\Mux58~4_combout ) # ((\registerArray[2][5]~q  & (!cuifregT_01 & cuifregT_1)))

	.dataa(\registerArray[2][5]~q ),
	.datab(cuifregT_0),
	.datac(cuifregT_1),
	.datad(\Mux58~4_combout ),
	.cin(gnd),
	.combout(\Mux58~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~5 .lut_mask = 16'hFF20;
defparam \Mux58~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N5
dffeas \registerArray[9][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][5] .is_wysiwyg = "true";
defparam \registerArray[9][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N1
dffeas \registerArray[8][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][5] .is_wysiwyg = "true";
defparam \registerArray[8][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N0
cycloneive_lcell_comb \Mux58~2 (
// Equation(s):
// \Mux58~2_combout  = (cuifregT_1 & ((\registerArray[10][5]~q ) # ((cuifregT_01)))) # (!cuifregT_1 & (((\registerArray[8][5]~q  & !cuifregT_01))))

	.dataa(\registerArray[10][5]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[8][5]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux58~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~2 .lut_mask = 16'hCCB8;
defparam \Mux58~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N28
cycloneive_lcell_comb \Mux58~3 (
// Equation(s):
// \Mux58~3_combout  = (cuifregT_01 & ((\Mux58~2_combout  & (\registerArray[11][5]~q )) # (!\Mux58~2_combout  & ((\registerArray[9][5]~q ))))) # (!cuifregT_01 & (((\Mux58~2_combout ))))

	.dataa(\registerArray[11][5]~q ),
	.datab(\registerArray[9][5]~q ),
	.datac(cuifregT_0),
	.datad(\Mux58~2_combout ),
	.cin(gnd),
	.combout(\Mux58~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~3 .lut_mask = 16'hAFC0;
defparam \Mux58~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N2
cycloneive_lcell_comb \Mux58~6 (
// Equation(s):
// \Mux58~6_combout  = (cuifregT_2 & (cuifregT_3)) # (!cuifregT_2 & ((cuifregT_3 & ((\Mux58~3_combout ))) # (!cuifregT_3 & (\Mux58~5_combout ))))

	.dataa(cuifregT_2),
	.datab(cuifregT_3),
	.datac(\Mux58~5_combout ),
	.datad(\Mux58~3_combout ),
	.cin(gnd),
	.combout(\Mux58~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~6 .lut_mask = 16'hDC98;
defparam \Mux58~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N21
dffeas \registerArray[23][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][5] .is_wysiwyg = "true";
defparam \registerArray[23][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N11
dffeas \registerArray[27][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][5] .is_wysiwyg = "true";
defparam \registerArray[27][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N15
dffeas \registerArray[19][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][5] .is_wysiwyg = "true";
defparam \registerArray[19][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N14
cycloneive_lcell_comb \Mux58~17 (
// Equation(s):
// \Mux58~17_combout  = (cuifregT_3 & ((\registerArray[27][5]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[19][5]~q  & !cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[27][5]~q ),
	.datac(\registerArray[19][5]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux58~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~17 .lut_mask = 16'hAAD8;
defparam \Mux58~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y30_N1
dffeas \registerArray[31][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][5] .is_wysiwyg = "true";
defparam \registerArray[31][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N0
cycloneive_lcell_comb \Mux58~18 (
// Equation(s):
// \Mux58~18_combout  = (\Mux58~17_combout  & (((\registerArray[31][5]~q ) # (!cuifregT_2)))) # (!\Mux58~17_combout  & (\registerArray[23][5]~q  & ((cuifregT_2))))

	.dataa(\registerArray[23][5]~q ),
	.datab(\Mux58~17_combout ),
	.datac(\registerArray[31][5]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux58~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~18 .lut_mask = 16'hE2CC;
defparam \Mux58~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N8
cycloneive_lcell_comb \registerArray[28][5]~feeder (
// Equation(s):
// \registerArray[28][5]~feeder_combout  = \Mux63~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux632),
	.cin(gnd),
	.combout(\registerArray[28][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[28][5]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[28][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y31_N9
dffeas \registerArray[28][5] (
	.clk(clk),
	.d(\registerArray[28][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][5] .is_wysiwyg = "true";
defparam \registerArray[28][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N20
cycloneive_lcell_comb \registerArray[16][5]~feeder (
// Equation(s):
// \registerArray[16][5]~feeder_combout  = \Mux63~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux632),
	.cin(gnd),
	.combout(\registerArray[16][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[16][5]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[16][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y31_N21
dffeas \registerArray[16][5] (
	.clk(clk),
	.d(\registerArray[16][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][5] .is_wysiwyg = "true";
defparam \registerArray[16][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y43_N11
dffeas \registerArray[20][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][5] .is_wysiwyg = "true";
defparam \registerArray[20][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N14
cycloneive_lcell_comb \Mux58~14 (
// Equation(s):
// \Mux58~14_combout  = (cuifregT_2 & (((\registerArray[20][5]~q ) # (cuifregT_3)))) # (!cuifregT_2 & (\registerArray[16][5]~q  & ((!cuifregT_3))))

	.dataa(cuifregT_2),
	.datab(\registerArray[16][5]~q ),
	.datac(\registerArray[20][5]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux58~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~14 .lut_mask = 16'hAAE4;
defparam \Mux58~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N30
cycloneive_lcell_comb \Mux58~15 (
// Equation(s):
// \Mux58~15_combout  = (\Mux58~14_combout  & (((\registerArray[28][5]~q ) # (!cuifregT_3)))) # (!\Mux58~14_combout  & (\registerArray[24][5]~q  & ((cuifregT_3))))

	.dataa(\registerArray[24][5]~q ),
	.datab(\registerArray[28][5]~q ),
	.datac(\Mux58~14_combout ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux58~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~15 .lut_mask = 16'hCAF0;
defparam \Mux58~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N31
dffeas \registerArray[30][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][5] .is_wysiwyg = "true";
defparam \registerArray[30][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N21
dffeas \registerArray[18][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][5] .is_wysiwyg = "true";
defparam \registerArray[18][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N20
cycloneive_lcell_comb \Mux58~12 (
// Equation(s):
// \Mux58~12_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[22][5]~q )) # (!cuifregT_2 & ((\registerArray[18][5]~q )))))

	.dataa(\registerArray[22][5]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[18][5]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux58~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~12 .lut_mask = 16'hEE30;
defparam \Mux58~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N30
cycloneive_lcell_comb \Mux58~13 (
// Equation(s):
// \Mux58~13_combout  = (cuifregT_3 & ((\Mux58~12_combout  & ((\registerArray[30][5]~q ))) # (!\Mux58~12_combout  & (\registerArray[26][5]~q )))) # (!cuifregT_3 & (((\Mux58~12_combout ))))

	.dataa(\registerArray[26][5]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[30][5]~q ),
	.datad(\Mux58~12_combout ),
	.cin(gnd),
	.combout(\Mux58~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~13 .lut_mask = 16'hF388;
defparam \Mux58~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N4
cycloneive_lcell_comb \Mux58~16 (
// Equation(s):
// \Mux58~16_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & ((\Mux58~13_combout ))) # (!cuifregT_1 & (\Mux58~15_combout ))))

	.dataa(\Mux58~15_combout ),
	.datab(cuifregT_0),
	.datac(cuifregT_1),
	.datad(\Mux58~13_combout ),
	.cin(gnd),
	.combout(\Mux58~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~16 .lut_mask = 16'hF2C2;
defparam \Mux58~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y41_N1
dffeas \registerArray[21][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][5] .is_wysiwyg = "true";
defparam \registerArray[21][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N15
dffeas \registerArray[17][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][5] .is_wysiwyg = "true";
defparam \registerArray[17][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N14
cycloneive_lcell_comb \Mux58~10 (
// Equation(s):
// \Mux58~10_combout  = (cuifregT_3 & ((\registerArray[25][5]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[17][5]~q  & !cuifregT_2))))

	.dataa(\registerArray[25][5]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[17][5]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux58~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~10 .lut_mask = 16'hCCB8;
defparam \Mux58~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N25
dffeas \registerArray[29][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][5] .is_wysiwyg = "true";
defparam \registerArray[29][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N24
cycloneive_lcell_comb \Mux58~11 (
// Equation(s):
// \Mux58~11_combout  = (\Mux58~10_combout  & (((\registerArray[29][5]~q ) # (!cuifregT_2)))) # (!\Mux58~10_combout  & (\registerArray[21][5]~q  & ((cuifregT_2))))

	.dataa(\registerArray[21][5]~q ),
	.datab(\Mux58~10_combout ),
	.datac(\registerArray[29][5]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux58~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~11 .lut_mask = 16'hE2CC;
defparam \Mux58~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N20
cycloneive_lcell_comb \registerArray[15][19]~feeder (
// Equation(s):
// \registerArray[15][19]~feeder_combout  = \Mux49~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux492),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[15][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[15][19]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[15][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y32_N21
dffeas \registerArray[15][19] (
	.clk(clk),
	.d(\registerArray[15][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][19] .is_wysiwyg = "true";
defparam \registerArray[15][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N14
cycloneive_lcell_comb \registerArray[14][19]~feeder (
// Equation(s):
// \registerArray[14][19]~feeder_combout  = \Mux49~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux492),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[14][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][19]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[14][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y32_N15
dffeas \registerArray[14][19] (
	.clk(clk),
	.d(\registerArray[14][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][19] .is_wysiwyg = "true";
defparam \registerArray[14][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N29
dffeas \registerArray[12][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][19] .is_wysiwyg = "true";
defparam \registerArray[12][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N28
cycloneive_lcell_comb \Mux44~7 (
// Equation(s):
// \Mux44~7_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[13][19]~q )) # (!cuifregT_01 & ((\registerArray[12][19]~q )))))

	.dataa(\registerArray[13][19]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[12][19]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux44~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~7 .lut_mask = 16'hEE30;
defparam \Mux44~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N10
cycloneive_lcell_comb \Mux44~8 (
// Equation(s):
// \Mux44~8_combout  = (cuifregT_1 & ((\Mux44~7_combout  & (\registerArray[15][19]~q )) # (!\Mux44~7_combout  & ((\registerArray[14][19]~q ))))) # (!cuifregT_1 & (((\Mux44~7_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[15][19]~q ),
	.datac(\registerArray[14][19]~q ),
	.datad(\Mux44~7_combout ),
	.cin(gnd),
	.combout(\Mux44~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~8 .lut_mask = 16'hDDA0;
defparam \Mux44~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N11
dffeas \registerArray[6][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][19] .is_wysiwyg = "true";
defparam \registerArray[6][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N9
dffeas \registerArray[7][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][19] .is_wysiwyg = "true";
defparam \registerArray[7][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N11
dffeas \registerArray[4][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][19] .is_wysiwyg = "true";
defparam \registerArray[4][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N10
cycloneive_lcell_comb \Mux44~0 (
// Equation(s):
// \Mux44~0_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[5][19]~q )) # (!cuifregT_01 & ((\registerArray[4][19]~q )))))

	.dataa(\registerArray[5][19]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[4][19]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux44~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~0 .lut_mask = 16'hEE30;
defparam \Mux44~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N8
cycloneive_lcell_comb \Mux44~1 (
// Equation(s):
// \Mux44~1_combout  = (cuifregT_1 & ((\Mux44~0_combout  & ((\registerArray[7][19]~q ))) # (!\Mux44~0_combout  & (\registerArray[6][19]~q )))) # (!cuifregT_1 & (((\Mux44~0_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[6][19]~q ),
	.datac(\registerArray[7][19]~q ),
	.datad(\Mux44~0_combout ),
	.cin(gnd),
	.combout(\Mux44~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~1 .lut_mask = 16'hF588;
defparam \Mux44~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y42_N15
dffeas \registerArray[11][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][19] .is_wysiwyg = "true";
defparam \registerArray[11][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N10
cycloneive_lcell_comb \registerArray[8][19]~feeder (
// Equation(s):
// \registerArray[8][19]~feeder_combout  = \Mux49~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux492),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[8][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[8][19]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[8][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y43_N11
dffeas \registerArray[8][19] (
	.clk(clk),
	.d(\registerArray[8][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][19] .is_wysiwyg = "true";
defparam \registerArray[8][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N16
cycloneive_lcell_comb \Mux44~2 (
// Equation(s):
// \Mux44~2_combout  = (cuifregT_1 & ((\registerArray[10][19]~q ) # ((cuifregT_01)))) # (!cuifregT_1 & (((\registerArray[8][19]~q  & !cuifregT_01))))

	.dataa(\registerArray[10][19]~q ),
	.datab(\registerArray[8][19]~q ),
	.datac(cuifregT_1),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux44~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~2 .lut_mask = 16'hF0AC;
defparam \Mux44~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N14
cycloneive_lcell_comb \Mux44~3 (
// Equation(s):
// \Mux44~3_combout  = (cuifregT_01 & ((\Mux44~2_combout  & ((\registerArray[11][19]~q ))) # (!\Mux44~2_combout  & (\registerArray[9][19]~q )))) # (!cuifregT_01 & (((\Mux44~2_combout ))))

	.dataa(\registerArray[9][19]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[11][19]~q ),
	.datad(\Mux44~2_combout ),
	.cin(gnd),
	.combout(\Mux44~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~3 .lut_mask = 16'hF388;
defparam \Mux44~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y42_N29
dffeas \registerArray[2][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][19] .is_wysiwyg = "true";
defparam \registerArray[2][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N25
dffeas \registerArray[3][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][19] .is_wysiwyg = "true";
defparam \registerArray[3][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N24
cycloneive_lcell_comb \Mux44~4 (
// Equation(s):
// \Mux44~4_combout  = (cuifregT_01 & ((cuifregT_1 & ((\registerArray[3][19]~q ))) # (!cuifregT_1 & (\registerArray[1][19]~q ))))

	.dataa(\registerArray[1][19]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[3][19]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux44~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~4 .lut_mask = 16'hC088;
defparam \Mux44~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N28
cycloneive_lcell_comb \Mux44~5 (
// Equation(s):
// \Mux44~5_combout  = (\Mux44~4_combout ) # ((!cuifregT_01 & (cuifregT_1 & \registerArray[2][19]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[2][19]~q ),
	.datad(\Mux44~4_combout ),
	.cin(gnd),
	.combout(\Mux44~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~5 .lut_mask = 16'hFF40;
defparam \Mux44~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N12
cycloneive_lcell_comb \Mux44~6 (
// Equation(s):
// \Mux44~6_combout  = (cuifregT_2 & (cuifregT_3)) # (!cuifregT_2 & ((cuifregT_3 & (\Mux44~3_combout )) # (!cuifregT_3 & ((\Mux44~5_combout )))))

	.dataa(cuifregT_2),
	.datab(cuifregT_3),
	.datac(\Mux44~3_combout ),
	.datad(\Mux44~5_combout ),
	.cin(gnd),
	.combout(\Mux44~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~6 .lut_mask = 16'hD9C8;
defparam \Mux44~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N27
dffeas \registerArray[28][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][19] .is_wysiwyg = "true";
defparam \registerArray[28][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N29
dffeas \registerArray[16][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][19] .is_wysiwyg = "true";
defparam \registerArray[16][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N28
cycloneive_lcell_comb \Mux44~14 (
// Equation(s):
// \Mux44~14_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[20][19]~q )) # (!cuifregT_2 & ((\registerArray[16][19]~q )))))

	.dataa(\registerArray[20][19]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[16][19]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux44~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~14 .lut_mask = 16'hEE30;
defparam \Mux44~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N26
cycloneive_lcell_comb \Mux44~15 (
// Equation(s):
// \Mux44~15_combout  = (cuifregT_3 & ((\Mux44~14_combout  & ((\registerArray[28][19]~q ))) # (!\Mux44~14_combout  & (\registerArray[24][19]~q )))) # (!cuifregT_3 & (((\Mux44~14_combout ))))

	.dataa(\registerArray[24][19]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[28][19]~q ),
	.datad(\Mux44~14_combout ),
	.cin(gnd),
	.combout(\Mux44~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~15 .lut_mask = 16'hF388;
defparam \Mux44~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N24
cycloneive_lcell_comb \registerArray[26][19]~feeder (
// Equation(s):
// \registerArray[26][19]~feeder_combout  = \Mux49~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux492),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[26][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[26][19]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[26][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N25
dffeas \registerArray[26][19] (
	.clk(clk),
	.d(\registerArray[26][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][19] .is_wysiwyg = "true";
defparam \registerArray[26][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N15
dffeas \registerArray[30][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][19] .is_wysiwyg = "true";
defparam \registerArray[30][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N30
cycloneive_lcell_comb \registerArray[22][19]~feeder (
// Equation(s):
// \registerArray[22][19]~feeder_combout  = \Mux49~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux492),
	.cin(gnd),
	.combout(\registerArray[22][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[22][19]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[22][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y40_N31
dffeas \registerArray[22][19] (
	.clk(clk),
	.d(\registerArray[22][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][19] .is_wysiwyg = "true";
defparam \registerArray[22][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N25
dffeas \registerArray[18][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][19] .is_wysiwyg = "true";
defparam \registerArray[18][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N24
cycloneive_lcell_comb \Mux44~12 (
// Equation(s):
// \Mux44~12_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[22][19]~q )) # (!cuifregT_2 & ((\registerArray[18][19]~q )))))

	.dataa(cuifregT_3),
	.datab(\registerArray[22][19]~q ),
	.datac(\registerArray[18][19]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux44~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~12 .lut_mask = 16'hEE50;
defparam \Mux44~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N14
cycloneive_lcell_comb \Mux44~13 (
// Equation(s):
// \Mux44~13_combout  = (cuifregT_3 & ((\Mux44~12_combout  & ((\registerArray[30][19]~q ))) # (!\Mux44~12_combout  & (\registerArray[26][19]~q )))) # (!cuifregT_3 & (((\Mux44~12_combout ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[26][19]~q ),
	.datac(\registerArray[30][19]~q ),
	.datad(\Mux44~12_combout ),
	.cin(gnd),
	.combout(\Mux44~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~13 .lut_mask = 16'hF588;
defparam \Mux44~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N8
cycloneive_lcell_comb \Mux44~16 (
// Equation(s):
// \Mux44~16_combout  = (cuifregT_1 & ((cuifregT_01) # ((\Mux44~13_combout )))) # (!cuifregT_1 & (!cuifregT_01 & (\Mux44~15_combout )))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\Mux44~15_combout ),
	.datad(\Mux44~13_combout ),
	.cin(gnd),
	.combout(\Mux44~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~16 .lut_mask = 16'hBA98;
defparam \Mux44~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N13
dffeas \registerArray[23][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][19] .is_wysiwyg = "true";
defparam \registerArray[23][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N13
dffeas \registerArray[31][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][19] .is_wysiwyg = "true";
defparam \registerArray[31][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N15
dffeas \registerArray[27][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][19] .is_wysiwyg = "true";
defparam \registerArray[27][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N3
dffeas \registerArray[19][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][19] .is_wysiwyg = "true";
defparam \registerArray[19][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N2
cycloneive_lcell_comb \Mux44~17 (
// Equation(s):
// \Mux44~17_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[27][19]~q )) # (!cuifregT_3 & ((\registerArray[19][19]~q )))))

	.dataa(cuifregT_2),
	.datab(\registerArray[27][19]~q ),
	.datac(\registerArray[19][19]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux44~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~17 .lut_mask = 16'hEE50;
defparam \Mux44~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N12
cycloneive_lcell_comb \Mux44~18 (
// Equation(s):
// \Mux44~18_combout  = (cuifregT_2 & ((\Mux44~17_combout  & ((\registerArray[31][19]~q ))) # (!\Mux44~17_combout  & (\registerArray[23][19]~q )))) # (!cuifregT_2 & (((\Mux44~17_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[23][19]~q ),
	.datac(\registerArray[31][19]~q ),
	.datad(\Mux44~17_combout ),
	.cin(gnd),
	.combout(\Mux44~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~18 .lut_mask = 16'hF588;
defparam \Mux44~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N25
dffeas \registerArray[21][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][19] .is_wysiwyg = "true";
defparam \registerArray[21][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y31_N19
dffeas \registerArray[29][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][19] .is_wysiwyg = "true";
defparam \registerArray[29][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N8
cycloneive_lcell_comb \registerArray[25][19]~feeder (
// Equation(s):
// \registerArray[25][19]~feeder_combout  = \Mux49~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux492),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[25][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[25][19]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[25][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N9
dffeas \registerArray[25][19] (
	.clk(clk),
	.d(\registerArray[25][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][19] .is_wysiwyg = "true";
defparam \registerArray[25][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N27
dffeas \registerArray[17][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][19] .is_wysiwyg = "true";
defparam \registerArray[17][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N26
cycloneive_lcell_comb \Mux44~10 (
// Equation(s):
// \Mux44~10_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[25][19]~q )) # (!cuifregT_3 & ((\registerArray[17][19]~q )))))

	.dataa(cuifregT_2),
	.datab(\registerArray[25][19]~q ),
	.datac(\registerArray[17][19]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux44~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~10 .lut_mask = 16'hEE50;
defparam \Mux44~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N18
cycloneive_lcell_comb \Mux44~11 (
// Equation(s):
// \Mux44~11_combout  = (cuifregT_2 & ((\Mux44~10_combout  & ((\registerArray[29][19]~q ))) # (!\Mux44~10_combout  & (\registerArray[21][19]~q )))) # (!cuifregT_2 & (((\Mux44~10_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[21][19]~q ),
	.datac(\registerArray[29][19]~q ),
	.datad(\Mux44~10_combout ),
	.cin(gnd),
	.combout(\Mux44~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~11 .lut_mask = 16'hF588;
defparam \Mux44~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N16
cycloneive_lcell_comb \registerArray[9][18]~feeder (
// Equation(s):
// \registerArray[9][18]~feeder_combout  = \Mux50~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux502),
	.cin(gnd),
	.combout(\registerArray[9][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[9][18]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[9][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y41_N17
dffeas \registerArray[9][18] (
	.clk(clk),
	.d(\registerArray[9][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][18] .is_wysiwyg = "true";
defparam \registerArray[9][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N31
dffeas \registerArray[11][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][18] .is_wysiwyg = "true";
defparam \registerArray[11][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N25
dffeas \registerArray[8][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][18] .is_wysiwyg = "true";
defparam \registerArray[8][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N24
cycloneive_lcell_comb \Mux45~0 (
// Equation(s):
// \Mux45~0_combout  = (cuifregT_1 & ((\registerArray[10][18]~q ) # ((cuifregT_01)))) # (!cuifregT_1 & (((\registerArray[8][18]~q  & !cuifregT_01))))

	.dataa(\registerArray[10][18]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[8][18]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux45~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~0 .lut_mask = 16'hCCB8;
defparam \Mux45~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N30
cycloneive_lcell_comb \Mux45~1 (
// Equation(s):
// \Mux45~1_combout  = (cuifregT_01 & ((\Mux45~0_combout  & ((\registerArray[11][18]~q ))) # (!\Mux45~0_combout  & (\registerArray[9][18]~q )))) # (!cuifregT_01 & (((\Mux45~0_combout ))))

	.dataa(\registerArray[9][18]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[11][18]~q ),
	.datad(\Mux45~0_combout ),
	.cin(gnd),
	.combout(\Mux45~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~1 .lut_mask = 16'hF388;
defparam \Mux45~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N4
cycloneive_lcell_comb \registerArray[14][18]~feeder (
// Equation(s):
// \registerArray[14][18]~feeder_combout  = \Mux50~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux502),
	.cin(gnd),
	.combout(\registerArray[14][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][18]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[14][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y42_N5
dffeas \registerArray[14][18] (
	.clk(clk),
	.d(\registerArray[14][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][18] .is_wysiwyg = "true";
defparam \registerArray[14][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N17
dffeas \registerArray[15][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][18] .is_wysiwyg = "true";
defparam \registerArray[15][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N7
dffeas \registerArray[12][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][18] .is_wysiwyg = "true";
defparam \registerArray[12][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N6
cycloneive_lcell_comb \Mux45~7 (
// Equation(s):
// \Mux45~7_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[13][18]~q )) # (!cuifregT_01 & ((\registerArray[12][18]~q )))))

	.dataa(\registerArray[13][18]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[12][18]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux45~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~7 .lut_mask = 16'hEE30;
defparam \Mux45~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N16
cycloneive_lcell_comb \Mux45~8 (
// Equation(s):
// \Mux45~8_combout  = (cuifregT_1 & ((\Mux45~7_combout  & ((\registerArray[15][18]~q ))) # (!\Mux45~7_combout  & (\registerArray[14][18]~q )))) # (!cuifregT_1 & (((\Mux45~7_combout ))))

	.dataa(\registerArray[14][18]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[15][18]~q ),
	.datad(\Mux45~7_combout ),
	.cin(gnd),
	.combout(\Mux45~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~8 .lut_mask = 16'hF388;
defparam \Mux45~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y31_N13
dffeas \registerArray[7][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][18] .is_wysiwyg = "true";
defparam \registerArray[7][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N19
dffeas \registerArray[4][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][18] .is_wysiwyg = "true";
defparam \registerArray[4][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N18
cycloneive_lcell_comb \Mux45~2 (
// Equation(s):
// \Mux45~2_combout  = (cuifregT_01 & ((\registerArray[5][18]~q ) # ((cuifregT_1)))) # (!cuifregT_01 & (((\registerArray[4][18]~q  & !cuifregT_1))))

	.dataa(\registerArray[5][18]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[4][18]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux45~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~2 .lut_mask = 16'hCCB8;
defparam \Mux45~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N12
cycloneive_lcell_comb \Mux45~3 (
// Equation(s):
// \Mux45~3_combout  = (cuifregT_1 & ((\Mux45~2_combout  & ((\registerArray[7][18]~q ))) # (!\Mux45~2_combout  & (\registerArray[6][18]~q )))) # (!cuifregT_1 & (((\Mux45~2_combout ))))

	.dataa(\registerArray[6][18]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[7][18]~q ),
	.datad(\Mux45~2_combout ),
	.cin(gnd),
	.combout(\Mux45~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~3 .lut_mask = 16'hF388;
defparam \Mux45~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y42_N7
dffeas \registerArray[1][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][18] .is_wysiwyg = "true";
defparam \registerArray[1][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N6
cycloneive_lcell_comb \Mux45~4 (
// Equation(s):
// \Mux45~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][18]~q )) # (!cuifregT_1 & ((\registerArray[1][18]~q )))))

	.dataa(\registerArray[3][18]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[1][18]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux45~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~4 .lut_mask = 16'hB800;
defparam \Mux45~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N24
cycloneive_lcell_comb \Mux45~5 (
// Equation(s):
// \Mux45~5_combout  = (\Mux45~4_combout ) # ((\registerArray[2][18]~q  & (!cuifregT_01 & cuifregT_1)))

	.dataa(\registerArray[2][18]~q ),
	.datab(cuifregT_0),
	.datac(cuifregT_1),
	.datad(\Mux45~4_combout ),
	.cin(gnd),
	.combout(\Mux45~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~5 .lut_mask = 16'hFF20;
defparam \Mux45~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y34_N6
cycloneive_lcell_comb \Mux45~6 (
// Equation(s):
// \Mux45~6_combout  = (cuifregT_2 & ((cuifregT_3) # ((\Mux45~3_combout )))) # (!cuifregT_2 & (!cuifregT_3 & ((\Mux45~5_combout ))))

	.dataa(cuifregT_2),
	.datab(cuifregT_3),
	.datac(\Mux45~3_combout ),
	.datad(\Mux45~5_combout ),
	.cin(gnd),
	.combout(\Mux45~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~6 .lut_mask = 16'hB9A8;
defparam \Mux45~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N15
dffeas \registerArray[22][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][18] .is_wysiwyg = "true";
defparam \registerArray[22][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N19
dffeas \registerArray[30][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][18] .is_wysiwyg = "true";
defparam \registerArray[30][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y33_N25
dffeas \registerArray[18][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][18] .is_wysiwyg = "true";
defparam \registerArray[18][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N24
cycloneive_lcell_comb \Mux45~12 (
// Equation(s):
// \Mux45~12_combout  = (cuifregT_3 & ((\registerArray[26][18]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[18][18]~q  & !cuifregT_2))))

	.dataa(\registerArray[26][18]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[18][18]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux45~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~12 .lut_mask = 16'hCCB8;
defparam \Mux45~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N18
cycloneive_lcell_comb \Mux45~13 (
// Equation(s):
// \Mux45~13_combout  = (cuifregT_2 & ((\Mux45~12_combout  & ((\registerArray[30][18]~q ))) # (!\Mux45~12_combout  & (\registerArray[22][18]~q )))) # (!cuifregT_2 & (((\Mux45~12_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[22][18]~q ),
	.datac(\registerArray[30][18]~q ),
	.datad(\Mux45~12_combout ),
	.cin(gnd),
	.combout(\Mux45~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~13 .lut_mask = 16'hF588;
defparam \Mux45~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y33_N3
dffeas \registerArray[28][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][18] .is_wysiwyg = "true";
defparam \registerArray[28][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y41_N3
dffeas \registerArray[24][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][18] .is_wysiwyg = "true";
defparam \registerArray[24][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N13
dffeas \registerArray[16][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][18] .is_wysiwyg = "true";
defparam \registerArray[16][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N12
cycloneive_lcell_comb \Mux45~14 (
// Equation(s):
// \Mux45~14_combout  = (cuifregT_3 & ((\registerArray[24][18]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[16][18]~q  & !cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[24][18]~q ),
	.datac(\registerArray[16][18]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux45~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~14 .lut_mask = 16'hAAD8;
defparam \Mux45~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N2
cycloneive_lcell_comb \Mux45~15 (
// Equation(s):
// \Mux45~15_combout  = (cuifregT_2 & ((\Mux45~14_combout  & ((\registerArray[28][18]~q ))) # (!\Mux45~14_combout  & (\registerArray[20][18]~q )))) # (!cuifregT_2 & (((\Mux45~14_combout ))))

	.dataa(\registerArray[20][18]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[28][18]~q ),
	.datad(\Mux45~14_combout ),
	.cin(gnd),
	.combout(\Mux45~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~15 .lut_mask = 16'hF388;
defparam \Mux45~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N16
cycloneive_lcell_comb \Mux45~16 (
// Equation(s):
// \Mux45~16_combout  = (cuifregT_1 & ((cuifregT_01) # ((\Mux45~13_combout )))) # (!cuifregT_1 & (!cuifregT_01 & ((\Mux45~15_combout ))))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\Mux45~13_combout ),
	.datad(\Mux45~15_combout ),
	.cin(gnd),
	.combout(\Mux45~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~16 .lut_mask = 16'hB9A8;
defparam \Mux45~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N6
cycloneive_lcell_comb \registerArray[27][18]~feeder (
// Equation(s):
// \registerArray[27][18]~feeder_combout  = \Mux50~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux502),
	.cin(gnd),
	.combout(\registerArray[27][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[27][18]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[27][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N7
dffeas \registerArray[27][18] (
	.clk(clk),
	.d(\registerArray[27][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][18] .is_wysiwyg = "true";
defparam \registerArray[27][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N7
dffeas \registerArray[31][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][18] .is_wysiwyg = "true";
defparam \registerArray[31][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N1
dffeas \registerArray[19][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][18] .is_wysiwyg = "true";
defparam \registerArray[19][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N0
cycloneive_lcell_comb \Mux45~17 (
// Equation(s):
// \Mux45~17_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[23][18]~q )) # (!cuifregT_2 & ((\registerArray[19][18]~q )))))

	.dataa(\registerArray[23][18]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[19][18]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux45~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~17 .lut_mask = 16'hEE30;
defparam \Mux45~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N6
cycloneive_lcell_comb \Mux45~18 (
// Equation(s):
// \Mux45~18_combout  = (cuifregT_3 & ((\Mux45~17_combout  & ((\registerArray[31][18]~q ))) # (!\Mux45~17_combout  & (\registerArray[27][18]~q )))) # (!cuifregT_3 & (((\Mux45~17_combout ))))

	.dataa(\registerArray[27][18]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[31][18]~q ),
	.datad(\Mux45~17_combout ),
	.cin(gnd),
	.combout(\Mux45~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~18 .lut_mask = 16'hF388;
defparam \Mux45~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N28
cycloneive_lcell_comb \registerArray[25][18]~feeder (
// Equation(s):
// \registerArray[25][18]~feeder_combout  = \Mux50~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux502),
	.cin(gnd),
	.combout(\registerArray[25][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[25][18]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[25][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y41_N29
dffeas \registerArray[25][18] (
	.clk(clk),
	.d(\registerArray[25][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][18] .is_wysiwyg = "true";
defparam \registerArray[25][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N11
dffeas \registerArray[29][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][18] .is_wysiwyg = "true";
defparam \registerArray[29][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N18
cycloneive_lcell_comb \registerArray[21][18]~feeder (
// Equation(s):
// \registerArray[21][18]~feeder_combout  = \Mux50~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux502),
	.cin(gnd),
	.combout(\registerArray[21][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[21][18]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[21][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y41_N19
dffeas \registerArray[21][18] (
	.clk(clk),
	.d(\registerArray[21][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][18] .is_wysiwyg = "true";
defparam \registerArray[21][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N28
cycloneive_lcell_comb \Mux45~10 (
// Equation(s):
// \Mux45~10_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & ((\registerArray[21][18]~q ))) # (!cuifregT_2 & (\registerArray[17][18]~q ))))

	.dataa(\registerArray[17][18]~q ),
	.datab(\registerArray[21][18]~q ),
	.datac(cuifregT_3),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux45~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~10 .lut_mask = 16'hFC0A;
defparam \Mux45~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N10
cycloneive_lcell_comb \Mux45~11 (
// Equation(s):
// \Mux45~11_combout  = (cuifregT_3 & ((\Mux45~10_combout  & ((\registerArray[29][18]~q ))) # (!\Mux45~10_combout  & (\registerArray[25][18]~q )))) # (!cuifregT_3 & (((\Mux45~10_combout ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[25][18]~q ),
	.datac(\registerArray[29][18]~q ),
	.datad(\Mux45~10_combout ),
	.cin(gnd),
	.combout(\Mux45~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~11 .lut_mask = 16'hF588;
defparam \Mux45~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N16
cycloneive_lcell_comb \registerArray[14][17]~feeder (
// Equation(s):
// \registerArray[14][17]~feeder_combout  = \Mux51~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux512),
	.cin(gnd),
	.combout(\registerArray[14][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][17]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[14][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N17
dffeas \registerArray[14][17] (
	.clk(clk),
	.d(\registerArray[14][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][17] .is_wysiwyg = "true";
defparam \registerArray[14][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N9
dffeas \registerArray[15][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][17] .is_wysiwyg = "true";
defparam \registerArray[15][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N19
dffeas \registerArray[12][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][17] .is_wysiwyg = "true";
defparam \registerArray[12][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N18
cycloneive_lcell_comb \Mux46~7 (
// Equation(s):
// \Mux46~7_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[13][17]~q )) # (!cuifregT_01 & ((\registerArray[12][17]~q )))))

	.dataa(\registerArray[13][17]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[12][17]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux46~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~7 .lut_mask = 16'hEE30;
defparam \Mux46~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N8
cycloneive_lcell_comb \Mux46~8 (
// Equation(s):
// \Mux46~8_combout  = (cuifregT_1 & ((\Mux46~7_combout  & ((\registerArray[15][17]~q ))) # (!\Mux46~7_combout  & (\registerArray[14][17]~q )))) # (!cuifregT_1 & (((\Mux46~7_combout ))))

	.dataa(\registerArray[14][17]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[15][17]~q ),
	.datad(\Mux46~7_combout ),
	.cin(gnd),
	.combout(\Mux46~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~8 .lut_mask = 16'hF388;
defparam \Mux46~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N25
dffeas \registerArray[6][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][17] .is_wysiwyg = "true";
defparam \registerArray[6][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N27
dffeas \registerArray[7][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][17] .is_wysiwyg = "true";
defparam \registerArray[7][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N5
dffeas \registerArray[5][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][17] .is_wysiwyg = "true";
defparam \registerArray[5][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N12
cycloneive_lcell_comb \Mux46~0 (
// Equation(s):
// \Mux46~0_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & ((\registerArray[5][17]~q ))) # (!cuifregT_01 & (\registerArray[4][17]~q ))))

	.dataa(\registerArray[4][17]~q ),
	.datab(\registerArray[5][17]~q ),
	.datac(cuifregT_1),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux46~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~0 .lut_mask = 16'hFC0A;
defparam \Mux46~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N26
cycloneive_lcell_comb \Mux46~1 (
// Equation(s):
// \Mux46~1_combout  = (cuifregT_1 & ((\Mux46~0_combout  & ((\registerArray[7][17]~q ))) # (!\Mux46~0_combout  & (\registerArray[6][17]~q )))) # (!cuifregT_1 & (((\Mux46~0_combout ))))

	.dataa(\registerArray[6][17]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[7][17]~q ),
	.datad(\Mux46~0_combout ),
	.cin(gnd),
	.combout(\Mux46~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~1 .lut_mask = 16'hF388;
defparam \Mux46~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N5
dffeas \registerArray[9][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][17] .is_wysiwyg = "true";
defparam \registerArray[9][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N19
dffeas \registerArray[11][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][17] .is_wysiwyg = "true";
defparam \registerArray[11][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N17
dffeas \registerArray[8][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][17] .is_wysiwyg = "true";
defparam \registerArray[8][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N16
cycloneive_lcell_comb \Mux46~2 (
// Equation(s):
// \Mux46~2_combout  = (cuifregT_1 & ((\registerArray[10][17]~q ) # ((cuifregT_01)))) # (!cuifregT_1 & (((\registerArray[8][17]~q  & !cuifregT_01))))

	.dataa(\registerArray[10][17]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[8][17]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux46~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~2 .lut_mask = 16'hCCB8;
defparam \Mux46~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N18
cycloneive_lcell_comb \Mux46~3 (
// Equation(s):
// \Mux46~3_combout  = (cuifregT_01 & ((\Mux46~2_combout  & ((\registerArray[11][17]~q ))) # (!\Mux46~2_combout  & (\registerArray[9][17]~q )))) # (!cuifregT_01 & (((\Mux46~2_combout ))))

	.dataa(cuifregT_0),
	.datab(\registerArray[9][17]~q ),
	.datac(\registerArray[11][17]~q ),
	.datad(\Mux46~2_combout ),
	.cin(gnd),
	.combout(\Mux46~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~3 .lut_mask = 16'hF588;
defparam \Mux46~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y40_N7
dffeas \registerArray[2][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][17] .is_wysiwyg = "true";
defparam \registerArray[2][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y40_N25
dffeas \registerArray[1][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][17] .is_wysiwyg = "true";
defparam \registerArray[1][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N24
cycloneive_lcell_comb \Mux46~4 (
// Equation(s):
// \Mux46~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][17]~q )) # (!cuifregT_1 & ((\registerArray[1][17]~q )))))

	.dataa(\registerArray[3][17]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[1][17]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux46~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~4 .lut_mask = 16'hB800;
defparam \Mux46~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N6
cycloneive_lcell_comb \Mux46~5 (
// Equation(s):
// \Mux46~5_combout  = (\Mux46~4_combout ) # ((!cuifregT_01 & (cuifregT_1 & \registerArray[2][17]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[2][17]~q ),
	.datad(\Mux46~4_combout ),
	.cin(gnd),
	.combout(\Mux46~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~5 .lut_mask = 16'hFF40;
defparam \Mux46~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N14
cycloneive_lcell_comb \Mux46~6 (
// Equation(s):
// \Mux46~6_combout  = (cuifregT_2 & (cuifregT_3)) # (!cuifregT_2 & ((cuifregT_3 & (\Mux46~3_combout )) # (!cuifregT_3 & ((\Mux46~5_combout )))))

	.dataa(cuifregT_2),
	.datab(cuifregT_3),
	.datac(\Mux46~3_combout ),
	.datad(\Mux46~5_combout ),
	.cin(gnd),
	.combout(\Mux46~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~6 .lut_mask = 16'hD9C8;
defparam \Mux46~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N11
dffeas \registerArray[24][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][17] .is_wysiwyg = "true";
defparam \registerArray[24][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N15
dffeas \registerArray[28][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][17] .is_wysiwyg = "true";
defparam \registerArray[28][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N21
dffeas \registerArray[16][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][17] .is_wysiwyg = "true";
defparam \registerArray[16][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N20
cycloneive_lcell_comb \Mux46~14 (
// Equation(s):
// \Mux46~14_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[20][17]~q )) # (!cuifregT_2 & ((\registerArray[16][17]~q )))))

	.dataa(\registerArray[20][17]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[16][17]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux46~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~14 .lut_mask = 16'hEE30;
defparam \Mux46~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N14
cycloneive_lcell_comb \Mux46~15 (
// Equation(s):
// \Mux46~15_combout  = (cuifregT_3 & ((\Mux46~14_combout  & ((\registerArray[28][17]~q ))) # (!\Mux46~14_combout  & (\registerArray[24][17]~q )))) # (!cuifregT_3 & (((\Mux46~14_combout ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[24][17]~q ),
	.datac(\registerArray[28][17]~q ),
	.datad(\Mux46~14_combout ),
	.cin(gnd),
	.combout(\Mux46~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~15 .lut_mask = 16'hF588;
defparam \Mux46~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N11
dffeas \registerArray[30][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][17] .is_wysiwyg = "true";
defparam \registerArray[30][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N29
dffeas \registerArray[18][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][17] .is_wysiwyg = "true";
defparam \registerArray[18][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N28
cycloneive_lcell_comb \Mux46~12 (
// Equation(s):
// \Mux46~12_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[22][17]~q )) # (!cuifregT_2 & ((\registerArray[18][17]~q )))))

	.dataa(\registerArray[22][17]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[18][17]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux46~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~12 .lut_mask = 16'hEE30;
defparam \Mux46~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N10
cycloneive_lcell_comb \Mux46~13 (
// Equation(s):
// \Mux46~13_combout  = (cuifregT_3 & ((\Mux46~12_combout  & ((\registerArray[30][17]~q ))) # (!\Mux46~12_combout  & (\registerArray[26][17]~q )))) # (!cuifregT_3 & (((\Mux46~12_combout ))))

	.dataa(\registerArray[26][17]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[30][17]~q ),
	.datad(\Mux46~12_combout ),
	.cin(gnd),
	.combout(\Mux46~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~13 .lut_mask = 16'hF388;
defparam \Mux46~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N0
cycloneive_lcell_comb \Mux46~16 (
// Equation(s):
// \Mux46~16_combout  = (cuifregT_1 & ((cuifregT_01) # ((\Mux46~13_combout )))) # (!cuifregT_1 & (!cuifregT_01 & (\Mux46~15_combout )))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\Mux46~15_combout ),
	.datad(\Mux46~13_combout ),
	.cin(gnd),
	.combout(\Mux46~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~16 .lut_mask = 16'hBA98;
defparam \Mux46~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y41_N25
dffeas \registerArray[21][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][17] .is_wysiwyg = "true";
defparam \registerArray[21][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y37_N3
dffeas \registerArray[29][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][17] .is_wysiwyg = "true";
defparam \registerArray[29][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y41_N7
dffeas \registerArray[25][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][17] .is_wysiwyg = "true";
defparam \registerArray[25][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N0
cycloneive_lcell_comb \Mux46~10 (
// Equation(s):
// \Mux46~10_combout  = (cuifregT_3 & (((\registerArray[25][17]~q ) # (cuifregT_2)))) # (!cuifregT_3 & (\registerArray[17][17]~q  & ((!cuifregT_2))))

	.dataa(\registerArray[17][17]~q ),
	.datab(\registerArray[25][17]~q ),
	.datac(cuifregT_3),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux46~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~10 .lut_mask = 16'hF0CA;
defparam \Mux46~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N2
cycloneive_lcell_comb \Mux46~11 (
// Equation(s):
// \Mux46~11_combout  = (cuifregT_2 & ((\Mux46~10_combout  & ((\registerArray[29][17]~q ))) # (!\Mux46~10_combout  & (\registerArray[21][17]~q )))) # (!cuifregT_2 & (((\Mux46~10_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[21][17]~q ),
	.datac(\registerArray[29][17]~q ),
	.datad(\Mux46~10_combout ),
	.cin(gnd),
	.combout(\Mux46~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~11 .lut_mask = 16'hF588;
defparam \Mux46~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y37_N31
dffeas \registerArray[31][17] (
	.clk(clk),
	.d(Mux512),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][17] .is_wysiwyg = "true";
defparam \registerArray[31][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N15
dffeas \registerArray[23][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][17] .is_wysiwyg = "true";
defparam \registerArray[23][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y41_N5
dffeas \registerArray[19][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][17] .is_wysiwyg = "true";
defparam \registerArray[19][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N4
cycloneive_lcell_comb \Mux46~17 (
// Equation(s):
// \Mux46~17_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[27][17]~q )) # (!cuifregT_3 & ((\registerArray[19][17]~q )))))

	.dataa(\registerArray[27][17]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[19][17]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux46~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~17 .lut_mask = 16'hEE30;
defparam \Mux46~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N14
cycloneive_lcell_comb \Mux46~18 (
// Equation(s):
// \Mux46~18_combout  = (cuifregT_2 & ((\Mux46~17_combout  & (\registerArray[31][17]~q )) # (!\Mux46~17_combout  & ((\registerArray[23][17]~q ))))) # (!cuifregT_2 & (((\Mux46~17_combout ))))

	.dataa(\registerArray[31][17]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[23][17]~q ),
	.datad(\Mux46~17_combout ),
	.cin(gnd),
	.combout(\Mux46~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~18 .lut_mask = 16'hBBC0;
defparam \Mux46~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N28
cycloneive_lcell_comb \registerArray[27][16]~feeder (
// Equation(s):
// \registerArray[27][16]~feeder_combout  = \Mux52~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux522),
	.cin(gnd),
	.combout(\registerArray[27][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[27][16]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[27][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y40_N29
dffeas \registerArray[27][16] (
	.clk(clk),
	.d(\registerArray[27][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][16] .is_wysiwyg = "true";
defparam \registerArray[27][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N17
dffeas \registerArray[31][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][16] .is_wysiwyg = "true";
defparam \registerArray[31][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N20
cycloneive_lcell_comb \registerArray[19][16]~feeder (
// Equation(s):
// \registerArray[19][16]~feeder_combout  = \Mux52~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux522),
	.cin(gnd),
	.combout(\registerArray[19][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[19][16]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[19][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y31_N21
dffeas \registerArray[19][16] (
	.clk(clk),
	.d(\registerArray[19][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][16] .is_wysiwyg = "true";
defparam \registerArray[19][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N10
cycloneive_lcell_comb \Mux47~7 (
// Equation(s):
// \Mux47~7_combout  = (cuifregT_2 & ((\registerArray[23][16]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[19][16]~q  & !cuifregT_3))))

	.dataa(\registerArray[23][16]~q ),
	.datab(\registerArray[19][16]~q ),
	.datac(cuifregT_2),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux47~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~7 .lut_mask = 16'hF0AC;
defparam \Mux47~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N16
cycloneive_lcell_comb \Mux47~8 (
// Equation(s):
// \Mux47~8_combout  = (cuifregT_3 & ((\Mux47~7_combout  & ((\registerArray[31][16]~q ))) # (!\Mux47~7_combout  & (\registerArray[27][16]~q )))) # (!cuifregT_3 & (((\Mux47~7_combout ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[27][16]~q ),
	.datac(\registerArray[31][16]~q ),
	.datad(\Mux47~7_combout ),
	.cin(gnd),
	.combout(\Mux47~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~8 .lut_mask = 16'hF588;
defparam \Mux47~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N16
cycloneive_lcell_comb \registerArray[29][16]~feeder (
// Equation(s):
// \registerArray[29][16]~feeder_combout  = \Mux52~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux522),
	.cin(gnd),
	.combout(\registerArray[29][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[29][16]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[29][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N17
dffeas \registerArray[29][16] (
	.clk(clk),
	.d(\registerArray[29][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][16] .is_wysiwyg = "true";
defparam \registerArray[29][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y37_N15
dffeas \registerArray[25][16] (
	.clk(clk),
	.d(Mux522),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][16] .is_wysiwyg = "true";
defparam \registerArray[25][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N24
cycloneive_lcell_comb \registerArray[17][16]~feeder (
// Equation(s):
// \registerArray[17][16]~feeder_combout  = \Mux52~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux522),
	.cin(gnd),
	.combout(\registerArray[17][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[17][16]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[17][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N25
dffeas \registerArray[17][16] (
	.clk(clk),
	.d(\registerArray[17][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][16] .is_wysiwyg = "true";
defparam \registerArray[17][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N2
cycloneive_lcell_comb \Mux47~0 (
// Equation(s):
// \Mux47~0_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[21][16]~q )) # (!cuifregT_2 & ((\registerArray[17][16]~q )))))

	.dataa(\registerArray[21][16]~q ),
	.datab(\registerArray[17][16]~q ),
	.datac(cuifregT_3),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux47~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~0 .lut_mask = 16'hFA0C;
defparam \Mux47~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N10
cycloneive_lcell_comb \Mux47~1 (
// Equation(s):
// \Mux47~1_combout  = (cuifregT_3 & ((\Mux47~0_combout  & (\registerArray[29][16]~q )) # (!\Mux47~0_combout  & ((\registerArray[25][16]~q ))))) # (!cuifregT_3 & (((\Mux47~0_combout ))))

	.dataa(\registerArray[29][16]~q ),
	.datab(\registerArray[25][16]~q ),
	.datac(cuifregT_3),
	.datad(\Mux47~0_combout ),
	.cin(gnd),
	.combout(\Mux47~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~1 .lut_mask = 16'hAFC0;
defparam \Mux47~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N17
dffeas \registerArray[20][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][16] .is_wysiwyg = "true";
defparam \registerArray[20][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y33_N5
dffeas \registerArray[28][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][16] .is_wysiwyg = "true";
defparam \registerArray[28][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N4
cycloneive_lcell_comb \Mux47~5 (
// Equation(s):
// \Mux47~5_combout  = (\Mux47~4_combout  & (((\registerArray[28][16]~q ) # (!cuifregT_2)))) # (!\Mux47~4_combout  & (\registerArray[20][16]~q  & ((cuifregT_2))))

	.dataa(\Mux47~4_combout ),
	.datab(\registerArray[20][16]~q ),
	.datac(\registerArray[28][16]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux47~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~5 .lut_mask = 16'hE4AA;
defparam \Mux47~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y33_N11
dffeas \registerArray[30][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][16] .is_wysiwyg = "true";
defparam \registerArray[30][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N3
dffeas \registerArray[26][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][16] .is_wysiwyg = "true";
defparam \registerArray[26][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N13
dffeas \registerArray[18][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][16] .is_wysiwyg = "true";
defparam \registerArray[18][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N12
cycloneive_lcell_comb \Mux47~2 (
// Equation(s):
// \Mux47~2_combout  = (cuifregT_3 & ((\registerArray[26][16]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[18][16]~q  & !cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[26][16]~q ),
	.datac(\registerArray[18][16]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux47~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~2 .lut_mask = 16'hAAD8;
defparam \Mux47~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N10
cycloneive_lcell_comb \Mux47~3 (
// Equation(s):
// \Mux47~3_combout  = (cuifregT_2 & ((\Mux47~2_combout  & ((\registerArray[30][16]~q ))) # (!\Mux47~2_combout  & (\registerArray[22][16]~q )))) # (!cuifregT_2 & (((\Mux47~2_combout ))))

	.dataa(\registerArray[22][16]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[30][16]~q ),
	.datad(\Mux47~2_combout ),
	.cin(gnd),
	.combout(\Mux47~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~3 .lut_mask = 16'hF388;
defparam \Mux47~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N18
cycloneive_lcell_comb \Mux47~6 (
// Equation(s):
// \Mux47~6_combout  = (cuifregT_1 & ((cuifregT_01) # ((\Mux47~3_combout )))) # (!cuifregT_1 & (!cuifregT_01 & (\Mux47~5_combout )))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\Mux47~5_combout ),
	.datad(\Mux47~3_combout ),
	.cin(gnd),
	.combout(\Mux47~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~6 .lut_mask = 16'hBA98;
defparam \Mux47~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N4
cycloneive_lcell_comb \registerArray[14][16]~feeder (
// Equation(s):
// \registerArray[14][16]~feeder_combout  = \Mux52~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux522),
	.cin(gnd),
	.combout(\registerArray[14][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][16]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[14][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y40_N5
dffeas \registerArray[14][16] (
	.clk(clk),
	.d(\registerArray[14][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][16] .is_wysiwyg = "true";
defparam \registerArray[14][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N5
dffeas \registerArray[15][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][16] .is_wysiwyg = "true";
defparam \registerArray[15][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N11
dffeas \registerArray[12][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][16] .is_wysiwyg = "true";
defparam \registerArray[12][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N10
cycloneive_lcell_comb \Mux47~17 (
// Equation(s):
// \Mux47~17_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[13][16]~q )) # (!cuifregT_01 & ((\registerArray[12][16]~q )))))

	.dataa(\registerArray[13][16]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[12][16]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux47~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~17 .lut_mask = 16'hEE30;
defparam \Mux47~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N4
cycloneive_lcell_comb \Mux47~18 (
// Equation(s):
// \Mux47~18_combout  = (cuifregT_1 & ((\Mux47~17_combout  & ((\registerArray[15][16]~q ))) # (!\Mux47~17_combout  & (\registerArray[14][16]~q )))) # (!cuifregT_1 & (((\Mux47~17_combout ))))

	.dataa(\registerArray[14][16]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[15][16]~q ),
	.datad(\Mux47~17_combout ),
	.cin(gnd),
	.combout(\Mux47~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~18 .lut_mask = 16'hF388;
defparam \Mux47~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y37_N15
dffeas \registerArray[2][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][16] .is_wysiwyg = "true";
defparam \registerArray[2][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y40_N21
dffeas \registerArray[1][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][16] .is_wysiwyg = "true";
defparam \registerArray[1][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N20
cycloneive_lcell_comb \Mux47~14 (
// Equation(s):
// \Mux47~14_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][16]~q )) # (!cuifregT_1 & ((\registerArray[1][16]~q )))))

	.dataa(\registerArray[3][16]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[1][16]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux47~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~14 .lut_mask = 16'hB800;
defparam \Mux47~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N14
cycloneive_lcell_comb \Mux47~15 (
// Equation(s):
// \Mux47~15_combout  = (\Mux47~14_combout ) # ((cuifregT_1 & (!cuifregT_01 & \registerArray[2][16]~q )))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\registerArray[2][16]~q ),
	.datad(\Mux47~14_combout ),
	.cin(gnd),
	.combout(\Mux47~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~15 .lut_mask = 16'hFF20;
defparam \Mux47~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N17
dffeas \registerArray[6][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][16] .is_wysiwyg = "true";
defparam \registerArray[6][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N27
dffeas \registerArray[4][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][16] .is_wysiwyg = "true";
defparam \registerArray[4][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N26
cycloneive_lcell_comb \Mux47~12 (
// Equation(s):
// \Mux47~12_combout  = (cuifregT_01 & ((\registerArray[5][16]~q ) # ((cuifregT_1)))) # (!cuifregT_01 & (((\registerArray[4][16]~q  & !cuifregT_1))))

	.dataa(\registerArray[5][16]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[4][16]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux47~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~12 .lut_mask = 16'hCCB8;
defparam \Mux47~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N24
cycloneive_lcell_comb \Mux47~13 (
// Equation(s):
// \Mux47~13_combout  = (cuifregT_1 & ((\Mux47~12_combout  & (\registerArray[7][16]~q )) # (!\Mux47~12_combout  & ((\registerArray[6][16]~q ))))) # (!cuifregT_1 & (((\Mux47~12_combout ))))

	.dataa(\registerArray[7][16]~q ),
	.datab(\registerArray[6][16]~q ),
	.datac(cuifregT_1),
	.datad(\Mux47~12_combout ),
	.cin(gnd),
	.combout(\Mux47~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~13 .lut_mask = 16'hAFC0;
defparam \Mux47~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N8
cycloneive_lcell_comb \Mux47~16 (
// Equation(s):
// \Mux47~16_combout  = (cuifregT_2 & ((cuifregT_3) # ((\Mux47~13_combout )))) # (!cuifregT_2 & (!cuifregT_3 & (\Mux47~15_combout )))

	.dataa(cuifregT_2),
	.datab(cuifregT_3),
	.datac(\Mux47~15_combout ),
	.datad(\Mux47~13_combout ),
	.cin(gnd),
	.combout(\Mux47~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~16 .lut_mask = 16'hBA98;
defparam \Mux47~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N1
dffeas \registerArray[9][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][16] .is_wysiwyg = "true";
defparam \registerArray[9][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N9
dffeas \registerArray[8][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][16] .is_wysiwyg = "true";
defparam \registerArray[8][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N8
cycloneive_lcell_comb \Mux47~10 (
// Equation(s):
// \Mux47~10_combout  = (cuifregT_1 & ((\registerArray[10][16]~q ) # ((cuifregT_01)))) # (!cuifregT_1 & (((\registerArray[8][16]~q  & !cuifregT_01))))

	.dataa(\registerArray[10][16]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[8][16]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux47~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~10 .lut_mask = 16'hCCB8;
defparam \Mux47~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y43_N3
dffeas \registerArray[11][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][16] .is_wysiwyg = "true";
defparam \registerArray[11][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N2
cycloneive_lcell_comb \Mux47~11 (
// Equation(s):
// \Mux47~11_combout  = (\Mux47~10_combout  & (((\registerArray[11][16]~q ) # (!cuifregT_01)))) # (!\Mux47~10_combout  & (\registerArray[9][16]~q  & ((cuifregT_01))))

	.dataa(\registerArray[9][16]~q ),
	.datab(\Mux47~10_combout ),
	.datac(\registerArray[11][16]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux47~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~11 .lut_mask = 16'hE2CC;
defparam \Mux47~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N2
cycloneive_lcell_comb \registerArray[6][15]~feeder (
// Equation(s):
// \registerArray[6][15]~feeder_combout  = \Mux53~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux532),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[6][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[6][15]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[6][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N3
dffeas \registerArray[6][15] (
	.clk(clk),
	.d(\registerArray[6][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][15] .is_wysiwyg = "true";
defparam \registerArray[6][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N31
dffeas \registerArray[7][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][15] .is_wysiwyg = "true";
defparam \registerArray[7][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N1
dffeas \registerArray[4][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][15] .is_wysiwyg = "true";
defparam \registerArray[4][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N0
cycloneive_lcell_comb \Mux48~0 (
// Equation(s):
// \Mux48~0_combout  = (cuifregT_01 & ((\registerArray[5][15]~q ) # ((cuifregT_1)))) # (!cuifregT_01 & (((\registerArray[4][15]~q  & !cuifregT_1))))

	.dataa(\registerArray[5][15]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[4][15]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux48~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~0 .lut_mask = 16'hCCB8;
defparam \Mux48~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N30
cycloneive_lcell_comb \Mux48~1 (
// Equation(s):
// \Mux48~1_combout  = (cuifregT_1 & ((\Mux48~0_combout  & ((\registerArray[7][15]~q ))) # (!\Mux48~0_combout  & (\registerArray[6][15]~q )))) # (!cuifregT_1 & (((\Mux48~0_combout ))))

	.dataa(\registerArray[6][15]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[7][15]~q ),
	.datad(\Mux48~0_combout ),
	.cin(gnd),
	.combout(\Mux48~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~1 .lut_mask = 16'hF388;
defparam \Mux48~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N14
cycloneive_lcell_comb \registerArray[14][15]~feeder (
// Equation(s):
// \registerArray[14][15]~feeder_combout  = \Mux53~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux532),
	.cin(gnd),
	.combout(\registerArray[14][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][15]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[14][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N15
dffeas \registerArray[14][15] (
	.clk(clk),
	.d(\registerArray[14][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][15] .is_wysiwyg = "true";
defparam \registerArray[14][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N25
dffeas \registerArray[15][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][15] .is_wysiwyg = "true";
defparam \registerArray[15][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N3
dffeas \registerArray[12][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][15] .is_wysiwyg = "true";
defparam \registerArray[12][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N2
cycloneive_lcell_comb \Mux48~7 (
// Equation(s):
// \Mux48~7_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[13][15]~q )) # (!cuifregT_01 & ((\registerArray[12][15]~q )))))

	.dataa(\registerArray[13][15]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[12][15]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux48~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~7 .lut_mask = 16'hEE30;
defparam \Mux48~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N24
cycloneive_lcell_comb \Mux48~8 (
// Equation(s):
// \Mux48~8_combout  = (cuifregT_1 & ((\Mux48~7_combout  & ((\registerArray[15][15]~q ))) # (!\Mux48~7_combout  & (\registerArray[14][15]~q )))) # (!cuifregT_1 & (((\Mux48~7_combout ))))

	.dataa(\registerArray[14][15]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[15][15]~q ),
	.datad(\Mux48~7_combout ),
	.cin(gnd),
	.combout(\Mux48~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~8 .lut_mask = 16'hF388;
defparam \Mux48~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y40_N1
dffeas \registerArray[2][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][15] .is_wysiwyg = "true";
defparam \registerArray[2][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y40_N19
dffeas \registerArray[1][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][15] .is_wysiwyg = "true";
defparam \registerArray[1][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N2
cycloneive_lcell_comb \registerArray[3][15]~feeder (
// Equation(s):
// \registerArray[3][15]~feeder_combout  = \Mux53~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux532),
	.cin(gnd),
	.combout(\registerArray[3][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[3][15]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[3][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N3
dffeas \registerArray[3][15] (
	.clk(clk),
	.d(\registerArray[3][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][15] .is_wysiwyg = "true";
defparam \registerArray[3][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N18
cycloneive_lcell_comb \Mux48~4 (
// Equation(s):
// \Mux48~4_combout  = (cuifregT_01 & ((cuifregT_1 & ((\registerArray[3][15]~q ))) # (!cuifregT_1 & (\registerArray[1][15]~q ))))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[1][15]~q ),
	.datad(\registerArray[3][15]~q ),
	.cin(gnd),
	.combout(\Mux48~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~4 .lut_mask = 16'hA820;
defparam \Mux48~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N0
cycloneive_lcell_comb \Mux48~5 (
// Equation(s):
// \Mux48~5_combout  = (\Mux48~4_combout ) # ((!cuifregT_01 & (cuifregT_1 & \registerArray[2][15]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[2][15]~q ),
	.datad(\Mux48~4_combout ),
	.cin(gnd),
	.combout(\Mux48~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~5 .lut_mask = 16'hFF40;
defparam \Mux48~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y31_N27
dffeas \registerArray[11][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][15] .is_wysiwyg = "true";
defparam \registerArray[11][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N13
dffeas \registerArray[8][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][15] .is_wysiwyg = "true";
defparam \registerArray[8][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N12
cycloneive_lcell_comb \Mux48~2 (
// Equation(s):
// \Mux48~2_combout  = (cuifregT_1 & ((\registerArray[10][15]~q ) # ((cuifregT_01)))) # (!cuifregT_1 & (((\registerArray[8][15]~q  & !cuifregT_01))))

	.dataa(\registerArray[10][15]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[8][15]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux48~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~2 .lut_mask = 16'hCCB8;
defparam \Mux48~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N26
cycloneive_lcell_comb \Mux48~3 (
// Equation(s):
// \Mux48~3_combout  = (cuifregT_01 & ((\Mux48~2_combout  & ((\registerArray[11][15]~q ))) # (!\Mux48~2_combout  & (\registerArray[9][15]~q )))) # (!cuifregT_01 & (((\Mux48~2_combout ))))

	.dataa(\registerArray[9][15]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[11][15]~q ),
	.datad(\Mux48~2_combout ),
	.cin(gnd),
	.combout(\Mux48~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~3 .lut_mask = 16'hF388;
defparam \Mux48~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N20
cycloneive_lcell_comb \Mux48~6 (
// Equation(s):
// \Mux48~6_combout  = (cuifregT_3 & ((cuifregT_2) # ((\Mux48~3_combout )))) # (!cuifregT_3 & (!cuifregT_2 & (\Mux48~5_combout )))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\Mux48~5_combout ),
	.datad(\Mux48~3_combout ),
	.cin(gnd),
	.combout(\Mux48~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~6 .lut_mask = 16'hBA98;
defparam \Mux48~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y30_N21
dffeas \registerArray[21][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][15] .is_wysiwyg = "true";
defparam \registerArray[21][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N31
dffeas \registerArray[29][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][15] .is_wysiwyg = "true";
defparam \registerArray[29][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N29
dffeas \registerArray[17][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][15] .is_wysiwyg = "true";
defparam \registerArray[17][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N28
cycloneive_lcell_comb \Mux48~10 (
// Equation(s):
// \Mux48~10_combout  = (cuifregT_3 & ((\registerArray[25][15]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[17][15]~q  & !cuifregT_2))))

	.dataa(\registerArray[25][15]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[17][15]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux48~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~10 .lut_mask = 16'hCCB8;
defparam \Mux48~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N30
cycloneive_lcell_comb \Mux48~11 (
// Equation(s):
// \Mux48~11_combout  = (cuifregT_2 & ((\Mux48~10_combout  & ((\registerArray[29][15]~q ))) # (!\Mux48~10_combout  & (\registerArray[21][15]~q )))) # (!cuifregT_2 & (((\Mux48~10_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[21][15]~q ),
	.datac(\registerArray[29][15]~q ),
	.datad(\Mux48~10_combout ),
	.cin(gnd),
	.combout(\Mux48~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~11 .lut_mask = 16'hF588;
defparam \Mux48~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N0
cycloneive_lcell_comb \registerArray[23][15]~feeder (
// Equation(s):
// \registerArray[23][15]~feeder_combout  = \Mux53~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux532),
	.cin(gnd),
	.combout(\registerArray[23][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[23][15]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[23][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y44_N1
dffeas \registerArray[23][15] (
	.clk(clk),
	.d(\registerArray[23][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][15] .is_wysiwyg = "true";
defparam \registerArray[23][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N3
dffeas \registerArray[31][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][15] .is_wysiwyg = "true";
defparam \registerArray[31][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N30
cycloneive_lcell_comb \registerArray[27][15]~feeder (
// Equation(s):
// \registerArray[27][15]~feeder_combout  = \Mux53~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux532),
	.cin(gnd),
	.combout(\registerArray[27][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[27][15]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[27][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y44_N31
dffeas \registerArray[27][15] (
	.clk(clk),
	.d(\registerArray[27][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][15] .is_wysiwyg = "true";
defparam \registerArray[27][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N12
cycloneive_lcell_comb \Mux48~17 (
// Equation(s):
// \Mux48~17_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & ((\registerArray[27][15]~q ))) # (!cuifregT_3 & (\registerArray[19][15]~q ))))

	.dataa(\registerArray[19][15]~q ),
	.datab(\registerArray[27][15]~q ),
	.datac(cuifregT_2),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux48~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~17 .lut_mask = 16'hFC0A;
defparam \Mux48~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N2
cycloneive_lcell_comb \Mux48~18 (
// Equation(s):
// \Mux48~18_combout  = (cuifregT_2 & ((\Mux48~17_combout  & ((\registerArray[31][15]~q ))) # (!\Mux48~17_combout  & (\registerArray[23][15]~q )))) # (!cuifregT_2 & (((\Mux48~17_combout ))))

	.dataa(\registerArray[23][15]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[31][15]~q ),
	.datad(\Mux48~17_combout ),
	.cin(gnd),
	.combout(\Mux48~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~18 .lut_mask = 16'hF388;
defparam \Mux48~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N28
cycloneive_lcell_comb \registerArray[28][15]~feeder (
// Equation(s):
// \registerArray[28][15]~feeder_combout  = \Mux53~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux532),
	.cin(gnd),
	.combout(\registerArray[28][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[28][15]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[28][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N29
dffeas \registerArray[28][15] (
	.clk(clk),
	.d(\registerArray[28][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][15] .is_wysiwyg = "true";
defparam \registerArray[28][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N4
cycloneive_lcell_comb \registerArray[16][15]~feeder (
// Equation(s):
// \registerArray[16][15]~feeder_combout  = \Mux53~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux532),
	.cin(gnd),
	.combout(\registerArray[16][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[16][15]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[16][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y41_N5
dffeas \registerArray[16][15] (
	.clk(clk),
	.d(\registerArray[16][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][15] .is_wysiwyg = "true";
defparam \registerArray[16][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N10
cycloneive_lcell_comb \Mux48~14 (
// Equation(s):
// \Mux48~14_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[20][15]~q )) # (!cuifregT_2 & ((\registerArray[16][15]~q )))))

	.dataa(\registerArray[20][15]~q ),
	.datab(\registerArray[16][15]~q ),
	.datac(cuifregT_3),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux48~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~14 .lut_mask = 16'hFA0C;
defparam \Mux48~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N26
cycloneive_lcell_comb \Mux48~15 (
// Equation(s):
// \Mux48~15_combout  = (cuifregT_3 & ((\Mux48~14_combout  & ((\registerArray[28][15]~q ))) # (!\Mux48~14_combout  & (\registerArray[24][15]~q )))) # (!cuifregT_3 & (((\Mux48~14_combout ))))

	.dataa(\registerArray[24][15]~q ),
	.datab(\registerArray[28][15]~q ),
	.datac(cuifregT_3),
	.datad(\Mux48~14_combout ),
	.cin(gnd),
	.combout(\Mux48~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~15 .lut_mask = 16'hCFA0;
defparam \Mux48~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N12
cycloneive_lcell_comb \registerArray[26][15]~feeder (
// Equation(s):
// \registerArray[26][15]~feeder_combout  = \Mux53~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux532),
	.cin(gnd),
	.combout(\registerArray[26][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[26][15]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[26][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N13
dffeas \registerArray[26][15] (
	.clk(clk),
	.d(\registerArray[26][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][15] .is_wysiwyg = "true";
defparam \registerArray[26][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N23
dffeas \registerArray[30][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][15] .is_wysiwyg = "true";
defparam \registerArray[30][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y37_N11
dffeas \registerArray[18][15] (
	.clk(clk),
	.d(Mux532),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][15] .is_wysiwyg = "true";
defparam \registerArray[18][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y40_N21
dffeas \registerArray[22][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][15] .is_wysiwyg = "true";
defparam \registerArray[22][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N20
cycloneive_lcell_comb \Mux48~12 (
// Equation(s):
// \Mux48~12_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & ((\registerArray[22][15]~q ))) # (!cuifregT_2 & (\registerArray[18][15]~q ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[18][15]~q ),
	.datac(\registerArray[22][15]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux48~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~12 .lut_mask = 16'hFA44;
defparam \Mux48~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N22
cycloneive_lcell_comb \Mux48~13 (
// Equation(s):
// \Mux48~13_combout  = (cuifregT_3 & ((\Mux48~12_combout  & ((\registerArray[30][15]~q ))) # (!\Mux48~12_combout  & (\registerArray[26][15]~q )))) # (!cuifregT_3 & (((\Mux48~12_combout ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[26][15]~q ),
	.datac(\registerArray[30][15]~q ),
	.datad(\Mux48~12_combout ),
	.cin(gnd),
	.combout(\Mux48~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~13 .lut_mask = 16'hF588;
defparam \Mux48~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y41_N16
cycloneive_lcell_comb \Mux48~16 (
// Equation(s):
// \Mux48~16_combout  = (cuifregT_1 & ((cuifregT_01) # ((\Mux48~13_combout )))) # (!cuifregT_1 & (!cuifregT_01 & (\Mux48~15_combout )))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\Mux48~15_combout ),
	.datad(\Mux48~13_combout ),
	.cin(gnd),
	.combout(\Mux48~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~16 .lut_mask = 16'hBA98;
defparam \Mux48~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N23
dffeas \registerArray[12][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][14] .is_wysiwyg = "true";
defparam \registerArray[12][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N22
cycloneive_lcell_comb \Mux49~7 (
// Equation(s):
// \Mux49~7_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[13][14]~q )) # (!cuifregT_01 & ((\registerArray[12][14]~q )))))

	.dataa(\registerArray[13][14]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[12][14]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux49~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~7 .lut_mask = 16'hEE30;
defparam \Mux49~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N1
dffeas \registerArray[15][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][14] .is_wysiwyg = "true";
defparam \registerArray[15][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N24
cycloneive_lcell_comb \registerArray[14][14]~feeder (
// Equation(s):
// \registerArray[14][14]~feeder_combout  = \Mux54~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux542),
	.cin(gnd),
	.combout(\registerArray[14][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][14]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[14][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y32_N25
dffeas \registerArray[14][14] (
	.clk(clk),
	.d(\registerArray[14][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][14] .is_wysiwyg = "true";
defparam \registerArray[14][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N0
cycloneive_lcell_comb \Mux49~8 (
// Equation(s):
// \Mux49~8_combout  = (\Mux49~7_combout  & (((\registerArray[15][14]~q )) # (!cuifregT_1))) # (!\Mux49~7_combout  & (cuifregT_1 & ((\registerArray[14][14]~q ))))

	.dataa(\Mux49~7_combout ),
	.datab(cuifregT_1),
	.datac(\registerArray[15][14]~q ),
	.datad(\registerArray[14][14]~q ),
	.cin(gnd),
	.combout(\Mux49~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~8 .lut_mask = 16'hE6A2;
defparam \Mux49~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N29
dffeas \registerArray[9][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][14] .is_wysiwyg = "true";
defparam \registerArray[9][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N31
dffeas \registerArray[11][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][14] .is_wysiwyg = "true";
defparam \registerArray[11][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N17
dffeas \registerArray[8][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][14] .is_wysiwyg = "true";
defparam \registerArray[8][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N16
cycloneive_lcell_comb \Mux49~0 (
// Equation(s):
// \Mux49~0_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & (\registerArray[10][14]~q )) # (!cuifregT_1 & ((\registerArray[8][14]~q )))))

	.dataa(\registerArray[10][14]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[8][14]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux49~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~0 .lut_mask = 16'hEE30;
defparam \Mux49~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N30
cycloneive_lcell_comb \Mux49~1 (
// Equation(s):
// \Mux49~1_combout  = (cuifregT_01 & ((\Mux49~0_combout  & ((\registerArray[11][14]~q ))) # (!\Mux49~0_combout  & (\registerArray[9][14]~q )))) # (!cuifregT_01 & (((\Mux49~0_combout ))))

	.dataa(\registerArray[9][14]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[11][14]~q ),
	.datad(\Mux49~0_combout ),
	.cin(gnd),
	.combout(\Mux49~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~1 .lut_mask = 16'hF388;
defparam \Mux49~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y31_N23
dffeas \registerArray[7][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][14] .is_wysiwyg = "true";
defparam \registerArray[7][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N25
dffeas \registerArray[4][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][14] .is_wysiwyg = "true";
defparam \registerArray[4][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N24
cycloneive_lcell_comb \Mux49~2 (
// Equation(s):
// \Mux49~2_combout  = (cuifregT_01 & ((\registerArray[5][14]~q ) # ((cuifregT_1)))) # (!cuifregT_01 & (((\registerArray[4][14]~q  & !cuifregT_1))))

	.dataa(\registerArray[5][14]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[4][14]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux49~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~2 .lut_mask = 16'hCCB8;
defparam \Mux49~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N22
cycloneive_lcell_comb \Mux49~3 (
// Equation(s):
// \Mux49~3_combout  = (cuifregT_1 & ((\Mux49~2_combout  & ((\registerArray[7][14]~q ))) # (!\Mux49~2_combout  & (\registerArray[6][14]~q )))) # (!cuifregT_1 & (((\Mux49~2_combout ))))

	.dataa(\registerArray[6][14]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[7][14]~q ),
	.datad(\Mux49~2_combout ),
	.cin(gnd),
	.combout(\Mux49~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~3 .lut_mask = 16'hF388;
defparam \Mux49~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y43_N27
dffeas \registerArray[2][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][14] .is_wysiwyg = "true";
defparam \registerArray[2][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y37_N5
dffeas \registerArray[3][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][14] .is_wysiwyg = "true";
defparam \registerArray[3][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y43_N25
dffeas \registerArray[1][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][14] .is_wysiwyg = "true";
defparam \registerArray[1][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N24
cycloneive_lcell_comb \Mux49~4 (
// Equation(s):
// \Mux49~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][14]~q )) # (!cuifregT_1 & ((\registerArray[1][14]~q )))))

	.dataa(cuifregT_0),
	.datab(\registerArray[3][14]~q ),
	.datac(\registerArray[1][14]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux49~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~4 .lut_mask = 16'h88A0;
defparam \Mux49~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N26
cycloneive_lcell_comb \Mux49~5 (
// Equation(s):
// \Mux49~5_combout  = (\Mux49~4_combout ) # ((!cuifregT_01 & (cuifregT_1 & \registerArray[2][14]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[2][14]~q ),
	.datad(\Mux49~4_combout ),
	.cin(gnd),
	.combout(\Mux49~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~5 .lut_mask = 16'hFF40;
defparam \Mux49~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N20
cycloneive_lcell_comb \Mux49~6 (
// Equation(s):
// \Mux49~6_combout  = (cuifregT_3 & (cuifregT_2)) # (!cuifregT_3 & ((cuifregT_2 & (\Mux49~3_combout )) # (!cuifregT_2 & ((\Mux49~5_combout )))))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\Mux49~3_combout ),
	.datad(\Mux49~5_combout ),
	.cin(gnd),
	.combout(\Mux49~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~6 .lut_mask = 16'hD9C8;
defparam \Mux49~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N18
cycloneive_lcell_comb \registerArray[27][14]~feeder (
// Equation(s):
// \registerArray[27][14]~feeder_combout  = \Mux54~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux542),
	.cin(gnd),
	.combout(\registerArray[27][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[27][14]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[27][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y37_N19
dffeas \registerArray[27][14] (
	.clk(clk),
	.d(\registerArray[27][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][14] .is_wysiwyg = "true";
defparam \registerArray[27][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N7
dffeas \registerArray[31][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][14] .is_wysiwyg = "true";
defparam \registerArray[31][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N29
dffeas \registerArray[19][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][14] .is_wysiwyg = "true";
defparam \registerArray[19][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N28
cycloneive_lcell_comb \Mux49~17 (
// Equation(s):
// \Mux49~17_combout  = (cuifregT_2 & ((\registerArray[23][14]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[19][14]~q  & !cuifregT_3))))

	.dataa(\registerArray[23][14]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[19][14]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux49~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~17 .lut_mask = 16'hCCB8;
defparam \Mux49~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N6
cycloneive_lcell_comb \Mux49~18 (
// Equation(s):
// \Mux49~18_combout  = (cuifregT_3 & ((\Mux49~17_combout  & ((\registerArray[31][14]~q ))) # (!\Mux49~17_combout  & (\registerArray[27][14]~q )))) # (!cuifregT_3 & (((\Mux49~17_combout ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[27][14]~q ),
	.datac(\registerArray[31][14]~q ),
	.datad(\Mux49~17_combout ),
	.cin(gnd),
	.combout(\Mux49~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~18 .lut_mask = 16'hF588;
defparam \Mux49~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N29
dffeas \registerArray[20][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][14] .is_wysiwyg = "true";
defparam \registerArray[20][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y37_N27
dffeas \registerArray[28][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][14] .is_wysiwyg = "true";
defparam \registerArray[28][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N2
cycloneive_lcell_comb \registerArray[16][14]~feeder (
// Equation(s):
// \registerArray[16][14]~feeder_combout  = \Mux54~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux542),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[16][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[16][14]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[16][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y37_N3
dffeas \registerArray[16][14] (
	.clk(clk),
	.d(\registerArray[16][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][14] .is_wysiwyg = "true";
defparam \registerArray[16][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N31
dffeas \registerArray[24][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][14] .is_wysiwyg = "true";
defparam \registerArray[24][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N16
cycloneive_lcell_comb \Mux49~14 (
// Equation(s):
// \Mux49~14_combout  = (cuifregT_3 & (((\registerArray[24][14]~q ) # (cuifregT_2)))) # (!cuifregT_3 & (\registerArray[16][14]~q  & ((!cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[16][14]~q ),
	.datac(\registerArray[24][14]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux49~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~14 .lut_mask = 16'hAAE4;
defparam \Mux49~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N26
cycloneive_lcell_comb \Mux49~15 (
// Equation(s):
// \Mux49~15_combout  = (cuifregT_2 & ((\Mux49~14_combout  & ((\registerArray[28][14]~q ))) # (!\Mux49~14_combout  & (\registerArray[20][14]~q )))) # (!cuifregT_2 & (((\Mux49~14_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[20][14]~q ),
	.datac(\registerArray[28][14]~q ),
	.datad(\Mux49~14_combout ),
	.cin(gnd),
	.combout(\Mux49~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~15 .lut_mask = 16'hF588;
defparam \Mux49~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y33_N7
dffeas \registerArray[30][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][14] .is_wysiwyg = "true";
defparam \registerArray[30][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N29
dffeas \registerArray[18][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][14] .is_wysiwyg = "true";
defparam \registerArray[18][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N23
dffeas \registerArray[26][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][14] .is_wysiwyg = "true";
defparam \registerArray[26][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N28
cycloneive_lcell_comb \Mux49~12 (
// Equation(s):
// \Mux49~12_combout  = (cuifregT_3 & ((cuifregT_2) # ((\registerArray[26][14]~q )))) # (!cuifregT_3 & (!cuifregT_2 & (\registerArray[18][14]~q )))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\registerArray[18][14]~q ),
	.datad(\registerArray[26][14]~q ),
	.cin(gnd),
	.combout(\Mux49~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~12 .lut_mask = 16'hBA98;
defparam \Mux49~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N6
cycloneive_lcell_comb \Mux49~13 (
// Equation(s):
// \Mux49~13_combout  = (cuifregT_2 & ((\Mux49~12_combout  & ((\registerArray[30][14]~q ))) # (!\Mux49~12_combout  & (\registerArray[22][14]~q )))) # (!cuifregT_2 & (((\Mux49~12_combout ))))

	.dataa(\registerArray[22][14]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[30][14]~q ),
	.datad(\Mux49~12_combout ),
	.cin(gnd),
	.combout(\Mux49~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~13 .lut_mask = 16'hF388;
defparam \Mux49~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y37_N4
cycloneive_lcell_comb \Mux49~16 (
// Equation(s):
// \Mux49~16_combout  = (cuifregT_01 & (cuifregT_1)) # (!cuifregT_01 & ((cuifregT_1 & ((\Mux49~13_combout ))) # (!cuifregT_1 & (\Mux49~15_combout ))))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\Mux49~15_combout ),
	.datad(\Mux49~13_combout ),
	.cin(gnd),
	.combout(\Mux49~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~16 .lut_mask = 16'hDC98;
defparam \Mux49~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y41_N13
dffeas \registerArray[25][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][14] .is_wysiwyg = "true";
defparam \registerArray[25][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N11
dffeas \registerArray[29][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][14] .is_wysiwyg = "true";
defparam \registerArray[29][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N1
dffeas \registerArray[17][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][14] .is_wysiwyg = "true";
defparam \registerArray[17][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N0
cycloneive_lcell_comb \Mux49~10 (
// Equation(s):
// \Mux49~10_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[21][14]~q )) # (!cuifregT_2 & ((\registerArray[17][14]~q )))))

	.dataa(\registerArray[21][14]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[17][14]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux49~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~10 .lut_mask = 16'hEE30;
defparam \Mux49~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N10
cycloneive_lcell_comb \Mux49~11 (
// Equation(s):
// \Mux49~11_combout  = (cuifregT_3 & ((\Mux49~10_combout  & ((\registerArray[29][14]~q ))) # (!\Mux49~10_combout  & (\registerArray[25][14]~q )))) # (!cuifregT_3 & (((\Mux49~10_combout ))))

	.dataa(\registerArray[25][14]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[29][14]~q ),
	.datad(\Mux49~10_combout ),
	.cin(gnd),
	.combout(\Mux49~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~11 .lut_mask = 16'hF388;
defparam \Mux49~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N18
cycloneive_lcell_comb \registerArray[14][13]~feeder (
// Equation(s):
// \registerArray[14][13]~feeder_combout  = \Mux55~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux552),
	.cin(gnd),
	.combout(\registerArray[14][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][13]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[14][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N19
dffeas \registerArray[14][13] (
	.clk(clk),
	.d(\registerArray[14][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][13] .is_wysiwyg = "true";
defparam \registerArray[14][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N4
cycloneive_lcell_comb \registerArray[15][13]~feeder (
// Equation(s):
// \registerArray[15][13]~feeder_combout  = \Mux55~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux552),
	.cin(gnd),
	.combout(\registerArray[15][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[15][13]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[15][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y32_N5
dffeas \registerArray[15][13] (
	.clk(clk),
	.d(\registerArray[15][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][13] .is_wysiwyg = "true";
defparam \registerArray[15][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N0
cycloneive_lcell_comb \registerArray[12][13]~feeder (
// Equation(s):
// \registerArray[12][13]~feeder_combout  = \Mux55~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux552),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[12][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[12][13]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[12][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N1
dffeas \registerArray[12][13] (
	.clk(clk),
	.d(\registerArray[12][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][13] .is_wysiwyg = "true";
defparam \registerArray[12][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N11
dffeas \registerArray[13][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][13] .is_wysiwyg = "true";
defparam \registerArray[13][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N18
cycloneive_lcell_comb \Mux50~7 (
// Equation(s):
// \Mux50~7_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & ((\registerArray[13][13]~q ))) # (!cuifregT_01 & (\registerArray[12][13]~q ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[12][13]~q ),
	.datac(cuifregT_0),
	.datad(\registerArray[13][13]~q ),
	.cin(gnd),
	.combout(\Mux50~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~7 .lut_mask = 16'hF4A4;
defparam \Mux50~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N14
cycloneive_lcell_comb \Mux50~8 (
// Equation(s):
// \Mux50~8_combout  = (cuifregT_1 & ((\Mux50~7_combout  & ((\registerArray[15][13]~q ))) # (!\Mux50~7_combout  & (\registerArray[14][13]~q )))) # (!cuifregT_1 & (((\Mux50~7_combout ))))

	.dataa(\registerArray[14][13]~q ),
	.datab(\registerArray[15][13]~q ),
	.datac(cuifregT_1),
	.datad(\Mux50~7_combout ),
	.cin(gnd),
	.combout(\Mux50~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~8 .lut_mask = 16'hCFA0;
defparam \Mux50~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N7
dffeas \registerArray[6][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][13] .is_wysiwyg = "true";
defparam \registerArray[6][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N5
dffeas \registerArray[4][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][13] .is_wysiwyg = "true";
defparam \registerArray[4][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N4
cycloneive_lcell_comb \Mux50~0 (
// Equation(s):
// \Mux50~0_combout  = (cuifregT_01 & ((\registerArray[5][13]~q ) # ((cuifregT_1)))) # (!cuifregT_01 & (((\registerArray[4][13]~q  & !cuifregT_1))))

	.dataa(\registerArray[5][13]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[4][13]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux50~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~0 .lut_mask = 16'hCCB8;
defparam \Mux50~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y31_N3
dffeas \registerArray[7][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][13] .is_wysiwyg = "true";
defparam \registerArray[7][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N2
cycloneive_lcell_comb \Mux50~1 (
// Equation(s):
// \Mux50~1_combout  = (\Mux50~0_combout  & (((\registerArray[7][13]~q ) # (!cuifregT_1)))) # (!\Mux50~0_combout  & (\registerArray[6][13]~q  & ((cuifregT_1))))

	.dataa(\registerArray[6][13]~q ),
	.datab(\Mux50~0_combout ),
	.datac(\registerArray[7][13]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux50~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~1 .lut_mask = 16'hE2CC;
defparam \Mux50~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y43_N3
dffeas \registerArray[2][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][13] .is_wysiwyg = "true";
defparam \registerArray[2][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N28
cycloneive_lcell_comb \registerArray[3][13]~feeder (
// Equation(s):
// \registerArray[3][13]~feeder_combout  = \Mux55~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux552),
	.cin(gnd),
	.combout(\registerArray[3][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[3][13]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[3][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y43_N29
dffeas \registerArray[3][13] (
	.clk(clk),
	.d(\registerArray[3][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][13] .is_wysiwyg = "true";
defparam \registerArray[3][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y43_N21
dffeas \registerArray[1][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][13] .is_wysiwyg = "true";
defparam \registerArray[1][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N20
cycloneive_lcell_comb \Mux50~4 (
// Equation(s):
// \Mux50~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][13]~q )) # (!cuifregT_1 & ((\registerArray[1][13]~q )))))

	.dataa(cuifregT_0),
	.datab(\registerArray[3][13]~q ),
	.datac(\registerArray[1][13]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux50~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~4 .lut_mask = 16'h88A0;
defparam \Mux50~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N2
cycloneive_lcell_comb \Mux50~5 (
// Equation(s):
// \Mux50~5_combout  = (\Mux50~4_combout ) # ((!cuifregT_01 & (cuifregT_1 & \registerArray[2][13]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[2][13]~q ),
	.datad(\Mux50~4_combout ),
	.cin(gnd),
	.combout(\Mux50~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~5 .lut_mask = 16'hFF40;
defparam \Mux50~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y31_N9
dffeas \registerArray[8][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][13] .is_wysiwyg = "true";
defparam \registerArray[8][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N8
cycloneive_lcell_comb \Mux50~2 (
// Equation(s):
// \Mux50~2_combout  = (cuifregT_1 & ((\registerArray[10][13]~q ) # ((cuifregT_01)))) # (!cuifregT_1 & (((\registerArray[8][13]~q  & !cuifregT_01))))

	.dataa(\registerArray[10][13]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[8][13]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux50~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~2 .lut_mask = 16'hCCB8;
defparam \Mux50~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y31_N19
dffeas \registerArray[11][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][13] .is_wysiwyg = "true";
defparam \registerArray[11][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N18
cycloneive_lcell_comb \Mux50~3 (
// Equation(s):
// \Mux50~3_combout  = (\Mux50~2_combout  & (((\registerArray[11][13]~q ) # (!cuifregT_01)))) # (!\Mux50~2_combout  & (\registerArray[9][13]~q  & ((cuifregT_01))))

	.dataa(\registerArray[9][13]~q ),
	.datab(\Mux50~2_combout ),
	.datac(\registerArray[11][13]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux50~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~3 .lut_mask = 16'hE2CC;
defparam \Mux50~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N28
cycloneive_lcell_comb \Mux50~6 (
// Equation(s):
// \Mux50~6_combout  = (cuifregT_3 & ((cuifregT_2) # ((\Mux50~3_combout )))) # (!cuifregT_3 & (!cuifregT_2 & (\Mux50~5_combout )))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\Mux50~5_combout ),
	.datad(\Mux50~3_combout ),
	.cin(gnd),
	.combout(\Mux50~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~6 .lut_mask = 16'hBA98;
defparam \Mux50~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N31
dffeas \registerArray[27][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][13] .is_wysiwyg = "true";
defparam \registerArray[27][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N27
dffeas \registerArray[19][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][13] .is_wysiwyg = "true";
defparam \registerArray[19][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N26
cycloneive_lcell_comb \Mux50~17 (
// Equation(s):
// \Mux50~17_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[27][13]~q )) # (!cuifregT_3 & ((\registerArray[19][13]~q )))))

	.dataa(cuifregT_2),
	.datab(\registerArray[27][13]~q ),
	.datac(\registerArray[19][13]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux50~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~17 .lut_mask = 16'hEE50;
defparam \Mux50~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N29
dffeas \registerArray[23][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][13] .is_wysiwyg = "true";
defparam \registerArray[23][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N21
dffeas \registerArray[31][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][13] .is_wysiwyg = "true";
defparam \registerArray[31][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N20
cycloneive_lcell_comb \Mux50~18 (
// Equation(s):
// \Mux50~18_combout  = (\Mux50~17_combout  & (((\registerArray[31][13]~q ) # (!cuifregT_2)))) # (!\Mux50~17_combout  & (\registerArray[23][13]~q  & ((cuifregT_2))))

	.dataa(\Mux50~17_combout ),
	.datab(\registerArray[23][13]~q ),
	.datac(\registerArray[31][13]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux50~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~18 .lut_mask = 16'hE4AA;
defparam \Mux50~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y33_N5
dffeas \registerArray[18][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][13] .is_wysiwyg = "true";
defparam \registerArray[18][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N7
dffeas \registerArray[22][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][13] .is_wysiwyg = "true";
defparam \registerArray[22][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N4
cycloneive_lcell_comb \Mux50~12 (
// Equation(s):
// \Mux50~12_combout  = (cuifregT_3 & (cuifregT_2)) # (!cuifregT_3 & ((cuifregT_2 & ((\registerArray[22][13]~q ))) # (!cuifregT_2 & (\registerArray[18][13]~q ))))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\registerArray[18][13]~q ),
	.datad(\registerArray[22][13]~q ),
	.cin(gnd),
	.combout(\Mux50~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~12 .lut_mask = 16'hDC98;
defparam \Mux50~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y33_N31
dffeas \registerArray[30][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][13] .is_wysiwyg = "true";
defparam \registerArray[30][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N25
dffeas \registerArray[26][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][13] .is_wysiwyg = "true";
defparam \registerArray[26][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N30
cycloneive_lcell_comb \Mux50~13 (
// Equation(s):
// \Mux50~13_combout  = (cuifregT_3 & ((\Mux50~12_combout  & (\registerArray[30][13]~q )) # (!\Mux50~12_combout  & ((\registerArray[26][13]~q ))))) # (!cuifregT_3 & (\Mux50~12_combout ))

	.dataa(cuifregT_3),
	.datab(\Mux50~12_combout ),
	.datac(\registerArray[30][13]~q ),
	.datad(\registerArray[26][13]~q ),
	.cin(gnd),
	.combout(\Mux50~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~13 .lut_mask = 16'hE6C4;
defparam \Mux50~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N9
dffeas \registerArray[28][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][13] .is_wysiwyg = "true";
defparam \registerArray[28][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N27
dffeas \registerArray[16][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][13] .is_wysiwyg = "true";
defparam \registerArray[16][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N26
cycloneive_lcell_comb \Mux50~14 (
// Equation(s):
// \Mux50~14_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[20][13]~q )) # (!cuifregT_2 & ((\registerArray[16][13]~q )))))

	.dataa(\registerArray[20][13]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[16][13]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux50~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~14 .lut_mask = 16'hEE30;
defparam \Mux50~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N8
cycloneive_lcell_comb \Mux50~15 (
// Equation(s):
// \Mux50~15_combout  = (cuifregT_3 & ((\Mux50~14_combout  & ((\registerArray[28][13]~q ))) # (!\Mux50~14_combout  & (\registerArray[24][13]~q )))) # (!cuifregT_3 & (((\Mux50~14_combout ))))

	.dataa(\registerArray[24][13]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[28][13]~q ),
	.datad(\Mux50~14_combout ),
	.cin(gnd),
	.combout(\Mux50~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~15 .lut_mask = 16'hF388;
defparam \Mux50~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N30
cycloneive_lcell_comb \Mux50~16 (
// Equation(s):
// \Mux50~16_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & (\Mux50~13_combout )) # (!cuifregT_1 & ((\Mux50~15_combout )))))

	.dataa(cuifregT_0),
	.datab(\Mux50~13_combout ),
	.datac(\Mux50~15_combout ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux50~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~16 .lut_mask = 16'hEE50;
defparam \Mux50~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N13
dffeas \registerArray[21][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][13] .is_wysiwyg = "true";
defparam \registerArray[21][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N24
cycloneive_lcell_comb \registerArray[29][13]~feeder (
// Equation(s):
// \registerArray[29][13]~feeder_combout  = \Mux55~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux552),
	.cin(gnd),
	.combout(\registerArray[29][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[29][13]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[29][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N25
dffeas \registerArray[29][13] (
	.clk(clk),
	.d(\registerArray[29][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][13] .is_wysiwyg = "true";
defparam \registerArray[29][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N21
dffeas \registerArray[25][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][13] .is_wysiwyg = "true";
defparam \registerArray[25][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N10
cycloneive_lcell_comb \registerArray[17][13]~feeder (
// Equation(s):
// \registerArray[17][13]~feeder_combout  = \Mux55~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux552),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[17][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[17][13]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[17][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N11
dffeas \registerArray[17][13] (
	.clk(clk),
	.d(\registerArray[17][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][13] .is_wysiwyg = "true";
defparam \registerArray[17][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N22
cycloneive_lcell_comb \Mux50~10 (
// Equation(s):
// \Mux50~10_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[25][13]~q )) # (!cuifregT_3 & ((\registerArray[17][13]~q )))))

	.dataa(cuifregT_2),
	.datab(\registerArray[25][13]~q ),
	.datac(\registerArray[17][13]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux50~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~10 .lut_mask = 16'hEE50;
defparam \Mux50~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N0
cycloneive_lcell_comb \Mux50~11 (
// Equation(s):
// \Mux50~11_combout  = (\Mux50~10_combout  & (((\registerArray[29][13]~q ) # (!cuifregT_2)))) # (!\Mux50~10_combout  & (\registerArray[21][13]~q  & ((cuifregT_2))))

	.dataa(\registerArray[21][13]~q ),
	.datab(\registerArray[29][13]~q ),
	.datac(\Mux50~10_combout ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux50~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~11 .lut_mask = 16'hCAF0;
defparam \Mux50~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N12
cycloneive_lcell_comb \registerArray[14][12]~feeder (
// Equation(s):
// \registerArray[14][12]~feeder_combout  = \Mux56~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux562),
	.cin(gnd),
	.combout(\registerArray[14][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][12]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[14][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y36_N13
dffeas \registerArray[14][12] (
	.clk(clk),
	.d(\registerArray[14][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][12] .is_wysiwyg = "true";
defparam \registerArray[14][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N29
dffeas \registerArray[15][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][12] .is_wysiwyg = "true";
defparam \registerArray[15][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N19
dffeas \registerArray[12][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][12] .is_wysiwyg = "true";
defparam \registerArray[12][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N18
cycloneive_lcell_comb \Mux51~7 (
// Equation(s):
// \Mux51~7_combout  = (cuifregT_01 & ((\registerArray[13][12]~q ) # ((cuifregT_1)))) # (!cuifregT_01 & (((\registerArray[12][12]~q  & !cuifregT_1))))

	.dataa(\registerArray[13][12]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[12][12]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux51~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~7 .lut_mask = 16'hCCB8;
defparam \Mux51~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N28
cycloneive_lcell_comb \Mux51~8 (
// Equation(s):
// \Mux51~8_combout  = (cuifregT_1 & ((\Mux51~7_combout  & ((\registerArray[15][12]~q ))) # (!\Mux51~7_combout  & (\registerArray[14][12]~q )))) # (!cuifregT_1 & (((\Mux51~7_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[14][12]~q ),
	.datac(\registerArray[15][12]~q ),
	.datad(\Mux51~7_combout ),
	.cin(gnd),
	.combout(\Mux51~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~8 .lut_mask = 16'hF588;
defparam \Mux51~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N0
cycloneive_lcell_comb \registerArray[9][12]~feeder (
// Equation(s):
// \registerArray[9][12]~feeder_combout  = \Mux56~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux562),
	.cin(gnd),
	.combout(\registerArray[9][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[9][12]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[9][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y39_N1
dffeas \registerArray[9][12] (
	.clk(clk),
	.d(\registerArray[9][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][12] .is_wysiwyg = "true";
defparam \registerArray[9][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N31
dffeas \registerArray[11][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][12] .is_wysiwyg = "true";
defparam \registerArray[11][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N2
cycloneive_lcell_comb \registerArray[8][12]~feeder (
// Equation(s):
// \registerArray[8][12]~feeder_combout  = \Mux56~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux562),
	.cin(gnd),
	.combout(\registerArray[8][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[8][12]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[8][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y39_N3
dffeas \registerArray[8][12] (
	.clk(clk),
	.d(\registerArray[8][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][12] .is_wysiwyg = "true";
defparam \registerArray[8][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N25
dffeas \registerArray[10][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][12] .is_wysiwyg = "true";
defparam \registerArray[10][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N24
cycloneive_lcell_comb \Mux51~0 (
// Equation(s):
// \Mux51~0_combout  = (cuifregT_1 & (((\registerArray[10][12]~q ) # (cuifregT_01)))) # (!cuifregT_1 & (\registerArray[8][12]~q  & ((!cuifregT_01))))

	.dataa(cuifregT_1),
	.datab(\registerArray[8][12]~q ),
	.datac(\registerArray[10][12]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux51~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~0 .lut_mask = 16'hAAE4;
defparam \Mux51~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N30
cycloneive_lcell_comb \Mux51~1 (
// Equation(s):
// \Mux51~1_combout  = (cuifregT_01 & ((\Mux51~0_combout  & ((\registerArray[11][12]~q ))) # (!\Mux51~0_combout  & (\registerArray[9][12]~q )))) # (!cuifregT_01 & (((\Mux51~0_combout ))))

	.dataa(cuifregT_0),
	.datab(\registerArray[9][12]~q ),
	.datac(\registerArray[11][12]~q ),
	.datad(\Mux51~0_combout ),
	.cin(gnd),
	.combout(\Mux51~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~1 .lut_mask = 16'hF588;
defparam \Mux51~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N8
cycloneive_lcell_comb \registerArray[7][12]~feeder (
// Equation(s):
// \registerArray[7][12]~feeder_combout  = \Mux56~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux562),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[7][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[7][12]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[7][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N9
dffeas \registerArray[7][12] (
	.clk(clk),
	.d(\registerArray[7][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][12] .is_wysiwyg = "true";
defparam \registerArray[7][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y42_N9
dffeas \registerArray[6][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][12] .is_wysiwyg = "true";
defparam \registerArray[6][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N21
dffeas \registerArray[5][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][12] .is_wysiwyg = "true";
defparam \registerArray[5][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N31
dffeas \registerArray[4][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][12] .is_wysiwyg = "true";
defparam \registerArray[4][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N30
cycloneive_lcell_comb \Mux51~2 (
// Equation(s):
// \Mux51~2_combout  = (cuifregT_01 & ((\registerArray[5][12]~q ) # ((cuifregT_1)))) # (!cuifregT_01 & (((\registerArray[4][12]~q  & !cuifregT_1))))

	.dataa(cuifregT_0),
	.datab(\registerArray[5][12]~q ),
	.datac(\registerArray[4][12]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux51~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~2 .lut_mask = 16'hAAD8;
defparam \Mux51~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N26
cycloneive_lcell_comb \Mux51~3 (
// Equation(s):
// \Mux51~3_combout  = (cuifregT_1 & ((\Mux51~2_combout  & (\registerArray[7][12]~q )) # (!\Mux51~2_combout  & ((\registerArray[6][12]~q ))))) # (!cuifregT_1 & (((\Mux51~2_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[7][12]~q ),
	.datac(\registerArray[6][12]~q ),
	.datad(\Mux51~2_combout ),
	.cin(gnd),
	.combout(\Mux51~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~3 .lut_mask = 16'hDDA0;
defparam \Mux51~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N24
cycloneive_lcell_comb \registerArray[2][12]~feeder (
// Equation(s):
// \registerArray[2][12]~feeder_combout  = \Mux56~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux562),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[2][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[2][12]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[2][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y34_N25
dffeas \registerArray[2][12] (
	.clk(clk),
	.d(\registerArray[2][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][12] .is_wysiwyg = "true";
defparam \registerArray[2][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y42_N13
dffeas \registerArray[3][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][12] .is_wysiwyg = "true";
defparam \registerArray[3][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y41_N24
cycloneive_lcell_comb \Mux51~4 (
// Equation(s):
// \Mux51~4_combout  = (cuifregT_01 & ((cuifregT_1 & ((\registerArray[3][12]~q ))) # (!cuifregT_1 & (\registerArray[1][12]~q ))))

	.dataa(\registerArray[1][12]~q ),
	.datab(\registerArray[3][12]~q ),
	.datac(cuifregT_1),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux51~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~4 .lut_mask = 16'hCA00;
defparam \Mux51~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N18
cycloneive_lcell_comb \Mux51~5 (
// Equation(s):
// \Mux51~5_combout  = (\Mux51~4_combout ) # ((cuifregT_1 & (!cuifregT_01 & \registerArray[2][12]~q )))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\registerArray[2][12]~q ),
	.datad(\Mux51~4_combout ),
	.cin(gnd),
	.combout(\Mux51~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~5 .lut_mask = 16'hFF20;
defparam \Mux51~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N16
cycloneive_lcell_comb \Mux51~6 (
// Equation(s):
// \Mux51~6_combout  = (cuifregT_3 & (cuifregT_2)) # (!cuifregT_3 & ((cuifregT_2 & (\Mux51~3_combout )) # (!cuifregT_2 & ((\Mux51~5_combout )))))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\Mux51~3_combout ),
	.datad(\Mux51~5_combout ),
	.cin(gnd),
	.combout(\Mux51~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~6 .lut_mask = 16'hD9C8;
defparam \Mux51~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N26
cycloneive_lcell_comb \registerArray[29][12]~feeder (
// Equation(s):
// \registerArray[29][12]~feeder_combout  = \Mux56~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux562),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[29][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[29][12]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[29][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N27
dffeas \registerArray[29][12] (
	.clk(clk),
	.d(\registerArray[29][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][12] .is_wysiwyg = "true";
defparam \registerArray[29][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N13
dffeas \registerArray[25][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][12] .is_wysiwyg = "true";
defparam \registerArray[25][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N7
dffeas \registerArray[17][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][12] .is_wysiwyg = "true";
defparam \registerArray[17][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N6
cycloneive_lcell_comb \Mux51~10 (
// Equation(s):
// \Mux51~10_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[21][12]~q )) # (!cuifregT_2 & ((\registerArray[17][12]~q )))))

	.dataa(\registerArray[21][12]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[17][12]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux51~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~10 .lut_mask = 16'hEE30;
defparam \Mux51~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N12
cycloneive_lcell_comb \Mux51~11 (
// Equation(s):
// \Mux51~11_combout  = (cuifregT_3 & ((\Mux51~10_combout  & (\registerArray[29][12]~q )) # (!\Mux51~10_combout  & ((\registerArray[25][12]~q ))))) # (!cuifregT_3 & (((\Mux51~10_combout ))))

	.dataa(\registerArray[29][12]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[25][12]~q ),
	.datad(\Mux51~10_combout ),
	.cin(gnd),
	.combout(\Mux51~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~11 .lut_mask = 16'hBBC0;
defparam \Mux51~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y33_N23
dffeas \registerArray[30][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][12] .is_wysiwyg = "true";
defparam \registerArray[30][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N22
cycloneive_lcell_comb \registerArray[26][12]~feeder (
// Equation(s):
// \registerArray[26][12]~feeder_combout  = \Mux56~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux562),
	.cin(gnd),
	.combout(\registerArray[26][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[26][12]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[26][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N23
dffeas \registerArray[26][12] (
	.clk(clk),
	.d(\registerArray[26][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][12] .is_wysiwyg = "true";
defparam \registerArray[26][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N17
dffeas \registerArray[18][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][12] .is_wysiwyg = "true";
defparam \registerArray[18][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N16
cycloneive_lcell_comb \Mux51~12 (
// Equation(s):
// \Mux51~12_combout  = (cuifregT_3 & ((\registerArray[26][12]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[18][12]~q  & !cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[26][12]~q ),
	.datac(\registerArray[18][12]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux51~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~12 .lut_mask = 16'hAAD8;
defparam \Mux51~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N22
cycloneive_lcell_comb \Mux51~13 (
// Equation(s):
// \Mux51~13_combout  = (cuifregT_2 & ((\Mux51~12_combout  & ((\registerArray[30][12]~q ))) # (!\Mux51~12_combout  & (\registerArray[22][12]~q )))) # (!cuifregT_2 & (((\Mux51~12_combout ))))

	.dataa(\registerArray[22][12]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[30][12]~q ),
	.datad(\Mux51~12_combout ),
	.cin(gnd),
	.combout(\Mux51~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~13 .lut_mask = 16'hF388;
defparam \Mux51~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N21
dffeas \registerArray[20][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][12] .is_wysiwyg = "true";
defparam \registerArray[20][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N31
dffeas \registerArray[28][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][12] .is_wysiwyg = "true";
defparam \registerArray[28][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N10
cycloneive_lcell_comb \registerArray[16][12]~feeder (
// Equation(s):
// \registerArray[16][12]~feeder_combout  = \Mux56~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux562),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[16][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[16][12]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[16][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N11
dffeas \registerArray[16][12] (
	.clk(clk),
	.d(\registerArray[16][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][12] .is_wysiwyg = "true";
defparam \registerArray[16][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N16
cycloneive_lcell_comb \Mux51~14 (
// Equation(s):
// \Mux51~14_combout  = (cuifregT_3 & ((\registerArray[24][12]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[16][12]~q  & !cuifregT_2))))

	.dataa(\registerArray[24][12]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[16][12]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux51~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~14 .lut_mask = 16'hCCB8;
defparam \Mux51~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N30
cycloneive_lcell_comb \Mux51~15 (
// Equation(s):
// \Mux51~15_combout  = (cuifregT_2 & ((\Mux51~14_combout  & ((\registerArray[28][12]~q ))) # (!\Mux51~14_combout  & (\registerArray[20][12]~q )))) # (!cuifregT_2 & (((\Mux51~14_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[20][12]~q ),
	.datac(\registerArray[28][12]~q ),
	.datad(\Mux51~14_combout ),
	.cin(gnd),
	.combout(\Mux51~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~15 .lut_mask = 16'hF588;
defparam \Mux51~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y34_N14
cycloneive_lcell_comb \Mux51~16 (
// Equation(s):
// \Mux51~16_combout  = (cuifregT_1 & ((cuifregT_01) # ((\Mux51~13_combout )))) # (!cuifregT_1 & (!cuifregT_01 & ((\Mux51~15_combout ))))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\Mux51~13_combout ),
	.datad(\Mux51~15_combout ),
	.cin(gnd),
	.combout(\Mux51~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~16 .lut_mask = 16'hB9A8;
defparam \Mux51~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N12
cycloneive_lcell_comb \registerArray[27][12]~feeder (
// Equation(s):
// \registerArray[27][12]~feeder_combout  = \Mux56~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux562),
	.cin(gnd),
	.combout(\registerArray[27][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[27][12]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[27][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N13
dffeas \registerArray[27][12] (
	.clk(clk),
	.d(\registerArray[27][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][12] .is_wysiwyg = "true";
defparam \registerArray[27][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N27
dffeas \registerArray[31][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][12] .is_wysiwyg = "true";
defparam \registerArray[31][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N25
dffeas \registerArray[19][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][12] .is_wysiwyg = "true";
defparam \registerArray[19][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N12
cycloneive_lcell_comb \registerArray[23][12]~feeder (
// Equation(s):
// \registerArray[23][12]~feeder_combout  = \Mux56~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux562),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[23][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[23][12]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[23][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y42_N13
dffeas \registerArray[23][12] (
	.clk(clk),
	.d(\registerArray[23][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][12] .is_wysiwyg = "true";
defparam \registerArray[23][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N24
cycloneive_lcell_comb \Mux51~17 (
// Equation(s):
// \Mux51~17_combout  = (cuifregT_3 & (cuifregT_2)) # (!cuifregT_3 & ((cuifregT_2 & ((\registerArray[23][12]~q ))) # (!cuifregT_2 & (\registerArray[19][12]~q ))))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\registerArray[19][12]~q ),
	.datad(\registerArray[23][12]~q ),
	.cin(gnd),
	.combout(\Mux51~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~17 .lut_mask = 16'hDC98;
defparam \Mux51~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N26
cycloneive_lcell_comb \Mux51~18 (
// Equation(s):
// \Mux51~18_combout  = (cuifregT_3 & ((\Mux51~17_combout  & ((\registerArray[31][12]~q ))) # (!\Mux51~17_combout  & (\registerArray[27][12]~q )))) # (!cuifregT_3 & (((\Mux51~17_combout ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[27][12]~q ),
	.datac(\registerArray[31][12]~q ),
	.datad(\Mux51~17_combout ),
	.cin(gnd),
	.combout(\Mux51~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~18 .lut_mask = 16'hF588;
defparam \Mux51~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N27
dffeas \registerArray[12][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][11] .is_wysiwyg = "true";
defparam \registerArray[12][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N26
cycloneive_lcell_comb \Mux52~7 (
// Equation(s):
// \Mux52~7_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[13][11]~q )) # (!cuifregT_01 & ((\registerArray[12][11]~q )))))

	.dataa(\registerArray[13][11]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[12][11]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux52~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~7 .lut_mask = 16'hEE30;
defparam \Mux52~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N21
dffeas \registerArray[15][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][11] .is_wysiwyg = "true";
defparam \registerArray[15][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N19
dffeas \registerArray[14][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][11] .is_wysiwyg = "true";
defparam \registerArray[14][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N20
cycloneive_lcell_comb \Mux52~8 (
// Equation(s):
// \Mux52~8_combout  = (\Mux52~7_combout  & (((\registerArray[15][11]~q )) # (!cuifregT_1))) # (!\Mux52~7_combout  & (cuifregT_1 & ((\registerArray[14][11]~q ))))

	.dataa(\Mux52~7_combout ),
	.datab(cuifregT_1),
	.datac(\registerArray[15][11]~q ),
	.datad(\registerArray[14][11]~q ),
	.cin(gnd),
	.combout(\Mux52~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~8 .lut_mask = 16'hE6A2;
defparam \Mux52~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y40_N7
dffeas \registerArray[2][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][11] .is_wysiwyg = "true";
defparam \registerArray[2][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N18
cycloneive_lcell_comb \registerArray[3][11]~feeder (
// Equation(s):
// \registerArray[3][11]~feeder_combout  = \Mux57~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux572),
	.cin(gnd),
	.combout(\registerArray[3][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[3][11]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[3][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y39_N19
dffeas \registerArray[3][11] (
	.clk(clk),
	.d(\registerArray[3][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][11] .is_wysiwyg = "true";
defparam \registerArray[3][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y40_N21
dffeas \registerArray[1][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][11] .is_wysiwyg = "true";
defparam \registerArray[1][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N20
cycloneive_lcell_comb \Mux52~4 (
// Equation(s):
// \Mux52~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][11]~q )) # (!cuifregT_1 & ((\registerArray[1][11]~q )))))

	.dataa(cuifregT_0),
	.datab(\registerArray[3][11]~q ),
	.datac(\registerArray[1][11]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux52~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~4 .lut_mask = 16'h88A0;
defparam \Mux52~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N6
cycloneive_lcell_comb \Mux52~5 (
// Equation(s):
// \Mux52~5_combout  = (\Mux52~4_combout ) # ((!cuifregT_01 & (cuifregT_1 & \registerArray[2][11]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[2][11]~q ),
	.datad(\Mux52~4_combout ),
	.cin(gnd),
	.combout(\Mux52~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~5 .lut_mask = 16'hFF40;
defparam \Mux52~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y43_N15
dffeas \registerArray[11][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][11] .is_wysiwyg = "true";
defparam \registerArray[11][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y43_N21
dffeas \registerArray[8][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][11] .is_wysiwyg = "true";
defparam \registerArray[8][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N20
cycloneive_lcell_comb \Mux52~2 (
// Equation(s):
// \Mux52~2_combout  = (cuifregT_1 & ((\registerArray[10][11]~q ) # ((cuifregT_01)))) # (!cuifregT_1 & (((\registerArray[8][11]~q  & !cuifregT_01))))

	.dataa(\registerArray[10][11]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[8][11]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux52~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~2 .lut_mask = 16'hCCB8;
defparam \Mux52~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y43_N14
cycloneive_lcell_comb \Mux52~3 (
// Equation(s):
// \Mux52~3_combout  = (cuifregT_01 & ((\Mux52~2_combout  & ((\registerArray[11][11]~q ))) # (!\Mux52~2_combout  & (\registerArray[9][11]~q )))) # (!cuifregT_01 & (((\Mux52~2_combout ))))

	.dataa(\registerArray[9][11]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[11][11]~q ),
	.datad(\Mux52~2_combout ),
	.cin(gnd),
	.combout(\Mux52~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~3 .lut_mask = 16'hF388;
defparam \Mux52~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N4
cycloneive_lcell_comb \Mux52~6 (
// Equation(s):
// \Mux52~6_combout  = (cuifregT_3 & ((cuifregT_2) # ((\Mux52~3_combout )))) # (!cuifregT_3 & (!cuifregT_2 & (\Mux52~5_combout )))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\Mux52~5_combout ),
	.datad(\Mux52~3_combout ),
	.cin(gnd),
	.combout(\Mux52~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~6 .lut_mask = 16'hBA98;
defparam \Mux52~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N13
dffeas \registerArray[5][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][11] .is_wysiwyg = "true";
defparam \registerArray[5][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N19
dffeas \registerArray[4][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][11] .is_wysiwyg = "true";
defparam \registerArray[4][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N18
cycloneive_lcell_comb \Mux52~0 (
// Equation(s):
// \Mux52~0_combout  = (cuifregT_01 & ((\registerArray[5][11]~q ) # ((cuifregT_1)))) # (!cuifregT_01 & (((\registerArray[4][11]~q  & !cuifregT_1))))

	.dataa(cuifregT_0),
	.datab(\registerArray[5][11]~q ),
	.datac(\registerArray[4][11]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux52~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~0 .lut_mask = 16'hAAD8;
defparam \Mux52~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N31
dffeas \registerArray[7][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][11] .is_wysiwyg = "true";
defparam \registerArray[7][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y38_N21
dffeas \registerArray[6][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][11] .is_wysiwyg = "true";
defparam \registerArray[6][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N30
cycloneive_lcell_comb \Mux52~1 (
// Equation(s):
// \Mux52~1_combout  = (\Mux52~0_combout  & (((\registerArray[7][11]~q )) # (!cuifregT_1))) # (!\Mux52~0_combout  & (cuifregT_1 & ((\registerArray[6][11]~q ))))

	.dataa(\Mux52~0_combout ),
	.datab(cuifregT_1),
	.datac(\registerArray[7][11]~q ),
	.datad(\registerArray[6][11]~q ),
	.cin(gnd),
	.combout(\Mux52~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~1 .lut_mask = 16'hE6A2;
defparam \Mux52~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N14
cycloneive_lcell_comb \registerArray[23][11]~feeder (
// Equation(s):
// \registerArray[23][11]~feeder_combout  = \Mux57~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux572),
	.cin(gnd),
	.combout(\registerArray[23][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[23][11]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[23][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y44_N15
dffeas \registerArray[23][11] (
	.clk(clk),
	.d(\registerArray[23][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][11] .is_wysiwyg = "true";
defparam \registerArray[23][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N23
dffeas \registerArray[31][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][11] .is_wysiwyg = "true";
defparam \registerArray[31][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N1
dffeas \registerArray[19][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][11] .is_wysiwyg = "true";
defparam \registerArray[19][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N8
cycloneive_lcell_comb \registerArray[27][11]~feeder (
// Equation(s):
// \registerArray[27][11]~feeder_combout  = \Mux57~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux572),
	.cin(gnd),
	.combout(\registerArray[27][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[27][11]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[27][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y44_N9
dffeas \registerArray[27][11] (
	.clk(clk),
	.d(\registerArray[27][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][11] .is_wysiwyg = "true";
defparam \registerArray[27][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N0
cycloneive_lcell_comb \Mux52~17 (
// Equation(s):
// \Mux52~17_combout  = (cuifregT_3 & ((cuifregT_2) # ((\registerArray[27][11]~q )))) # (!cuifregT_3 & (!cuifregT_2 & (\registerArray[19][11]~q )))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\registerArray[19][11]~q ),
	.datad(\registerArray[27][11]~q ),
	.cin(gnd),
	.combout(\Mux52~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~17 .lut_mask = 16'hBA98;
defparam \Mux52~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N22
cycloneive_lcell_comb \Mux52~18 (
// Equation(s):
// \Mux52~18_combout  = (cuifregT_2 & ((\Mux52~17_combout  & ((\registerArray[31][11]~q ))) # (!\Mux52~17_combout  & (\registerArray[23][11]~q )))) # (!cuifregT_2 & (((\Mux52~17_combout ))))

	.dataa(\registerArray[23][11]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[31][11]~q ),
	.datad(\Mux52~17_combout ),
	.cin(gnd),
	.combout(\Mux52~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~18 .lut_mask = 16'hF388;
defparam \Mux52~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N15
dffeas \registerArray[21][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][11] .is_wysiwyg = "true";
defparam \registerArray[21][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y31_N31
dffeas \registerArray[29][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][11] .is_wysiwyg = "true";
defparam \registerArray[29][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N26
cycloneive_lcell_comb \registerArray[17][11]~feeder (
// Equation(s):
// \registerArray[17][11]~feeder_combout  = \Mux57~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux572),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[17][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[17][11]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[17][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N27
dffeas \registerArray[17][11] (
	.clk(clk),
	.d(\registerArray[17][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][11] .is_wysiwyg = "true";
defparam \registerArray[17][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N1
dffeas \registerArray[25][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][11] .is_wysiwyg = "true";
defparam \registerArray[25][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N20
cycloneive_lcell_comb \Mux52~10 (
// Equation(s):
// \Mux52~10_combout  = (cuifregT_3 & (((\registerArray[25][11]~q ) # (cuifregT_2)))) # (!cuifregT_3 & (\registerArray[17][11]~q  & ((!cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[17][11]~q ),
	.datac(\registerArray[25][11]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux52~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~10 .lut_mask = 16'hAAE4;
defparam \Mux52~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N30
cycloneive_lcell_comb \Mux52~11 (
// Equation(s):
// \Mux52~11_combout  = (cuifregT_2 & ((\Mux52~10_combout  & ((\registerArray[29][11]~q ))) # (!\Mux52~10_combout  & (\registerArray[21][11]~q )))) # (!cuifregT_2 & (((\Mux52~10_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[21][11]~q ),
	.datac(\registerArray[29][11]~q ),
	.datad(\Mux52~10_combout ),
	.cin(gnd),
	.combout(\Mux52~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~11 .lut_mask = 16'hF588;
defparam \Mux52~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N5
dffeas \registerArray[26][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][11] .is_wysiwyg = "true";
defparam \registerArray[26][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N3
dffeas \registerArray[30][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][11] .is_wysiwyg = "true";
defparam \registerArray[30][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N23
dffeas \registerArray[22][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][11] .is_wysiwyg = "true";
defparam \registerArray[22][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N21
dffeas \registerArray[18][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][11] .is_wysiwyg = "true";
defparam \registerArray[18][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N20
cycloneive_lcell_comb \Mux52~12 (
// Equation(s):
// \Mux52~12_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[22][11]~q )) # (!cuifregT_2 & ((\registerArray[18][11]~q )))))

	.dataa(cuifregT_3),
	.datab(\registerArray[22][11]~q ),
	.datac(\registerArray[18][11]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux52~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~12 .lut_mask = 16'hEE50;
defparam \Mux52~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N2
cycloneive_lcell_comb \Mux52~13 (
// Equation(s):
// \Mux52~13_combout  = (cuifregT_3 & ((\Mux52~12_combout  & ((\registerArray[30][11]~q ))) # (!\Mux52~12_combout  & (\registerArray[26][11]~q )))) # (!cuifregT_3 & (((\Mux52~12_combout ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[26][11]~q ),
	.datac(\registerArray[30][11]~q ),
	.datad(\Mux52~12_combout ),
	.cin(gnd),
	.combout(\Mux52~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~13 .lut_mask = 16'hF588;
defparam \Mux52~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N19
dffeas \registerArray[28][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][11] .is_wysiwyg = "true";
defparam \registerArray[28][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y43_N15
dffeas \registerArray[20][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][11] .is_wysiwyg = "true";
defparam \registerArray[20][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N25
dffeas \registerArray[16][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][11] .is_wysiwyg = "true";
defparam \registerArray[16][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N24
cycloneive_lcell_comb \Mux52~14 (
// Equation(s):
// \Mux52~14_combout  = (cuifregT_2 & ((\registerArray[20][11]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[16][11]~q  & !cuifregT_3))))

	.dataa(cuifregT_2),
	.datab(\registerArray[20][11]~q ),
	.datac(\registerArray[16][11]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux52~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~14 .lut_mask = 16'hAAD8;
defparam \Mux52~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N18
cycloneive_lcell_comb \Mux52~15 (
// Equation(s):
// \Mux52~15_combout  = (cuifregT_3 & ((\Mux52~14_combout  & ((\registerArray[28][11]~q ))) # (!\Mux52~14_combout  & (\registerArray[24][11]~q )))) # (!cuifregT_3 & (((\Mux52~14_combout ))))

	.dataa(\registerArray[24][11]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[28][11]~q ),
	.datad(\Mux52~14_combout ),
	.cin(gnd),
	.combout(\Mux52~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~15 .lut_mask = 16'hF388;
defparam \Mux52~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N12
cycloneive_lcell_comb \Mux52~16 (
// Equation(s):
// \Mux52~16_combout  = (cuifregT_1 & ((cuifregT_01) # ((\Mux52~13_combout )))) # (!cuifregT_1 & (!cuifregT_01 & ((\Mux52~15_combout ))))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\Mux52~13_combout ),
	.datad(\Mux52~15_combout ),
	.cin(gnd),
	.combout(\Mux52~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~16 .lut_mask = 16'hB9A8;
defparam \Mux52~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N28
cycloneive_lcell_comb \registerArray[14][10]~feeder (
// Equation(s):
// \registerArray[14][10]~feeder_combout  = \Mux58~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux582),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[14][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][10]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[14][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y42_N29
dffeas \registerArray[14][10] (
	.clk(clk),
	.d(\registerArray[14][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][10] .is_wysiwyg = "true";
defparam \registerArray[14][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N7
dffeas \registerArray[15][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][10] .is_wysiwyg = "true";
defparam \registerArray[15][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N6
cycloneive_lcell_comb \registerArray[13][10]~feeder (
// Equation(s):
// \registerArray[13][10]~feeder_combout  = \Mux58~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux582),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[13][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[13][10]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[13][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y42_N7
dffeas \registerArray[13][10] (
	.clk(clk),
	.d(\registerArray[13][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][10] .is_wysiwyg = "true";
defparam \registerArray[13][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N12
cycloneive_lcell_comb \Mux53~7 (
// Equation(s):
// \Mux53~7_combout  = (cuifregT_01 & (((\registerArray[13][10]~q ) # (cuifregT_1)))) # (!cuifregT_01 & (\registerArray[12][10]~q  & ((!cuifregT_1))))

	.dataa(\registerArray[12][10]~q ),
	.datab(\registerArray[13][10]~q ),
	.datac(cuifregT_0),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux53~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~7 .lut_mask = 16'hF0CA;
defparam \Mux53~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N6
cycloneive_lcell_comb \Mux53~8 (
// Equation(s):
// \Mux53~8_combout  = (cuifregT_1 & ((\Mux53~7_combout  & ((\registerArray[15][10]~q ))) # (!\Mux53~7_combout  & (\registerArray[14][10]~q )))) # (!cuifregT_1 & (((\Mux53~7_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[14][10]~q ),
	.datac(\registerArray[15][10]~q ),
	.datad(\Mux53~7_combout ),
	.cin(gnd),
	.combout(\Mux53~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~8 .lut_mask = 16'hF588;
defparam \Mux53~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N29
dffeas \registerArray[9][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][10] .is_wysiwyg = "true";
defparam \registerArray[9][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N3
dffeas \registerArray[11][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][10] .is_wysiwyg = "true";
defparam \registerArray[11][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N1
dffeas \registerArray[8][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][10] .is_wysiwyg = "true";
defparam \registerArray[8][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N0
cycloneive_lcell_comb \Mux53~0 (
// Equation(s):
// \Mux53~0_combout  = (cuifregT_1 & ((\registerArray[10][10]~q ) # ((cuifregT_01)))) # (!cuifregT_1 & (((\registerArray[8][10]~q  & !cuifregT_01))))

	.dataa(\registerArray[10][10]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[8][10]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux53~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~0 .lut_mask = 16'hCCB8;
defparam \Mux53~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N2
cycloneive_lcell_comb \Mux53~1 (
// Equation(s):
// \Mux53~1_combout  = (cuifregT_01 & ((\Mux53~0_combout  & ((\registerArray[11][10]~q ))) # (!\Mux53~0_combout  & (\registerArray[9][10]~q )))) # (!cuifregT_01 & (((\Mux53~0_combout ))))

	.dataa(\registerArray[9][10]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[11][10]~q ),
	.datad(\Mux53~0_combout ),
	.cin(gnd),
	.combout(\Mux53~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~1 .lut_mask = 16'hF388;
defparam \Mux53~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N24
cycloneive_lcell_comb \registerArray[2][10]~feeder (
// Equation(s):
// \registerArray[2][10]~feeder_combout  = \Mux58~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux582),
	.cin(gnd),
	.combout(\registerArray[2][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[2][10]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[2][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y43_N25
dffeas \registerArray[2][10] (
	.clk(clk),
	.d(\registerArray[2][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][10] .is_wysiwyg = "true";
defparam \registerArray[2][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N4
cycloneive_lcell_comb \registerArray[1][10]~feeder (
// Equation(s):
// \registerArray[1][10]~feeder_combout  = \Mux58~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux582),
	.cin(gnd),
	.combout(\registerArray[1][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[1][10]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[1][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y43_N5
dffeas \registerArray[1][10] (
	.clk(clk),
	.d(\registerArray[1][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][10] .is_wysiwyg = "true";
defparam \registerArray[1][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N10
cycloneive_lcell_comb \Mux53~4 (
// Equation(s):
// \Mux53~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][10]~q )) # (!cuifregT_1 & ((\registerArray[1][10]~q )))))

	.dataa(\registerArray[3][10]~q ),
	.datab(\registerArray[1][10]~q ),
	.datac(cuifregT_1),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux53~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~4 .lut_mask = 16'hAC00;
defparam \Mux53~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N26
cycloneive_lcell_comb \Mux53~5 (
// Equation(s):
// \Mux53~5_combout  = (\Mux53~4_combout ) # ((cuifregT_1 & (\registerArray[2][10]~q  & !cuifregT_01)))

	.dataa(cuifregT_1),
	.datab(\registerArray[2][10]~q ),
	.datac(cuifregT_0),
	.datad(\Mux53~4_combout ),
	.cin(gnd),
	.combout(\Mux53~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~5 .lut_mask = 16'hFF08;
defparam \Mux53~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N6
cycloneive_lcell_comb \registerArray[6][10]~feeder (
// Equation(s):
// \registerArray[6][10]~feeder_combout  = \Mux58~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux582),
	.cin(gnd),
	.combout(\registerArray[6][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[6][10]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[6][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y43_N7
dffeas \registerArray[6][10] (
	.clk(clk),
	.d(\registerArray[6][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][10] .is_wysiwyg = "true";
defparam \registerArray[6][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N12
cycloneive_lcell_comb \registerArray[7][10]~feeder (
// Equation(s):
// \registerArray[7][10]~feeder_combout  = \Mux58~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux582),
	.cin(gnd),
	.combout(\registerArray[7][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[7][10]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[7][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y43_N13
dffeas \registerArray[7][10] (
	.clk(clk),
	.d(\registerArray[7][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][10] .is_wysiwyg = "true";
defparam \registerArray[7][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N15
dffeas \registerArray[4][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][10] .is_wysiwyg = "true";
defparam \registerArray[4][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N14
cycloneive_lcell_comb \Mux53~2 (
// Equation(s):
// \Mux53~2_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[5][10]~q )) # (!cuifregT_01 & ((\registerArray[4][10]~q )))))

	.dataa(\registerArray[5][10]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[4][10]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux53~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~2 .lut_mask = 16'hEE30;
defparam \Mux53~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N10
cycloneive_lcell_comb \Mux53~3 (
// Equation(s):
// \Mux53~3_combout  = (cuifregT_1 & ((\Mux53~2_combout  & ((\registerArray[7][10]~q ))) # (!\Mux53~2_combout  & (\registerArray[6][10]~q )))) # (!cuifregT_1 & (((\Mux53~2_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[6][10]~q ),
	.datac(\registerArray[7][10]~q ),
	.datad(\Mux53~2_combout ),
	.cin(gnd),
	.combout(\Mux53~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~3 .lut_mask = 16'hF588;
defparam \Mux53~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N0
cycloneive_lcell_comb \Mux53~6 (
// Equation(s):
// \Mux53~6_combout  = (cuifregT_3 & (cuifregT_2)) # (!cuifregT_3 & ((cuifregT_2 & ((\Mux53~3_combout ))) # (!cuifregT_2 & (\Mux53~5_combout ))))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\Mux53~5_combout ),
	.datad(\Mux53~3_combout ),
	.cin(gnd),
	.combout(\Mux53~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~6 .lut_mask = 16'hDC98;
defparam \Mux53~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N4
cycloneive_lcell_comb \registerArray[27][10]~feeder (
// Equation(s):
// \registerArray[27][10]~feeder_combout  = \Mux58~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux582),
	.cin(gnd),
	.combout(\registerArray[27][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[27][10]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[27][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y43_N5
dffeas \registerArray[27][10] (
	.clk(clk),
	.d(\registerArray[27][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][10] .is_wysiwyg = "true";
defparam \registerArray[27][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N3
dffeas \registerArray[31][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][10] .is_wysiwyg = "true";
defparam \registerArray[31][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N21
dffeas \registerArray[19][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][10] .is_wysiwyg = "true";
defparam \registerArray[19][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N20
cycloneive_lcell_comb \Mux53~17 (
// Equation(s):
// \Mux53~17_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[23][10]~q )) # (!cuifregT_2 & ((\registerArray[19][10]~q )))))

	.dataa(\registerArray[23][10]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[19][10]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux53~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~17 .lut_mask = 16'hEE30;
defparam \Mux53~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N2
cycloneive_lcell_comb \Mux53~18 (
// Equation(s):
// \Mux53~18_combout  = (cuifregT_3 & ((\Mux53~17_combout  & ((\registerArray[31][10]~q ))) # (!\Mux53~17_combout  & (\registerArray[27][10]~q )))) # (!cuifregT_3 & (((\Mux53~17_combout ))))

	.dataa(\registerArray[27][10]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[31][10]~q ),
	.datad(\Mux53~17_combout ),
	.cin(gnd),
	.combout(\Mux53~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~18 .lut_mask = 16'hF388;
defparam \Mux53~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N17
dffeas \registerArray[25][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][10] .is_wysiwyg = "true";
defparam \registerArray[25][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y40_N11
dffeas \registerArray[29][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][10] .is_wysiwyg = "true";
defparam \registerArray[29][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N14
cycloneive_lcell_comb \registerArray[17][10]~feeder (
// Equation(s):
// \registerArray[17][10]~feeder_combout  = \Mux58~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux582),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[17][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[17][10]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[17][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N15
dffeas \registerArray[17][10] (
	.clk(clk),
	.d(\registerArray[17][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][10] .is_wysiwyg = "true";
defparam \registerArray[17][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N22
cycloneive_lcell_comb \Mux53~10 (
// Equation(s):
// \Mux53~10_combout  = (cuifregT_2 & ((\registerArray[21][10]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[17][10]~q  & !cuifregT_3))))

	.dataa(\registerArray[21][10]~q ),
	.datab(\registerArray[17][10]~q ),
	.datac(cuifregT_2),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux53~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~10 .lut_mask = 16'hF0AC;
defparam \Mux53~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y40_N10
cycloneive_lcell_comb \Mux53~11 (
// Equation(s):
// \Mux53~11_combout  = (cuifregT_3 & ((\Mux53~10_combout  & ((\registerArray[29][10]~q ))) # (!\Mux53~10_combout  & (\registerArray[25][10]~q )))) # (!cuifregT_3 & (((\Mux53~10_combout ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[25][10]~q ),
	.datac(\registerArray[29][10]~q ),
	.datad(\Mux53~10_combout ),
	.cin(gnd),
	.combout(\Mux53~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~11 .lut_mask = 16'hF588;
defparam \Mux53~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y33_N27
dffeas \registerArray[30][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][10] .is_wysiwyg = "true";
defparam \registerArray[30][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N27
dffeas \registerArray[26][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][10] .is_wysiwyg = "true";
defparam \registerArray[26][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N1
dffeas \registerArray[18][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][10] .is_wysiwyg = "true";
defparam \registerArray[18][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N0
cycloneive_lcell_comb \Mux53~12 (
// Equation(s):
// \Mux53~12_combout  = (cuifregT_3 & ((\registerArray[26][10]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[18][10]~q  & !cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[26][10]~q ),
	.datac(\registerArray[18][10]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux53~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~12 .lut_mask = 16'hAAD8;
defparam \Mux53~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N26
cycloneive_lcell_comb \Mux53~13 (
// Equation(s):
// \Mux53~13_combout  = (cuifregT_2 & ((\Mux53~12_combout  & ((\registerArray[30][10]~q ))) # (!\Mux53~12_combout  & (\registerArray[22][10]~q )))) # (!cuifregT_2 & (((\Mux53~12_combout ))))

	.dataa(\registerArray[22][10]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[30][10]~q ),
	.datad(\Mux53~12_combout ),
	.cin(gnd),
	.combout(\Mux53~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~13 .lut_mask = 16'hF388;
defparam \Mux53~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N13
dffeas \registerArray[20][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][10] .is_wysiwyg = "true";
defparam \registerArray[20][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y39_N3
dffeas \registerArray[28][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][10] .is_wysiwyg = "true";
defparam \registerArray[28][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N14
cycloneive_lcell_comb \registerArray[16][10]~feeder (
// Equation(s):
// \registerArray[16][10]~feeder_combout  = \Mux58~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux582),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[16][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[16][10]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[16][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y39_N15
dffeas \registerArray[16][10] (
	.clk(clk),
	.d(\registerArray[16][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][10] .is_wysiwyg = "true";
defparam \registerArray[16][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N0
cycloneive_lcell_comb \Mux53~14 (
// Equation(s):
// \Mux53~14_combout  = (cuifregT_3 & ((\registerArray[24][10]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[16][10]~q  & !cuifregT_2))))

	.dataa(\registerArray[24][10]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[16][10]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux53~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~14 .lut_mask = 16'hCCB8;
defparam \Mux53~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N2
cycloneive_lcell_comb \Mux53~15 (
// Equation(s):
// \Mux53~15_combout  = (cuifregT_2 & ((\Mux53~14_combout  & ((\registerArray[28][10]~q ))) # (!\Mux53~14_combout  & (\registerArray[20][10]~q )))) # (!cuifregT_2 & (((\Mux53~14_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[20][10]~q ),
	.datac(\registerArray[28][10]~q ),
	.datad(\Mux53~14_combout ),
	.cin(gnd),
	.combout(\Mux53~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~15 .lut_mask = 16'hF588;
defparam \Mux53~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y43_N6
cycloneive_lcell_comb \Mux53~16 (
// Equation(s):
// \Mux53~16_combout  = (cuifregT_1 & ((cuifregT_01) # ((\Mux53~13_combout )))) # (!cuifregT_1 & (!cuifregT_01 & ((\Mux53~15_combout ))))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\Mux53~13_combout ),
	.datad(\Mux53~15_combout ),
	.cin(gnd),
	.combout(\Mux53~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~16 .lut_mask = 16'hB9A8;
defparam \Mux53~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N31
dffeas \registerArray[14][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][9] .is_wysiwyg = "true";
defparam \registerArray[14][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N9
dffeas \registerArray[12][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][9] .is_wysiwyg = "true";
defparam \registerArray[12][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N8
cycloneive_lcell_comb \Mux54~7 (
// Equation(s):
// \Mux54~7_combout  = (cuifregT_01 & ((\registerArray[13][9]~q ) # ((cuifregT_1)))) # (!cuifregT_01 & (((\registerArray[12][9]~q  & !cuifregT_1))))

	.dataa(\registerArray[13][9]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[12][9]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux54~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~7 .lut_mask = 16'hCCB8;
defparam \Mux54~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N15
dffeas \registerArray[15][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][9] .is_wysiwyg = "true";
defparam \registerArray[15][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N14
cycloneive_lcell_comb \Mux54~8 (
// Equation(s):
// \Mux54~8_combout  = (\Mux54~7_combout  & (((\registerArray[15][9]~q ) # (!cuifregT_1)))) # (!\Mux54~7_combout  & (\registerArray[14][9]~q  & ((cuifregT_1))))

	.dataa(\registerArray[14][9]~q ),
	.datab(\Mux54~7_combout ),
	.datac(\registerArray[15][9]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux54~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~8 .lut_mask = 16'hE2CC;
defparam \Mux54~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N9
dffeas \registerArray[6][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][9] .is_wysiwyg = "true";
defparam \registerArray[6][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N27
dffeas \registerArray[7][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][9] .is_wysiwyg = "true";
defparam \registerArray[7][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N1
dffeas \registerArray[5][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][9] .is_wysiwyg = "true";
defparam \registerArray[5][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N3
dffeas \registerArray[4][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][9] .is_wysiwyg = "true";
defparam \registerArray[4][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N2
cycloneive_lcell_comb \Mux54~0 (
// Equation(s):
// \Mux54~0_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[5][9]~q )) # (!cuifregT_01 & ((\registerArray[4][9]~q )))))

	.dataa(cuifregT_1),
	.datab(\registerArray[5][9]~q ),
	.datac(\registerArray[4][9]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux54~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~0 .lut_mask = 16'hEE50;
defparam \Mux54~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N26
cycloneive_lcell_comb \Mux54~1 (
// Equation(s):
// \Mux54~1_combout  = (cuifregT_1 & ((\Mux54~0_combout  & ((\registerArray[7][9]~q ))) # (!\Mux54~0_combout  & (\registerArray[6][9]~q )))) # (!cuifregT_1 & (((\Mux54~0_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[6][9]~q ),
	.datac(\registerArray[7][9]~q ),
	.datad(\Mux54~0_combout ),
	.cin(gnd),
	.combout(\Mux54~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~1 .lut_mask = 16'hF588;
defparam \Mux54~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N24
cycloneive_lcell_comb \registerArray[2][9]~feeder (
// Equation(s):
// \registerArray[2][9]~feeder_combout  = \Mux59~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux592),
	.cin(gnd),
	.combout(\registerArray[2][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[2][9]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[2][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N25
dffeas \registerArray[2][9] (
	.clk(clk),
	.d(\registerArray[2][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][9] .is_wysiwyg = "true";
defparam \registerArray[2][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N28
cycloneive_lcell_comb \registerArray[1][9]~feeder (
// Equation(s):
// \registerArray[1][9]~feeder_combout  = \Mux59~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux592),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[1][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[1][9]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[1][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y42_N29
dffeas \registerArray[1][9] (
	.clk(clk),
	.d(\registerArray[1][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][9] .is_wysiwyg = "true";
defparam \registerArray[1][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N4
cycloneive_lcell_comb \Mux54~4 (
// Equation(s):
// \Mux54~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][9]~q )) # (!cuifregT_1 & ((\registerArray[1][9]~q )))))

	.dataa(\registerArray[3][9]~q ),
	.datab(\registerArray[1][9]~q ),
	.datac(cuifregT_1),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux54~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~4 .lut_mask = 16'hAC00;
defparam \Mux54~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N30
cycloneive_lcell_comb \Mux54~5 (
// Equation(s):
// \Mux54~5_combout  = (\Mux54~4_combout ) # ((cuifregT_1 & (\registerArray[2][9]~q  & !cuifregT_01)))

	.dataa(cuifregT_1),
	.datab(\registerArray[2][9]~q ),
	.datac(\Mux54~4_combout ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux54~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~5 .lut_mask = 16'hF0F8;
defparam \Mux54~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N21
dffeas \registerArray[9][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][9] .is_wysiwyg = "true";
defparam \registerArray[9][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N15
dffeas \registerArray[11][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][9] .is_wysiwyg = "true";
defparam \registerArray[11][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N29
dffeas \registerArray[8][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][9] .is_wysiwyg = "true";
defparam \registerArray[8][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N28
cycloneive_lcell_comb \Mux54~2 (
// Equation(s):
// \Mux54~2_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & (\registerArray[10][9]~q )) # (!cuifregT_1 & ((\registerArray[8][9]~q )))))

	.dataa(\registerArray[10][9]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[8][9]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux54~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~2 .lut_mask = 16'hEE30;
defparam \Mux54~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N14
cycloneive_lcell_comb \Mux54~3 (
// Equation(s):
// \Mux54~3_combout  = (cuifregT_01 & ((\Mux54~2_combout  & ((\registerArray[11][9]~q ))) # (!\Mux54~2_combout  & (\registerArray[9][9]~q )))) # (!cuifregT_01 & (((\Mux54~2_combout ))))

	.dataa(cuifregT_0),
	.datab(\registerArray[9][9]~q ),
	.datac(\registerArray[11][9]~q ),
	.datad(\Mux54~2_combout ),
	.cin(gnd),
	.combout(\Mux54~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~3 .lut_mask = 16'hF588;
defparam \Mux54~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N20
cycloneive_lcell_comb \Mux54~6 (
// Equation(s):
// \Mux54~6_combout  = (cuifregT_2 & (cuifregT_3)) # (!cuifregT_2 & ((cuifregT_3 & ((\Mux54~3_combout ))) # (!cuifregT_3 & (\Mux54~5_combout ))))

	.dataa(cuifregT_2),
	.datab(cuifregT_3),
	.datac(\Mux54~5_combout ),
	.datad(\Mux54~3_combout ),
	.cin(gnd),
	.combout(\Mux54~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~6 .lut_mask = 16'hDC98;
defparam \Mux54~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N25
dffeas \registerArray[24][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][9] .is_wysiwyg = "true";
defparam \registerArray[24][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N13
dffeas \registerArray[28][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][9] .is_wysiwyg = "true";
defparam \registerArray[28][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N12
cycloneive_lcell_comb \Mux54~15 (
// Equation(s):
// \Mux54~15_combout  = (\Mux54~14_combout  & (((\registerArray[28][9]~q ) # (!cuifregT_3)))) # (!\Mux54~14_combout  & (\registerArray[24][9]~q  & ((cuifregT_3))))

	.dataa(\Mux54~14_combout ),
	.datab(\registerArray[24][9]~q ),
	.datac(\registerArray[28][9]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux54~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~15 .lut_mask = 16'hE4AA;
defparam \Mux54~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N19
dffeas \registerArray[22][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][9] .is_wysiwyg = "true";
defparam \registerArray[22][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N9
dffeas \registerArray[18][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][9] .is_wysiwyg = "true";
defparam \registerArray[18][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N8
cycloneive_lcell_comb \Mux54~12 (
// Equation(s):
// \Mux54~12_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[22][9]~q )) # (!cuifregT_2 & ((\registerArray[18][9]~q )))))

	.dataa(cuifregT_3),
	.datab(\registerArray[22][9]~q ),
	.datac(\registerArray[18][9]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux54~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~12 .lut_mask = 16'hEE50;
defparam \Mux54~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y33_N19
dffeas \registerArray[30][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][9] .is_wysiwyg = "true";
defparam \registerArray[30][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N1
dffeas \registerArray[26][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][9] .is_wysiwyg = "true";
defparam \registerArray[26][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N18
cycloneive_lcell_comb \Mux54~13 (
// Equation(s):
// \Mux54~13_combout  = (cuifregT_3 & ((\Mux54~12_combout  & (\registerArray[30][9]~q )) # (!\Mux54~12_combout  & ((\registerArray[26][9]~q ))))) # (!cuifregT_3 & (\Mux54~12_combout ))

	.dataa(cuifregT_3),
	.datab(\Mux54~12_combout ),
	.datac(\registerArray[30][9]~q ),
	.datad(\registerArray[26][9]~q ),
	.cin(gnd),
	.combout(\Mux54~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~13 .lut_mask = 16'hE6C4;
defparam \Mux54~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N22
cycloneive_lcell_comb \Mux54~16 (
// Equation(s):
// \Mux54~16_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & ((\Mux54~13_combout ))) # (!cuifregT_1 & (\Mux54~15_combout ))))

	.dataa(\Mux54~15_combout ),
	.datab(cuifregT_0),
	.datac(cuifregT_1),
	.datad(\Mux54~13_combout ),
	.cin(gnd),
	.combout(\Mux54~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~16 .lut_mask = 16'hF2C2;
defparam \Mux54~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N17
dffeas \registerArray[21][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][9] .is_wysiwyg = "true";
defparam \registerArray[21][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N8
cycloneive_lcell_comb \registerArray[29][9]~feeder (
// Equation(s):
// \registerArray[29][9]~feeder_combout  = \Mux59~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux592),
	.cin(gnd),
	.combout(\registerArray[29][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[29][9]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[29][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y30_N9
dffeas \registerArray[29][9] (
	.clk(clk),
	.d(\registerArray[29][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][9] .is_wysiwyg = "true";
defparam \registerArray[29][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N28
cycloneive_lcell_comb \registerArray[25][9]~feeder (
// Equation(s):
// \registerArray[25][9]~feeder_combout  = \Mux59~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux592),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[25][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[25][9]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[25][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N29
dffeas \registerArray[25][9] (
	.clk(clk),
	.d(\registerArray[25][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][9] .is_wysiwyg = "true";
defparam \registerArray[25][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N23
dffeas \registerArray[17][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][9] .is_wysiwyg = "true";
defparam \registerArray[17][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N22
cycloneive_lcell_comb \Mux54~10 (
// Equation(s):
// \Mux54~10_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[25][9]~q )) # (!cuifregT_3 & ((\registerArray[17][9]~q )))))

	.dataa(cuifregT_2),
	.datab(\registerArray[25][9]~q ),
	.datac(\registerArray[17][9]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux54~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~10 .lut_mask = 16'hEE50;
defparam \Mux54~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N10
cycloneive_lcell_comb \Mux54~11 (
// Equation(s):
// \Mux54~11_combout  = (cuifregT_2 & ((\Mux54~10_combout  & ((\registerArray[29][9]~q ))) # (!\Mux54~10_combout  & (\registerArray[21][9]~q )))) # (!cuifregT_2 & (((\Mux54~10_combout ))))

	.dataa(\registerArray[21][9]~q ),
	.datab(\registerArray[29][9]~q ),
	.datac(cuifregT_2),
	.datad(\Mux54~10_combout ),
	.cin(gnd),
	.combout(\Mux54~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~11 .lut_mask = 16'hCFA0;
defparam \Mux54~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N25
dffeas \registerArray[23][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][9] .is_wysiwyg = "true";
defparam \registerArray[23][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N11
dffeas \registerArray[31][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][9] .is_wysiwyg = "true";
defparam \registerArray[31][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N25
dffeas \registerArray[19][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][9] .is_wysiwyg = "true";
defparam \registerArray[19][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N24
cycloneive_lcell_comb \Mux54~17 (
// Equation(s):
// \Mux54~17_combout  = (cuifregT_3 & ((\registerArray[27][9]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[19][9]~q  & !cuifregT_2))))

	.dataa(\registerArray[27][9]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[19][9]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux54~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~17 .lut_mask = 16'hCCB8;
defparam \Mux54~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N10
cycloneive_lcell_comb \Mux54~18 (
// Equation(s):
// \Mux54~18_combout  = (cuifregT_2 & ((\Mux54~17_combout  & ((\registerArray[31][9]~q ))) # (!\Mux54~17_combout  & (\registerArray[23][9]~q )))) # (!cuifregT_2 & (((\Mux54~17_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[23][9]~q ),
	.datac(\registerArray[31][9]~q ),
	.datad(\Mux54~17_combout ),
	.cin(gnd),
	.combout(\Mux54~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~18 .lut_mask = 16'hF588;
defparam \Mux54~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N9
dffeas \registerArray[9][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][8] .is_wysiwyg = "true";
defparam \registerArray[9][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N5
dffeas \registerArray[8][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][8] .is_wysiwyg = "true";
defparam \registerArray[8][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N4
cycloneive_lcell_comb \Mux55~0 (
// Equation(s):
// \Mux55~0_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & (\registerArray[10][8]~q )) # (!cuifregT_1 & ((\registerArray[8][8]~q )))))

	.dataa(\registerArray[10][8]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[8][8]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux55~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~0 .lut_mask = 16'hEE30;
defparam \Mux55~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y31_N7
dffeas \registerArray[11][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][8] .is_wysiwyg = "true";
defparam \registerArray[11][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N6
cycloneive_lcell_comb \Mux55~1 (
// Equation(s):
// \Mux55~1_combout  = (\Mux55~0_combout  & (((\registerArray[11][8]~q ) # (!cuifregT_01)))) # (!\Mux55~0_combout  & (\registerArray[9][8]~q  & ((cuifregT_01))))

	.dataa(\registerArray[9][8]~q ),
	.datab(\Mux55~0_combout ),
	.datac(\registerArray[11][8]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux55~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~1 .lut_mask = 16'hE2CC;
defparam \Mux55~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N10
cycloneive_lcell_comb \registerArray[14][8]~feeder (
// Equation(s):
// \registerArray[14][8]~feeder_combout  = \Mux60~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux602),
	.cin(gnd),
	.combout(\registerArray[14][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][8]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[14][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N11
dffeas \registerArray[14][8] (
	.clk(clk),
	.d(\registerArray[14][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][8] .is_wysiwyg = "true";
defparam \registerArray[14][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N27
dffeas \registerArray[15][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][8] .is_wysiwyg = "true";
defparam \registerArray[15][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N17
dffeas \registerArray[12][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][8] .is_wysiwyg = "true";
defparam \registerArray[12][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N16
cycloneive_lcell_comb \Mux55~7 (
// Equation(s):
// \Mux55~7_combout  = (cuifregT_01 & ((\registerArray[13][8]~q ) # ((cuifregT_1)))) # (!cuifregT_01 & (((\registerArray[12][8]~q  & !cuifregT_1))))

	.dataa(\registerArray[13][8]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[12][8]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux55~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~7 .lut_mask = 16'hCCB8;
defparam \Mux55~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N26
cycloneive_lcell_comb \Mux55~8 (
// Equation(s):
// \Mux55~8_combout  = (cuifregT_1 & ((\Mux55~7_combout  & ((\registerArray[15][8]~q ))) # (!\Mux55~7_combout  & (\registerArray[14][8]~q )))) # (!cuifregT_1 & (((\Mux55~7_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[14][8]~q ),
	.datac(\registerArray[15][8]~q ),
	.datad(\Mux55~7_combout ),
	.cin(gnd),
	.combout(\Mux55~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~8 .lut_mask = 16'hF588;
defparam \Mux55~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N2
cycloneive_lcell_comb \registerArray[6][8]~feeder (
// Equation(s):
// \registerArray[6][8]~feeder_combout  = \Mux60~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux602),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[6][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[6][8]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[6][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y30_N3
dffeas \registerArray[6][8] (
	.clk(clk),
	.d(\registerArray[6][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][8] .is_wysiwyg = "true";
defparam \registerArray[6][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N15
dffeas \registerArray[7][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][8] .is_wysiwyg = "true";
defparam \registerArray[7][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N21
dffeas \registerArray[4][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][8] .is_wysiwyg = "true";
defparam \registerArray[4][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N20
cycloneive_lcell_comb \Mux55~2 (
// Equation(s):
// \Mux55~2_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[5][8]~q )) # (!cuifregT_01 & ((\registerArray[4][8]~q )))))

	.dataa(\registerArray[5][8]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[4][8]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux55~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~2 .lut_mask = 16'hEE30;
defparam \Mux55~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N14
cycloneive_lcell_comb \Mux55~3 (
// Equation(s):
// \Mux55~3_combout  = (cuifregT_1 & ((\Mux55~2_combout  & ((\registerArray[7][8]~q ))) # (!\Mux55~2_combout  & (\registerArray[6][8]~q )))) # (!cuifregT_1 & (((\Mux55~2_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[6][8]~q ),
	.datac(\registerArray[7][8]~q ),
	.datad(\Mux55~2_combout ),
	.cin(gnd),
	.combout(\Mux55~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~3 .lut_mask = 16'hF588;
defparam \Mux55~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y37_N7
dffeas \registerArray[2][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][8] .is_wysiwyg = "true";
defparam \registerArray[2][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y37_N21
dffeas \registerArray[1][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][8] .is_wysiwyg = "true";
defparam \registerArray[1][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N20
cycloneive_lcell_comb \Mux55~4 (
// Equation(s):
// \Mux55~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][8]~q )) # (!cuifregT_1 & ((\registerArray[1][8]~q )))))

	.dataa(\registerArray[3][8]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[1][8]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux55~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~4 .lut_mask = 16'hB800;
defparam \Mux55~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N6
cycloneive_lcell_comb \Mux55~5 (
// Equation(s):
// \Mux55~5_combout  = (\Mux55~4_combout ) # ((!cuifregT_01 & (cuifregT_1 & \registerArray[2][8]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[2][8]~q ),
	.datad(\Mux55~4_combout ),
	.cin(gnd),
	.combout(\Mux55~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~5 .lut_mask = 16'hFF40;
defparam \Mux55~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N0
cycloneive_lcell_comb \Mux55~6 (
// Equation(s):
// \Mux55~6_combout  = (cuifregT_3 & (cuifregT_2)) # (!cuifregT_3 & ((cuifregT_2 & (\Mux55~3_combout )) # (!cuifregT_2 & ((\Mux55~5_combout )))))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\Mux55~3_combout ),
	.datad(\Mux55~5_combout ),
	.cin(gnd),
	.combout(\Mux55~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~6 .lut_mask = 16'hD9C8;
defparam \Mux55~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N18
cycloneive_lcell_comb \registerArray[19][8]~feeder (
// Equation(s):
// \registerArray[19][8]~feeder_combout  = \Mux60~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux602),
	.cin(gnd),
	.combout(\registerArray[19][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[19][8]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[19][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y30_N19
dffeas \registerArray[19][8] (
	.clk(clk),
	.d(\registerArray[19][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][8] .is_wysiwyg = "true";
defparam \registerArray[19][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N2
cycloneive_lcell_comb \registerArray[23][8]~feeder (
// Equation(s):
// \registerArray[23][8]~feeder_combout  = \Mux60~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux602),
	.cin(gnd),
	.combout(\registerArray[23][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[23][8]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[23][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N3
dffeas \registerArray[23][8] (
	.clk(clk),
	.d(\registerArray[23][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][8] .is_wysiwyg = "true";
defparam \registerArray[23][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N30
cycloneive_lcell_comb \Mux55~17 (
// Equation(s):
// \Mux55~17_combout  = (cuifregT_2 & (((\registerArray[23][8]~q ) # (cuifregT_3)))) # (!cuifregT_2 & (\registerArray[19][8]~q  & ((!cuifregT_3))))

	.dataa(cuifregT_2),
	.datab(\registerArray[19][8]~q ),
	.datac(\registerArray[23][8]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux55~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~17 .lut_mask = 16'hAAE4;
defparam \Mux55~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N1
dffeas \registerArray[27][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][8] .is_wysiwyg = "true";
defparam \registerArray[27][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N25
dffeas \registerArray[31][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][8] .is_wysiwyg = "true";
defparam \registerArray[31][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N24
cycloneive_lcell_comb \Mux55~18 (
// Equation(s):
// \Mux55~18_combout  = (\Mux55~17_combout  & (((\registerArray[31][8]~q ) # (!cuifregT_3)))) # (!\Mux55~17_combout  & (\registerArray[27][8]~q  & ((cuifregT_3))))

	.dataa(\Mux55~17_combout ),
	.datab(\registerArray[27][8]~q ),
	.datac(\registerArray[31][8]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux55~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~18 .lut_mask = 16'hE4AA;
defparam \Mux55~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y31_N31
dffeas \registerArray[30][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][8] .is_wysiwyg = "true";
defparam \registerArray[30][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N25
dffeas \registerArray[18][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][8] .is_wysiwyg = "true";
defparam \registerArray[18][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N24
cycloneive_lcell_comb \Mux55~12 (
// Equation(s):
// \Mux55~12_combout  = (cuifregT_3 & ((\registerArray[26][8]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[18][8]~q  & !cuifregT_2))))

	.dataa(\registerArray[26][8]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[18][8]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux55~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~12 .lut_mask = 16'hCCB8;
defparam \Mux55~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N30
cycloneive_lcell_comb \Mux55~13 (
// Equation(s):
// \Mux55~13_combout  = (cuifregT_2 & ((\Mux55~12_combout  & ((\registerArray[30][8]~q ))) # (!\Mux55~12_combout  & (\registerArray[22][8]~q )))) # (!cuifregT_2 & (((\Mux55~12_combout ))))

	.dataa(\registerArray[22][8]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[30][8]~q ),
	.datad(\Mux55~12_combout ),
	.cin(gnd),
	.combout(\Mux55~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~13 .lut_mask = 16'hF388;
defparam \Mux55~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N9
dffeas \registerArray[20][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][8] .is_wysiwyg = "true";
defparam \registerArray[20][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y35_N21
dffeas \registerArray[28][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][8] .is_wysiwyg = "true";
defparam \registerArray[28][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N20
cycloneive_lcell_comb \Mux55~15 (
// Equation(s):
// \Mux55~15_combout  = (\Mux55~14_combout  & (((\registerArray[28][8]~q ) # (!cuifregT_2)))) # (!\Mux55~14_combout  & (\registerArray[20][8]~q  & ((cuifregT_2))))

	.dataa(\Mux55~14_combout ),
	.datab(\registerArray[20][8]~q ),
	.datac(\registerArray[28][8]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux55~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~15 .lut_mask = 16'hE4AA;
defparam \Mux55~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y35_N2
cycloneive_lcell_comb \Mux55~16 (
// Equation(s):
// \Mux55~16_combout  = (cuifregT_1 & ((cuifregT_01) # ((\Mux55~13_combout )))) # (!cuifregT_1 & (!cuifregT_01 & ((\Mux55~15_combout ))))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\Mux55~13_combout ),
	.datad(\Mux55~15_combout ),
	.cin(gnd),
	.combout(\Mux55~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~16 .lut_mask = 16'hB9A8;
defparam \Mux55~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N12
cycloneive_lcell_comb \registerArray[29][8]~feeder (
// Equation(s):
// \registerArray[29][8]~feeder_combout  = \Mux60~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux602),
	.cin(gnd),
	.combout(\registerArray[29][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[29][8]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[29][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N13
dffeas \registerArray[29][8] (
	.clk(clk),
	.d(\registerArray[29][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][8] .is_wysiwyg = "true";
defparam \registerArray[29][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N8
cycloneive_lcell_comb \registerArray[25][8]~feeder (
// Equation(s):
// \registerArray[25][8]~feeder_combout  = \Mux60~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux602),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[25][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[25][8]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[25][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N9
dffeas \registerArray[25][8] (
	.clk(clk),
	.d(\registerArray[25][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][8] .is_wysiwyg = "true";
defparam \registerArray[25][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N20
cycloneive_lcell_comb \registerArray[17][8]~feeder (
// Equation(s):
// \registerArray[17][8]~feeder_combout  = \Mux60~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux602),
	.cin(gnd),
	.combout(\registerArray[17][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[17][8]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[17][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N21
dffeas \registerArray[17][8] (
	.clk(clk),
	.d(\registerArray[17][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][8] .is_wysiwyg = "true";
defparam \registerArray[17][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N18
cycloneive_lcell_comb \Mux55~10 (
// Equation(s):
// \Mux55~10_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[21][8]~q )) # (!cuifregT_2 & ((\registerArray[17][8]~q )))))

	.dataa(\registerArray[21][8]~q ),
	.datab(\registerArray[17][8]~q ),
	.datac(cuifregT_3),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux55~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~10 .lut_mask = 16'hFA0C;
defparam \Mux55~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N30
cycloneive_lcell_comb \Mux55~11 (
// Equation(s):
// \Mux55~11_combout  = (cuifregT_3 & ((\Mux55~10_combout  & (\registerArray[29][8]~q )) # (!\Mux55~10_combout  & ((\registerArray[25][8]~q ))))) # (!cuifregT_3 & (((\Mux55~10_combout ))))

	.dataa(\registerArray[29][8]~q ),
	.datab(\registerArray[25][8]~q ),
	.datac(cuifregT_3),
	.datad(\Mux55~10_combout ),
	.cin(gnd),
	.combout(\Mux55~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~11 .lut_mask = 16'hAFC0;
defparam \Mux55~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N18
cycloneive_lcell_comb \registerArray[14][7]~feeder (
// Equation(s):
// \registerArray[14][7]~feeder_combout  = \Mux61~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux612),
	.cin(gnd),
	.combout(\registerArray[14][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][7]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[14][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y39_N19
dffeas \registerArray[14][7] (
	.clk(clk),
	.d(\registerArray[14][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][7] .is_wysiwyg = "true";
defparam \registerArray[14][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N31
dffeas \registerArray[15][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][7] .is_wysiwyg = "true";
defparam \registerArray[15][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N5
dffeas \registerArray[13][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][7] .is_wysiwyg = "true";
defparam \registerArray[13][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y36_N9
dffeas \registerArray[12][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][7] .is_wysiwyg = "true";
defparam \registerArray[12][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N8
cycloneive_lcell_comb \Mux56~7 (
// Equation(s):
// \Mux56~7_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[13][7]~q )) # (!cuifregT_01 & ((\registerArray[12][7]~q )))))

	.dataa(cuifregT_1),
	.datab(\registerArray[13][7]~q ),
	.datac(\registerArray[12][7]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux56~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~7 .lut_mask = 16'hEE50;
defparam \Mux56~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y36_N30
cycloneive_lcell_comb \Mux56~8 (
// Equation(s):
// \Mux56~8_combout  = (cuifregT_1 & ((\Mux56~7_combout  & ((\registerArray[15][7]~q ))) # (!\Mux56~7_combout  & (\registerArray[14][7]~q )))) # (!cuifregT_1 & (((\Mux56~7_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[14][7]~q ),
	.datac(\registerArray[15][7]~q ),
	.datad(\Mux56~7_combout ),
	.cin(gnd),
	.combout(\Mux56~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~8 .lut_mask = 16'hF588;
defparam \Mux56~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N21
dffeas \registerArray[6][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][7] .is_wysiwyg = "true";
defparam \registerArray[6][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N13
dffeas \registerArray[7][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][7] .is_wysiwyg = "true";
defparam \registerArray[7][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N14
cycloneive_lcell_comb \registerArray[4][7]~feeder (
// Equation(s):
// \registerArray[4][7]~feeder_combout  = \Mux61~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux612),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[4][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[4][7]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[4][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N15
dffeas \registerArray[4][7] (
	.clk(clk),
	.d(\registerArray[4][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][7] .is_wysiwyg = "true";
defparam \registerArray[4][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N2
cycloneive_lcell_comb \Mux56~0 (
// Equation(s):
// \Mux56~0_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[5][7]~q )) # (!cuifregT_01 & ((\registerArray[4][7]~q )))))

	.dataa(\registerArray[5][7]~q ),
	.datab(\registerArray[4][7]~q ),
	.datac(cuifregT_1),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux56~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~0 .lut_mask = 16'hFA0C;
defparam \Mux56~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N12
cycloneive_lcell_comb \Mux56~1 (
// Equation(s):
// \Mux56~1_combout  = (cuifregT_1 & ((\Mux56~0_combout  & ((\registerArray[7][7]~q ))) # (!\Mux56~0_combout  & (\registerArray[6][7]~q )))) # (!cuifregT_1 & (((\Mux56~0_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[6][7]~q ),
	.datac(\registerArray[7][7]~q ),
	.datad(\Mux56~0_combout ),
	.cin(gnd),
	.combout(\Mux56~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~1 .lut_mask = 16'hF588;
defparam \Mux56~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y35_N9
dffeas \registerArray[2][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][7] .is_wysiwyg = "true";
defparam \registerArray[2][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N8
cycloneive_lcell_comb \Mux56~5 (
// Equation(s):
// \Mux56~5_combout  = (\Mux56~4_combout ) # ((cuifregT_1 & (\registerArray[2][7]~q  & !cuifregT_01)))

	.dataa(\Mux56~4_combout ),
	.datab(cuifregT_1),
	.datac(\registerArray[2][7]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux56~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~5 .lut_mask = 16'hAAEA;
defparam \Mux56~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y36_N11
dffeas \registerArray[11][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][7] .is_wysiwyg = "true";
defparam \registerArray[11][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y36_N29
dffeas \registerArray[8][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][7] .is_wysiwyg = "true";
defparam \registerArray[8][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N28
cycloneive_lcell_comb \Mux56~2 (
// Equation(s):
// \Mux56~2_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & (\registerArray[10][7]~q )) # (!cuifregT_1 & ((\registerArray[8][7]~q )))))

	.dataa(\registerArray[10][7]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[8][7]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux56~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~2 .lut_mask = 16'hEE30;
defparam \Mux56~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y36_N10
cycloneive_lcell_comb \Mux56~3 (
// Equation(s):
// \Mux56~3_combout  = (cuifregT_01 & ((\Mux56~2_combout  & ((\registerArray[11][7]~q ))) # (!\Mux56~2_combout  & (\registerArray[9][7]~q )))) # (!cuifregT_01 & (((\Mux56~2_combout ))))

	.dataa(\registerArray[9][7]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[11][7]~q ),
	.datad(\Mux56~2_combout ),
	.cin(gnd),
	.combout(\Mux56~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~3 .lut_mask = 16'hF388;
defparam \Mux56~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N6
cycloneive_lcell_comb \Mux56~6 (
// Equation(s):
// \Mux56~6_combout  = (cuifregT_2 & (cuifregT_3)) # (!cuifregT_2 & ((cuifregT_3 & ((\Mux56~3_combout ))) # (!cuifregT_3 & (\Mux56~5_combout ))))

	.dataa(cuifregT_2),
	.datab(cuifregT_3),
	.datac(\Mux56~5_combout ),
	.datad(\Mux56~3_combout ),
	.cin(gnd),
	.combout(\Mux56~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~6 .lut_mask = 16'hDC98;
defparam \Mux56~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N17
dffeas \registerArray[23][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][7] .is_wysiwyg = "true";
defparam \registerArray[23][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N15
dffeas \registerArray[31][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][7] .is_wysiwyg = "true";
defparam \registerArray[31][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y39_N29
dffeas \registerArray[19][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][7] .is_wysiwyg = "true";
defparam \registerArray[19][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N28
cycloneive_lcell_comb \Mux56~17 (
// Equation(s):
// \Mux56~17_combout  = (cuifregT_3 & ((\registerArray[27][7]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[19][7]~q  & !cuifregT_2))))

	.dataa(\registerArray[27][7]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[19][7]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux56~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~17 .lut_mask = 16'hCCB8;
defparam \Mux56~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N14
cycloneive_lcell_comb \Mux56~18 (
// Equation(s):
// \Mux56~18_combout  = (cuifregT_2 & ((\Mux56~17_combout  & ((\registerArray[31][7]~q ))) # (!\Mux56~17_combout  & (\registerArray[23][7]~q )))) # (!cuifregT_2 & (((\Mux56~17_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[23][7]~q ),
	.datac(\registerArray[31][7]~q ),
	.datad(\Mux56~17_combout ),
	.cin(gnd),
	.combout(\Mux56~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~18 .lut_mask = 16'hF588;
defparam \Mux56~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y30_N1
dffeas \registerArray[21][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][7] .is_wysiwyg = "true";
defparam \registerArray[21][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y31_N23
dffeas \registerArray[29][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][7] .is_wysiwyg = "true";
defparam \registerArray[29][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y30_N19
dffeas \registerArray[25][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][7] .is_wysiwyg = "true";
defparam \registerArray[25][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N5
dffeas \registerArray[17][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][7] .is_wysiwyg = "true";
defparam \registerArray[17][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N4
cycloneive_lcell_comb \Mux56~10 (
// Equation(s):
// \Mux56~10_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[25][7]~q )) # (!cuifregT_3 & ((\registerArray[17][7]~q )))))

	.dataa(cuifregT_2),
	.datab(\registerArray[25][7]~q ),
	.datac(\registerArray[17][7]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux56~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~10 .lut_mask = 16'hEE50;
defparam \Mux56~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N22
cycloneive_lcell_comb \Mux56~11 (
// Equation(s):
// \Mux56~11_combout  = (cuifregT_2 & ((\Mux56~10_combout  & ((\registerArray[29][7]~q ))) # (!\Mux56~10_combout  & (\registerArray[21][7]~q )))) # (!cuifregT_2 & (((\Mux56~10_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[21][7]~q ),
	.datac(\registerArray[29][7]~q ),
	.datad(\Mux56~10_combout ),
	.cin(gnd),
	.combout(\Mux56~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~11 .lut_mask = 16'hF588;
defparam \Mux56~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y32_N11
dffeas \registerArray[28][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][7] .is_wysiwyg = "true";
defparam \registerArray[28][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N21
dffeas \registerArray[16][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][7] .is_wysiwyg = "true";
defparam \registerArray[16][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N20
cycloneive_lcell_comb \Mux56~14 (
// Equation(s):
// \Mux56~14_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[20][7]~q )) # (!cuifregT_2 & ((\registerArray[16][7]~q )))))

	.dataa(\registerArray[20][7]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[16][7]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux56~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~14 .lut_mask = 16'hEE30;
defparam \Mux56~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N10
cycloneive_lcell_comb \Mux56~15 (
// Equation(s):
// \Mux56~15_combout  = (cuifregT_3 & ((\Mux56~14_combout  & ((\registerArray[28][7]~q ))) # (!\Mux56~14_combout  & (\registerArray[24][7]~q )))) # (!cuifregT_3 & (((\Mux56~14_combout ))))

	.dataa(\registerArray[24][7]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[28][7]~q ),
	.datad(\Mux56~14_combout ),
	.cin(gnd),
	.combout(\Mux56~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~15 .lut_mask = 16'hF388;
defparam \Mux56~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y31_N27
dffeas \registerArray[30][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][7] .is_wysiwyg = "true";
defparam \registerArray[30][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N17
dffeas \registerArray[18][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][7] .is_wysiwyg = "true";
defparam \registerArray[18][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N16
cycloneive_lcell_comb \Mux56~12 (
// Equation(s):
// \Mux56~12_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[22][7]~q )) # (!cuifregT_2 & ((\registerArray[18][7]~q )))))

	.dataa(\registerArray[22][7]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[18][7]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux56~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~12 .lut_mask = 16'hEE30;
defparam \Mux56~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N26
cycloneive_lcell_comb \Mux56~13 (
// Equation(s):
// \Mux56~13_combout  = (cuifregT_3 & ((\Mux56~12_combout  & ((\registerArray[30][7]~q ))) # (!\Mux56~12_combout  & (\registerArray[26][7]~q )))) # (!cuifregT_3 & (((\Mux56~12_combout ))))

	.dataa(\registerArray[26][7]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[30][7]~q ),
	.datad(\Mux56~12_combout ),
	.cin(gnd),
	.combout(\Mux56~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~13 .lut_mask = 16'hF388;
defparam \Mux56~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y35_N16
cycloneive_lcell_comb \Mux56~16 (
// Equation(s):
// \Mux56~16_combout  = (cuifregT_1 & ((cuifregT_01) # ((\Mux56~13_combout )))) # (!cuifregT_1 & (!cuifregT_01 & (\Mux56~15_combout )))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\Mux56~15_combout ),
	.datad(\Mux56~13_combout ),
	.cin(gnd),
	.combout(\Mux56~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~16 .lut_mask = 16'hBA98;
defparam \Mux56~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N25
dffeas \registerArray[9][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][6] .is_wysiwyg = "true";
defparam \registerArray[9][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N11
dffeas \registerArray[11][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][6] .is_wysiwyg = "true";
defparam \registerArray[11][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N21
dffeas \registerArray[8][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][6] .is_wysiwyg = "true";
defparam \registerArray[8][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N20
cycloneive_lcell_comb \Mux57~0 (
// Equation(s):
// \Mux57~0_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & (\registerArray[10][6]~q )) # (!cuifregT_1 & ((\registerArray[8][6]~q )))))

	.dataa(\registerArray[10][6]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[8][6]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux57~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~0 .lut_mask = 16'hEE30;
defparam \Mux57~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N10
cycloneive_lcell_comb \Mux57~1 (
// Equation(s):
// \Mux57~1_combout  = (cuifregT_01 & ((\Mux57~0_combout  & ((\registerArray[11][6]~q ))) # (!\Mux57~0_combout  & (\registerArray[9][6]~q )))) # (!cuifregT_01 & (((\Mux57~0_combout ))))

	.dataa(\registerArray[9][6]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[11][6]~q ),
	.datad(\Mux57~0_combout ),
	.cin(gnd),
	.combout(\Mux57~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~1 .lut_mask = 16'hF388;
defparam \Mux57~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y32_N9
dffeas \registerArray[2][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][6] .is_wysiwyg = "true";
defparam \registerArray[2][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N4
cycloneive_lcell_comb \registerArray[3][6]~feeder (
// Equation(s):
// \registerArray[3][6]~feeder_combout  = \Mux62~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux622),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[3][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[3][6]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[3][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y43_N5
dffeas \registerArray[3][6] (
	.clk(clk),
	.d(\registerArray[3][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][6] .is_wysiwyg = "true";
defparam \registerArray[3][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N19
dffeas \registerArray[1][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][6] .is_wysiwyg = "true";
defparam \registerArray[1][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N18
cycloneive_lcell_comb \Mux57~4 (
// Equation(s):
// \Mux57~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][6]~q )) # (!cuifregT_1 & ((\registerArray[1][6]~q )))))

	.dataa(cuifregT_1),
	.datab(\registerArray[3][6]~q ),
	.datac(\registerArray[1][6]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux57~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~4 .lut_mask = 16'hD800;
defparam \Mux57~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N8
cycloneive_lcell_comb \Mux57~5 (
// Equation(s):
// \Mux57~5_combout  = (\Mux57~4_combout ) # ((!cuifregT_01 & (cuifregT_1 & \registerArray[2][6]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[2][6]~q ),
	.datad(\Mux57~4_combout ),
	.cin(gnd),
	.combout(\Mux57~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~5 .lut_mask = 16'hFF40;
defparam \Mux57~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y32_N11
dffeas \registerArray[7][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][6] .is_wysiwyg = "true";
defparam \registerArray[7][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N4
cycloneive_lcell_comb \registerArray[5][6]~feeder (
// Equation(s):
// \registerArray[5][6]~feeder_combout  = \Mux62~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux622),
	.cin(gnd),
	.combout(\registerArray[5][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[5][6]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[5][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y30_N5
dffeas \registerArray[5][6] (
	.clk(clk),
	.d(\registerArray[5][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][6] .is_wysiwyg = "true";
defparam \registerArray[5][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N20
cycloneive_lcell_comb \Mux57~2 (
// Equation(s):
// \Mux57~2_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & ((\registerArray[5][6]~q ))) # (!cuifregT_01 & (\registerArray[4][6]~q ))))

	.dataa(\registerArray[4][6]~q ),
	.datab(\registerArray[5][6]~q ),
	.datac(cuifregT_1),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux57~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~2 .lut_mask = 16'hFC0A;
defparam \Mux57~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N10
cycloneive_lcell_comb \Mux57~3 (
// Equation(s):
// \Mux57~3_combout  = (cuifregT_1 & ((\Mux57~2_combout  & ((\registerArray[7][6]~q ))) # (!\Mux57~2_combout  & (\registerArray[6][6]~q )))) # (!cuifregT_1 & (((\Mux57~2_combout ))))

	.dataa(\registerArray[6][6]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[7][6]~q ),
	.datad(\Mux57~2_combout ),
	.cin(gnd),
	.combout(\Mux57~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~3 .lut_mask = 16'hF388;
defparam \Mux57~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N26
cycloneive_lcell_comb \Mux57~6 (
// Equation(s):
// \Mux57~6_combout  = (cuifregT_2 & ((cuifregT_3) # ((\Mux57~3_combout )))) # (!cuifregT_2 & (!cuifregT_3 & (\Mux57~5_combout )))

	.dataa(cuifregT_2),
	.datab(cuifregT_3),
	.datac(\Mux57~5_combout ),
	.datad(\Mux57~3_combout ),
	.cin(gnd),
	.combout(\Mux57~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~6 .lut_mask = 16'hBA98;
defparam \Mux57~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N13
dffeas \registerArray[14][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][6] .is_wysiwyg = "true";
defparam \registerArray[14][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N7
dffeas \registerArray[15][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][6] .is_wysiwyg = "true";
defparam \registerArray[15][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y38_N17
dffeas \registerArray[12][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][6] .is_wysiwyg = "true";
defparam \registerArray[12][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y39_N19
dffeas \registerArray[13][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][6] .is_wysiwyg = "true";
defparam \registerArray[13][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N16
cycloneive_lcell_comb \Mux57~7 (
// Equation(s):
// \Mux57~7_combout  = (cuifregT_01 & ((cuifregT_1) # ((\registerArray[13][6]~q )))) # (!cuifregT_01 & (!cuifregT_1 & (\registerArray[12][6]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[12][6]~q ),
	.datad(\registerArray[13][6]~q ),
	.cin(gnd),
	.combout(\Mux57~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~7 .lut_mask = 16'hBA98;
defparam \Mux57~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y38_N6
cycloneive_lcell_comb \Mux57~8 (
// Equation(s):
// \Mux57~8_combout  = (cuifregT_1 & ((\Mux57~7_combout  & ((\registerArray[15][6]~q ))) # (!\Mux57~7_combout  & (\registerArray[14][6]~q )))) # (!cuifregT_1 & (((\Mux57~7_combout ))))

	.dataa(\registerArray[14][6]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[15][6]~q ),
	.datad(\Mux57~7_combout ),
	.cin(gnd),
	.combout(\Mux57~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~8 .lut_mask = 16'hF388;
defparam \Mux57~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y41_N5
dffeas \registerArray[25][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][6] .is_wysiwyg = "true";
defparam \registerArray[25][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N31
dffeas \registerArray[29][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][6] .is_wysiwyg = "true";
defparam \registerArray[29][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y41_N31
dffeas \registerArray[21][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][6] .is_wysiwyg = "true";
defparam \registerArray[21][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y41_N21
dffeas \registerArray[17][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][6] .is_wysiwyg = "true";
defparam \registerArray[17][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N20
cycloneive_lcell_comb \Mux57~10 (
// Equation(s):
// \Mux57~10_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[21][6]~q )) # (!cuifregT_2 & ((\registerArray[17][6]~q )))))

	.dataa(cuifregT_3),
	.datab(\registerArray[21][6]~q ),
	.datac(\registerArray[17][6]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux57~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~10 .lut_mask = 16'hEE50;
defparam \Mux57~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N30
cycloneive_lcell_comb \Mux57~11 (
// Equation(s):
// \Mux57~11_combout  = (cuifregT_3 & ((\Mux57~10_combout  & ((\registerArray[29][6]~q ))) # (!\Mux57~10_combout  & (\registerArray[25][6]~q )))) # (!cuifregT_3 & (((\Mux57~10_combout ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[25][6]~q ),
	.datac(\registerArray[29][6]~q ),
	.datad(\Mux57~10_combout ),
	.cin(gnd),
	.combout(\Mux57~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~11 .lut_mask = 16'hF588;
defparam \Mux57~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N0
cycloneive_lcell_comb \registerArray[27][6]~feeder (
// Equation(s):
// \registerArray[27][6]~feeder_combout  = \Mux62~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux622),
	.cin(gnd),
	.combout(\registerArray[27][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[27][6]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[27][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y30_N1
dffeas \registerArray[27][6] (
	.clk(clk),
	.d(\registerArray[27][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][6] .is_wysiwyg = "true";
defparam \registerArray[27][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N15
dffeas \registerArray[31][6] (
	.clk(clk),
	.d(Mux622),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][6] .is_wysiwyg = "true";
defparam \registerArray[31][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y40_N5
dffeas \registerArray[23][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][6] .is_wysiwyg = "true";
defparam \registerArray[23][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N10
cycloneive_lcell_comb \Mux57~17 (
// Equation(s):
// \Mux57~17_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & ((\registerArray[23][6]~q ))) # (!cuifregT_2 & (\registerArray[19][6]~q ))))

	.dataa(\registerArray[19][6]~q ),
	.datab(\registerArray[23][6]~q ),
	.datac(cuifregT_3),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux57~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~17 .lut_mask = 16'hFC0A;
defparam \Mux57~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N24
cycloneive_lcell_comb \Mux57~18 (
// Equation(s):
// \Mux57~18_combout  = (cuifregT_3 & ((\Mux57~17_combout  & ((\registerArray[31][6]~q ))) # (!\Mux57~17_combout  & (\registerArray[27][6]~q )))) # (!cuifregT_3 & (((\Mux57~17_combout ))))

	.dataa(\registerArray[27][6]~q ),
	.datab(\registerArray[31][6]~q ),
	.datac(cuifregT_3),
	.datad(\Mux57~17_combout ),
	.cin(gnd),
	.combout(\Mux57~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~18 .lut_mask = 16'hCFA0;
defparam \Mux57~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y32_N1
dffeas \registerArray[22][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][6] .is_wysiwyg = "true";
defparam \registerArray[22][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N23
dffeas \registerArray[30][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][6] .is_wysiwyg = "true";
defparam \registerArray[30][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N13
dffeas \registerArray[18][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][6] .is_wysiwyg = "true";
defparam \registerArray[18][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N12
cycloneive_lcell_comb \Mux57~12 (
// Equation(s):
// \Mux57~12_combout  = (cuifregT_3 & ((\registerArray[26][6]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[18][6]~q  & !cuifregT_2))))

	.dataa(\registerArray[26][6]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[18][6]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux57~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~12 .lut_mask = 16'hCCB8;
defparam \Mux57~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N22
cycloneive_lcell_comb \Mux57~13 (
// Equation(s):
// \Mux57~13_combout  = (cuifregT_2 & ((\Mux57~12_combout  & ((\registerArray[30][6]~q ))) # (!\Mux57~12_combout  & (\registerArray[22][6]~q )))) # (!cuifregT_2 & (((\Mux57~12_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[22][6]~q ),
	.datac(\registerArray[30][6]~q ),
	.datad(\Mux57~12_combout ),
	.cin(gnd),
	.combout(\Mux57~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~13 .lut_mask = 16'hF588;
defparam \Mux57~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N23
dffeas \registerArray[28][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][6] .is_wysiwyg = "true";
defparam \registerArray[28][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N7
dffeas \registerArray[24][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][6] .is_wysiwyg = "true";
defparam \registerArray[24][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N0
cycloneive_lcell_comb \Mux57~14 (
// Equation(s):
// \Mux57~14_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & ((\registerArray[24][6]~q ))) # (!cuifregT_3 & (\registerArray[16][6]~q ))))

	.dataa(\registerArray[16][6]~q ),
	.datab(\registerArray[24][6]~q ),
	.datac(cuifregT_2),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux57~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~14 .lut_mask = 16'hFC0A;
defparam \Mux57~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N22
cycloneive_lcell_comb \Mux57~15 (
// Equation(s):
// \Mux57~15_combout  = (cuifregT_2 & ((\Mux57~14_combout  & ((\registerArray[28][6]~q ))) # (!\Mux57~14_combout  & (\registerArray[20][6]~q )))) # (!cuifregT_2 & (((\Mux57~14_combout ))))

	.dataa(\registerArray[20][6]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[28][6]~q ),
	.datad(\Mux57~14_combout ),
	.cin(gnd),
	.combout(\Mux57~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~15 .lut_mask = 16'hF388;
defparam \Mux57~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N16
cycloneive_lcell_comb \Mux57~16 (
// Equation(s):
// \Mux57~16_combout  = (cuifregT_01 & (cuifregT_1)) # (!cuifregT_01 & ((cuifregT_1 & (\Mux57~13_combout )) # (!cuifregT_1 & ((\Mux57~15_combout )))))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\Mux57~13_combout ),
	.datad(\Mux57~15_combout ),
	.cin(gnd),
	.combout(\Mux57~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~16 .lut_mask = 16'hD9C8;
defparam \Mux57~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N29
dffeas \registerArray[31][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][2] .is_wysiwyg = "true";
defparam \registerArray[31][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N25
dffeas \registerArray[19][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][2] .is_wysiwyg = "true";
defparam \registerArray[19][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N15
dffeas \registerArray[27][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][2] .is_wysiwyg = "true";
defparam \registerArray[27][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N14
cycloneive_lcell_comb \Mux29~7 (
// Equation(s):
// \Mux29~7_combout  = (cuifregS_3 & (((\registerArray[27][2]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[19][2]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[19][2]~q ),
	.datac(\registerArray[27][2]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux29~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~7 .lut_mask = 16'hAAE4;
defparam \Mux29~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N22
cycloneive_lcell_comb \Mux29~8 (
// Equation(s):
// \Mux29~8_combout  = (\Mux29~7_combout  & (((\registerArray[31][2]~q ) # (!cuifregS_2)))) # (!\Mux29~7_combout  & (\registerArray[23][2]~q  & ((cuifregS_2))))

	.dataa(\registerArray[23][2]~q ),
	.datab(\registerArray[31][2]~q ),
	.datac(\Mux29~7_combout ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux29~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~8 .lut_mask = 16'hCAF0;
defparam \Mux29~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y31_N3
dffeas \registerArray[30][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][2] .is_wysiwyg = "true";
defparam \registerArray[30][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N13
dffeas \registerArray[26][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][2] .is_wysiwyg = "true";
defparam \registerArray[26][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N7
dffeas \registerArray[22][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][2] .is_wysiwyg = "true";
defparam \registerArray[22][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N6
cycloneive_lcell_comb \Mux29~2 (
// Equation(s):
// \Mux29~2_combout  = (cuifregS_2 & (((\registerArray[22][2]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[18][2]~q  & ((!cuifregS_3))))

	.dataa(\registerArray[18][2]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[22][2]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux29~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~2 .lut_mask = 16'hCCE2;
defparam \Mux29~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N12
cycloneive_lcell_comb \Mux29~3 (
// Equation(s):
// \Mux29~3_combout  = (cuifregS_3 & ((\Mux29~2_combout  & (\registerArray[30][2]~q )) # (!\Mux29~2_combout  & ((\registerArray[26][2]~q ))))) # (!cuifregS_3 & (((\Mux29~2_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[30][2]~q ),
	.datac(\registerArray[26][2]~q ),
	.datad(\Mux29~2_combout ),
	.cin(gnd),
	.combout(\Mux29~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~3 .lut_mask = 16'hDDA0;
defparam \Mux29~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y31_N15
dffeas \registerArray[28][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][2] .is_wysiwyg = "true";
defparam \registerArray[28][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N1
dffeas \registerArray[24][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][2] .is_wysiwyg = "true";
defparam \registerArray[24][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N13
dffeas \registerArray[16][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][2] .is_wysiwyg = "true";
defparam \registerArray[16][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N19
dffeas \registerArray[20][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][2] .is_wysiwyg = "true";
defparam \registerArray[20][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N18
cycloneive_lcell_comb \Mux29~4 (
// Equation(s):
// \Mux29~4_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[20][2]~q ))) # (!cuifregS_2 & (\registerArray[16][2]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[16][2]~q ),
	.datac(\registerArray[20][2]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux29~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~4 .lut_mask = 16'hFA44;
defparam \Mux29~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N0
cycloneive_lcell_comb \Mux29~5 (
// Equation(s):
// \Mux29~5_combout  = (cuifregS_3 & ((\Mux29~4_combout  & (\registerArray[28][2]~q )) # (!\Mux29~4_combout  & ((\registerArray[24][2]~q ))))) # (!cuifregS_3 & (((\Mux29~4_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[28][2]~q ),
	.datac(\registerArray[24][2]~q ),
	.datad(\Mux29~4_combout ),
	.cin(gnd),
	.combout(\Mux29~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~5 .lut_mask = 16'hDDA0;
defparam \Mux29~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N4
cycloneive_lcell_comb \Mux29~6 (
// Equation(s):
// \Mux29~6_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\Mux29~3_combout )) # (!cuifregS_1 & ((\Mux29~5_combout )))))

	.dataa(cuifregS_0),
	.datab(\Mux29~3_combout ),
	.datac(\Mux29~5_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux29~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~6 .lut_mask = 16'hEE50;
defparam \Mux29~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N20
cycloneive_lcell_comb \registerArray[21][2]~feeder (
// Equation(s):
// \registerArray[21][2]~feeder_combout  = \Mux66~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux66),
	.cin(gnd),
	.combout(\registerArray[21][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[21][2]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[21][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N21
dffeas \registerArray[21][2] (
	.clk(clk),
	.d(\registerArray[21][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][2] .is_wysiwyg = "true";
defparam \registerArray[21][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N9
dffeas \registerArray[17][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][2] .is_wysiwyg = "true";
defparam \registerArray[17][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N24
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & (\registerArray[25][2]~q )) # (!cuifregS_3 & ((\registerArray[17][2]~q )))))

	.dataa(\registerArray[25][2]~q ),
	.datab(\registerArray[17][2]~q ),
	.datac(cuifregS_2),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'hFA0C;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N12
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// \Mux29~1_combout  = (cuifregS_2 & ((\Mux29~0_combout  & (\registerArray[29][2]~q )) # (!\Mux29~0_combout  & ((\registerArray[21][2]~q ))))) # (!cuifregS_2 & (((\Mux29~0_combout ))))

	.dataa(\registerArray[29][2]~q ),
	.datab(\registerArray[21][2]~q ),
	.datac(cuifregS_2),
	.datad(\Mux29~0_combout ),
	.cin(gnd),
	.combout(\Mux29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'hAFC0;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N26
cycloneive_lcell_comb \Mux29~9 (
// Equation(s):
// \Mux29~9_combout  = (cuifregS_0 & ((\Mux29~6_combout  & (\Mux29~8_combout )) # (!\Mux29~6_combout  & ((\Mux29~1_combout ))))) # (!cuifregS_0 & (((\Mux29~6_combout ))))

	.dataa(\Mux29~8_combout ),
	.datab(cuifregS_0),
	.datac(\Mux29~6_combout ),
	.datad(\Mux29~1_combout ),
	.cin(gnd),
	.combout(\Mux29~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~9 .lut_mask = 16'hBCB0;
defparam \Mux29~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N28
cycloneive_lcell_comb \registerArray[7][2]~feeder (
// Equation(s):
// \registerArray[7][2]~feeder_combout  = \Mux66~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux66),
	.cin(gnd),
	.combout(\registerArray[7][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[7][2]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[7][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N29
dffeas \registerArray[7][2] (
	.clk(clk),
	.d(\registerArray[7][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][2] .is_wysiwyg = "true";
defparam \registerArray[7][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N23
dffeas \registerArray[6][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][2] .is_wysiwyg = "true";
defparam \registerArray[6][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N17
dffeas \registerArray[5][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][2] .is_wysiwyg = "true";
defparam \registerArray[5][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N16
cycloneive_lcell_comb \Mux29~10 (
// Equation(s):
// \Mux29~10_combout  = (cuifregS_0 & (((\registerArray[5][2]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[4][2]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[4][2]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[5][2]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux29~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~10 .lut_mask = 16'hCCE2;
defparam \Mux29~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N22
cycloneive_lcell_comb \Mux29~11 (
// Equation(s):
// \Mux29~11_combout  = (cuifregS_1 & ((\Mux29~10_combout  & (\registerArray[7][2]~q )) # (!\Mux29~10_combout  & ((\registerArray[6][2]~q ))))) # (!cuifregS_1 & (((\Mux29~10_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[7][2]~q ),
	.datac(\registerArray[6][2]~q ),
	.datad(\Mux29~10_combout ),
	.cin(gnd),
	.combout(\Mux29~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~11 .lut_mask = 16'hDDA0;
defparam \Mux29~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N24
cycloneive_lcell_comb \registerArray[12][2]~feeder (
// Equation(s):
// \registerArray[12][2]~feeder_combout  = \Mux66~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux66),
	.cin(gnd),
	.combout(\registerArray[12][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[12][2]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[12][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N25
dffeas \registerArray[12][2] (
	.clk(clk),
	.d(\registerArray[12][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][2] .is_wysiwyg = "true";
defparam \registerArray[12][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N9
dffeas \registerArray[13][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][2] .is_wysiwyg = "true";
defparam \registerArray[13][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N8
cycloneive_lcell_comb \Mux29~17 (
// Equation(s):
// \Mux29~17_combout  = (cuifregS_0 & (((\registerArray[13][2]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[12][2]~q  & ((!cuifregS_1))))

	.dataa(cuifregS_0),
	.datab(\registerArray[12][2]~q ),
	.datac(\registerArray[13][2]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux29~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~17 .lut_mask = 16'hAAE4;
defparam \Mux29~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N27
dffeas \registerArray[14][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][2] .is_wysiwyg = "true";
defparam \registerArray[14][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N26
cycloneive_lcell_comb \Mux29~18 (
// Equation(s):
// \Mux29~18_combout  = (\Mux29~17_combout  & ((\registerArray[15][2]~q ) # ((!cuifregS_1)))) # (!\Mux29~17_combout  & (((\registerArray[14][2]~q  & cuifregS_1))))

	.dataa(\registerArray[15][2]~q ),
	.datab(\Mux29~17_combout ),
	.datac(\registerArray[14][2]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux29~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~18 .lut_mask = 16'hB8CC;
defparam \Mux29~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N21
dffeas \registerArray[2][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][2] .is_wysiwyg = "true";
defparam \registerArray[2][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N26
cycloneive_lcell_comb \registerArray[1][2]~feeder (
// Equation(s):
// \registerArray[1][2]~feeder_combout  = \Mux66~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux66),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[1][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[1][2]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[1][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y42_N27
dffeas \registerArray[1][2] (
	.clk(clk),
	.d(\registerArray[1][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][2] .is_wysiwyg = "true";
defparam \registerArray[1][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N6
cycloneive_lcell_comb \Mux29~14 (
// Equation(s):
// \Mux29~14_combout  = (cuifregS_0 & ((cuifregS_1 & (\registerArray[3][2]~q )) # (!cuifregS_1 & ((\registerArray[1][2]~q )))))

	.dataa(\registerArray[3][2]~q ),
	.datab(\registerArray[1][2]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux29~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~14 .lut_mask = 16'hA0C0;
defparam \Mux29~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N20
cycloneive_lcell_comb \Mux29~15 (
// Equation(s):
// \Mux29~15_combout  = (\Mux29~14_combout ) # ((cuifregS_1 & (!cuifregS_0 & \registerArray[2][2]~q )))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\registerArray[2][2]~q ),
	.datad(\Mux29~14_combout ),
	.cin(gnd),
	.combout(\Mux29~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~15 .lut_mask = 16'hFF20;
defparam \Mux29~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N9
dffeas \registerArray[9][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][2] .is_wysiwyg = "true";
defparam \registerArray[9][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N27
dffeas \registerArray[11][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][2] .is_wysiwyg = "true";
defparam \registerArray[11][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N7
dffeas \registerArray[8][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][2] .is_wysiwyg = "true";
defparam \registerArray[8][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N6
cycloneive_lcell_comb \Mux29~12 (
// Equation(s):
// \Mux29~12_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\registerArray[10][2]~q )) # (!cuifregS_1 & ((\registerArray[8][2]~q )))))

	.dataa(\registerArray[10][2]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[8][2]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux29~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~12 .lut_mask = 16'hEE30;
defparam \Mux29~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N26
cycloneive_lcell_comb \Mux29~13 (
// Equation(s):
// \Mux29~13_combout  = (cuifregS_0 & ((\Mux29~12_combout  & ((\registerArray[11][2]~q ))) # (!\Mux29~12_combout  & (\registerArray[9][2]~q )))) # (!cuifregS_0 & (((\Mux29~12_combout ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[9][2]~q ),
	.datac(\registerArray[11][2]~q ),
	.datad(\Mux29~12_combout ),
	.cin(gnd),
	.combout(\Mux29~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~13 .lut_mask = 16'hF588;
defparam \Mux29~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N18
cycloneive_lcell_comb \Mux29~16 (
// Equation(s):
// \Mux29~16_combout  = (cuifregS_3 & ((cuifregS_2) # ((\Mux29~13_combout )))) # (!cuifregS_3 & (!cuifregS_2 & (\Mux29~15_combout )))

	.dataa(cuifregS_3),
	.datab(cuifregS_2),
	.datac(\Mux29~15_combout ),
	.datad(\Mux29~13_combout ),
	.cin(gnd),
	.combout(\Mux29~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~16 .lut_mask = 16'hBA98;
defparam \Mux29~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N16
cycloneive_lcell_comb \Mux29~19 (
// Equation(s):
// \Mux29~19_combout  = (cuifregS_2 & ((\Mux29~16_combout  & ((\Mux29~18_combout ))) # (!\Mux29~16_combout  & (\Mux29~11_combout )))) # (!cuifregS_2 & (((\Mux29~16_combout ))))

	.dataa(\Mux29~11_combout ),
	.datab(cuifregS_2),
	.datac(\Mux29~18_combout ),
	.datad(\Mux29~16_combout ),
	.cin(gnd),
	.combout(\Mux29~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~19 .lut_mask = 16'hF388;
defparam \Mux29~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N19
dffeas \registerArray[25][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][1] .is_wysiwyg = "true";
defparam \registerArray[25][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N0
cycloneive_lcell_comb \registerArray[21][1]~feeder (
// Equation(s):
// \registerArray[21][1]~feeder_combout  = \Mux67~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux67),
	.cin(gnd),
	.combout(\registerArray[21][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[21][1]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[21][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N1
dffeas \registerArray[21][1] (
	.clk(clk),
	.d(\registerArray[21][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][1] .is_wysiwyg = "true";
defparam \registerArray[21][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N10
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// \Mux30~0_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[21][1]~q ))) # (!cuifregS_2 & (\registerArray[17][1]~q ))))

	.dataa(\registerArray[17][1]~q ),
	.datab(cuifregS_3),
	.datac(cuifregS_2),
	.datad(\registerArray[21][1]~q ),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'hF2C2;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N18
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// \Mux30~1_combout  = (cuifregS_3 & ((\Mux30~0_combout  & (\registerArray[29][1]~q )) # (!\Mux30~0_combout  & ((\registerArray[25][1]~q ))))) # (!cuifregS_3 & (((\Mux30~0_combout ))))

	.dataa(\registerArray[29][1]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[25][1]~q ),
	.datad(\Mux30~0_combout ),
	.cin(gnd),
	.combout(\Mux30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'hBBC0;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y31_N19
dffeas \registerArray[30][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][1] .is_wysiwyg = "true";
defparam \registerArray[30][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N21
dffeas \registerArray[22][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][1] .is_wysiwyg = "true";
defparam \registerArray[22][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N4
cycloneive_lcell_comb \registerArray[18][1]~feeder (
// Equation(s):
// \registerArray[18][1]~feeder_combout  = \Mux67~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux67),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[18][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[18][1]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[18][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y31_N5
dffeas \registerArray[18][1] (
	.clk(clk),
	.d(\registerArray[18][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][1] .is_wysiwyg = "true";
defparam \registerArray[18][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N3
dffeas \registerArray[26][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][1] .is_wysiwyg = "true";
defparam \registerArray[26][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N2
cycloneive_lcell_comb \Mux30~2 (
// Equation(s):
// \Mux30~2_combout  = (cuifregS_3 & (((\registerArray[26][1]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[18][1]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[18][1]~q ),
	.datac(\registerArray[26][1]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~2 .lut_mask = 16'hAAE4;
defparam \Mux30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N20
cycloneive_lcell_comb \Mux30~3 (
// Equation(s):
// \Mux30~3_combout  = (cuifregS_2 & ((\Mux30~2_combout  & (\registerArray[30][1]~q )) # (!\Mux30~2_combout  & ((\registerArray[22][1]~q ))))) # (!cuifregS_2 & (((\Mux30~2_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[30][1]~q ),
	.datac(\registerArray[22][1]~q ),
	.datad(\Mux30~2_combout ),
	.cin(gnd),
	.combout(\Mux30~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~3 .lut_mask = 16'hDDA0;
defparam \Mux30~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y32_N27
dffeas \registerArray[28][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][1] .is_wysiwyg = "true";
defparam \registerArray[28][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N5
dffeas \registerArray[20][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][1] .is_wysiwyg = "true";
defparam \registerArray[20][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N1
dffeas \registerArray[16][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][1] .is_wysiwyg = "true";
defparam \registerArray[16][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N3
dffeas \registerArray[24][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][1] .is_wysiwyg = "true";
defparam \registerArray[24][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N2
cycloneive_lcell_comb \Mux30~4 (
// Equation(s):
// \Mux30~4_combout  = (cuifregS_3 & (((\registerArray[24][1]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[16][1]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[16][1]~q ),
	.datac(\registerArray[24][1]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux30~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~4 .lut_mask = 16'hAAE4;
defparam \Mux30~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N4
cycloneive_lcell_comb \Mux30~5 (
// Equation(s):
// \Mux30~5_combout  = (cuifregS_2 & ((\Mux30~4_combout  & (\registerArray[28][1]~q )) # (!\Mux30~4_combout  & ((\registerArray[20][1]~q ))))) # (!cuifregS_2 & (((\Mux30~4_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[28][1]~q ),
	.datac(\registerArray[20][1]~q ),
	.datad(\Mux30~4_combout ),
	.cin(gnd),
	.combout(\Mux30~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~5 .lut_mask = 16'hDDA0;
defparam \Mux30~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N8
cycloneive_lcell_comb \Mux30~6 (
// Equation(s):
// \Mux30~6_combout  = (cuifregS_1 & ((cuifregS_0) # ((\Mux30~3_combout )))) # (!cuifregS_1 & (!cuifregS_0 & ((\Mux30~5_combout ))))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\Mux30~3_combout ),
	.datad(\Mux30~5_combout ),
	.cin(gnd),
	.combout(\Mux30~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~6 .lut_mask = 16'hB9A8;
defparam \Mux30~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y30_N5
dffeas \registerArray[31][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][1] .is_wysiwyg = "true";
defparam \registerArray[31][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N24
cycloneive_lcell_comb \registerArray[27][1]~feeder (
// Equation(s):
// \registerArray[27][1]~feeder_combout  = \Mux67~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux67),
	.cin(gnd),
	.combout(\registerArray[27][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[27][1]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[27][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y37_N25
dffeas \registerArray[27][1] (
	.clk(clk),
	.d(\registerArray[27][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][1] .is_wysiwyg = "true";
defparam \registerArray[27][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N6
cycloneive_lcell_comb \Mux30~8 (
// Equation(s):
// \Mux30~8_combout  = (\Mux30~7_combout  & (((\registerArray[31][1]~q )) # (!cuifregS_3))) # (!\Mux30~7_combout  & (cuifregS_3 & ((\registerArray[27][1]~q ))))

	.dataa(\Mux30~7_combout ),
	.datab(cuifregS_3),
	.datac(\registerArray[31][1]~q ),
	.datad(\registerArray[27][1]~q ),
	.cin(gnd),
	.combout(\Mux30~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~8 .lut_mask = 16'hE6A2;
defparam \Mux30~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N28
cycloneive_lcell_comb \Mux30~9 (
// Equation(s):
// \Mux30~9_combout  = (cuifregS_0 & ((\Mux30~6_combout  & ((\Mux30~8_combout ))) # (!\Mux30~6_combout  & (\Mux30~1_combout )))) # (!cuifregS_0 & (((\Mux30~6_combout ))))

	.dataa(\Mux30~1_combout ),
	.datab(cuifregS_0),
	.datac(\Mux30~6_combout ),
	.datad(\Mux30~8_combout ),
	.cin(gnd),
	.combout(\Mux30~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~9 .lut_mask = 16'hF838;
defparam \Mux30~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N17
dffeas \registerArray[9][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][1] .is_wysiwyg = "true";
defparam \registerArray[9][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N23
dffeas \registerArray[11][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][1] .is_wysiwyg = "true";
defparam \registerArray[11][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N16
cycloneive_lcell_comb \Mux30~11 (
// Equation(s):
// \Mux30~11_combout  = (\Mux30~10_combout  & (((\registerArray[11][1]~q )) # (!cuifregS_0))) # (!\Mux30~10_combout  & (cuifregS_0 & (\registerArray[9][1]~q )))

	.dataa(\Mux30~10_combout ),
	.datab(cuifregS_0),
	.datac(\registerArray[9][1]~q ),
	.datad(\registerArray[11][1]~q ),
	.cin(gnd),
	.combout(\Mux30~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~11 .lut_mask = 16'hEA62;
defparam \Mux30~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N4
cycloneive_lcell_comb \registerArray[14][1]~feeder (
// Equation(s):
// \registerArray[14][1]~feeder_combout  = \Mux67~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux67),
	.cin(gnd),
	.combout(\registerArray[14][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][1]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[14][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N5
dffeas \registerArray[14][1] (
	.clk(clk),
	.d(\registerArray[14][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][1] .is_wysiwyg = "true";
defparam \registerArray[14][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N31
dffeas \registerArray[15][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][1] .is_wysiwyg = "true";
defparam \registerArray[15][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N22
cycloneive_lcell_comb \registerArray[13][1]~feeder (
// Equation(s):
// \registerArray[13][1]~feeder_combout  = \Mux67~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux67),
	.cin(gnd),
	.combout(\registerArray[13][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[13][1]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[13][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N23
dffeas \registerArray[13][1] (
	.clk(clk),
	.d(\registerArray[13][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][1] .is_wysiwyg = "true";
defparam \registerArray[13][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N4
cycloneive_lcell_comb \registerArray[12][1]~feeder (
// Equation(s):
// \registerArray[12][1]~feeder_combout  = \Mux67~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux67),
	.cin(gnd),
	.combout(\registerArray[12][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[12][1]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[12][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N5
dffeas \registerArray[12][1] (
	.clk(clk),
	.d(\registerArray[12][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][1] .is_wysiwyg = "true";
defparam \registerArray[12][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N12
cycloneive_lcell_comb \Mux30~17 (
// Equation(s):
// \Mux30~17_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & (\registerArray[13][1]~q )) # (!cuifregS_0 & ((\registerArray[12][1]~q )))))

	.dataa(cuifregS_1),
	.datab(\registerArray[13][1]~q ),
	.datac(\registerArray[12][1]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux30~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~17 .lut_mask = 16'hEE50;
defparam \Mux30~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N6
cycloneive_lcell_comb \Mux30~18 (
// Equation(s):
// \Mux30~18_combout  = (cuifregS_1 & ((\Mux30~17_combout  & ((\registerArray[15][1]~q ))) # (!\Mux30~17_combout  & (\registerArray[14][1]~q )))) # (!cuifregS_1 & (((\Mux30~17_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[14][1]~q ),
	.datac(\registerArray[15][1]~q ),
	.datad(\Mux30~17_combout ),
	.cin(gnd),
	.combout(\Mux30~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~18 .lut_mask = 16'hF588;
defparam \Mux30~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N11
dffeas \registerArray[1][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][1] .is_wysiwyg = "true";
defparam \registerArray[1][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N14
cycloneive_lcell_comb \registerArray[3][1]~feeder (
// Equation(s):
// \registerArray[3][1]~feeder_combout  = \Mux67~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux67),
	.cin(gnd),
	.combout(\registerArray[3][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[3][1]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[3][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y37_N15
dffeas \registerArray[3][1] (
	.clk(clk),
	.d(\registerArray[3][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][1] .is_wysiwyg = "true";
defparam \registerArray[3][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N4
cycloneive_lcell_comb \Mux30~14 (
// Equation(s):
// \Mux30~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][1]~q ))) # (!cuifregS_1 & (\registerArray[1][1]~q ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[1][1]~q ),
	.datac(\registerArray[3][1]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux30~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~14 .lut_mask = 16'hE400;
defparam \Mux30~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N30
cycloneive_lcell_comb \Mux30~15 (
// Equation(s):
// \Mux30~15_combout  = (\Mux30~14_combout ) # ((\registerArray[2][1]~q  & (cuifregS_1 & !cuifregS_0)))

	.dataa(\registerArray[2][1]~q ),
	.datab(\Mux30~14_combout ),
	.datac(cuifregS_1),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux30~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~15 .lut_mask = 16'hCCEC;
defparam \Mux30~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N18
cycloneive_lcell_comb \registerArray[6][1]~feeder (
// Equation(s):
// \registerArray[6][1]~feeder_combout  = \Mux67~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux67),
	.cin(gnd),
	.combout(\registerArray[6][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[6][1]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[6][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N19
dffeas \registerArray[6][1] (
	.clk(clk),
	.d(\registerArray[6][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][1] .is_wysiwyg = "true";
defparam \registerArray[6][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N29
dffeas \registerArray[7][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][1] .is_wysiwyg = "true";
defparam \registerArray[7][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N29
dffeas \registerArray[5][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][1] .is_wysiwyg = "true";
defparam \registerArray[5][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N28
cycloneive_lcell_comb \Mux30~12 (
// Equation(s):
// \Mux30~12_combout  = (cuifregS_0 & (((\registerArray[5][1]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[4][1]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[4][1]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[5][1]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux30~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~12 .lut_mask = 16'hCCE2;
defparam \Mux30~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N26
cycloneive_lcell_comb \Mux30~13 (
// Equation(s):
// \Mux30~13_combout  = (cuifregS_1 & ((\Mux30~12_combout  & ((\registerArray[7][1]~q ))) # (!\Mux30~12_combout  & (\registerArray[6][1]~q )))) # (!cuifregS_1 & (((\Mux30~12_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[6][1]~q ),
	.datac(\registerArray[7][1]~q ),
	.datad(\Mux30~12_combout ),
	.cin(gnd),
	.combout(\Mux30~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~13 .lut_mask = 16'hF588;
defparam \Mux30~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N16
cycloneive_lcell_comb \Mux30~16 (
// Equation(s):
// \Mux30~16_combout  = (cuifregS_2 & ((cuifregS_3) # ((\Mux30~13_combout )))) # (!cuifregS_2 & (!cuifregS_3 & (\Mux30~15_combout )))

	.dataa(cuifregS_2),
	.datab(cuifregS_3),
	.datac(\Mux30~15_combout ),
	.datad(\Mux30~13_combout ),
	.cin(gnd),
	.combout(\Mux30~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~16 .lut_mask = 16'hBA98;
defparam \Mux30~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N18
cycloneive_lcell_comb \Mux30~19 (
// Equation(s):
// \Mux30~19_combout  = (cuifregS_3 & ((\Mux30~16_combout  & ((\Mux30~18_combout ))) # (!\Mux30~16_combout  & (\Mux30~11_combout )))) # (!cuifregS_3 & (((\Mux30~16_combout ))))

	.dataa(\Mux30~11_combout ),
	.datab(cuifregS_3),
	.datac(\Mux30~18_combout ),
	.datad(\Mux30~16_combout ),
	.cin(gnd),
	.combout(\Mux30~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~19 .lut_mask = 16'hF388;
defparam \Mux30~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N20
cycloneive_lcell_comb \Mux62~7 (
// Equation(s):
// \Mux62~7_combout  = (cuifregT_01 & (((\registerArray[13][1]~q ) # (cuifregT_1)))) # (!cuifregT_01 & (\registerArray[12][1]~q  & ((!cuifregT_1))))

	.dataa(\registerArray[12][1]~q ),
	.datab(\registerArray[13][1]~q ),
	.datac(cuifregT_0),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux62~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~7 .lut_mask = 16'hF0CA;
defparam \Mux62~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N30
cycloneive_lcell_comb \Mux62~8 (
// Equation(s):
// \Mux62~8_combout  = (cuifregT_1 & ((\Mux62~7_combout  & ((\registerArray[15][1]~q ))) # (!\Mux62~7_combout  & (\registerArray[14][1]~q )))) # (!cuifregT_1 & (((\Mux62~7_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[14][1]~q ),
	.datac(\registerArray[15][1]~q ),
	.datad(\Mux62~7_combout ),
	.cin(gnd),
	.combout(\Mux62~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~8 .lut_mask = 16'hF588;
defparam \Mux62~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N7
dffeas \registerArray[4][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][1] .is_wysiwyg = "true";
defparam \registerArray[4][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N6
cycloneive_lcell_comb \Mux62~0 (
// Equation(s):
// \Mux62~0_combout  = (cuifregT_01 & ((\registerArray[5][1]~q ) # ((cuifregT_1)))) # (!cuifregT_01 & (((\registerArray[4][1]~q  & !cuifregT_1))))

	.dataa(cuifregT_0),
	.datab(\registerArray[5][1]~q ),
	.datac(\registerArray[4][1]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux62~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~0 .lut_mask = 16'hAAD8;
defparam \Mux62~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N28
cycloneive_lcell_comb \Mux62~1 (
// Equation(s):
// \Mux62~1_combout  = (cuifregT_1 & ((\Mux62~0_combout  & ((\registerArray[7][1]~q ))) # (!\Mux62~0_combout  & (\registerArray[6][1]~q )))) # (!cuifregT_1 & (((\Mux62~0_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[6][1]~q ),
	.datac(\registerArray[7][1]~q ),
	.datad(\Mux62~0_combout ),
	.cin(gnd),
	.combout(\Mux62~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~1 .lut_mask = 16'hF588;
defparam \Mux62~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y31_N25
dffeas \registerArray[8][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][1] .is_wysiwyg = "true";
defparam \registerArray[8][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N24
cycloneive_lcell_comb \Mux62~2 (
// Equation(s):
// \Mux62~2_combout  = (cuifregT_1 & ((\registerArray[10][1]~q ) # ((cuifregT_01)))) # (!cuifregT_1 & (((\registerArray[8][1]~q  & !cuifregT_01))))

	.dataa(\registerArray[10][1]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[8][1]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux62~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~2 .lut_mask = 16'hCCB8;
defparam \Mux62~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N22
cycloneive_lcell_comb \Mux62~3 (
// Equation(s):
// \Mux62~3_combout  = (cuifregT_01 & ((\Mux62~2_combout  & ((\registerArray[11][1]~q ))) # (!\Mux62~2_combout  & (\registerArray[9][1]~q )))) # (!cuifregT_01 & (((\Mux62~2_combout ))))

	.dataa(\registerArray[9][1]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[11][1]~q ),
	.datad(\Mux62~2_combout ),
	.cin(gnd),
	.combout(\Mux62~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~3 .lut_mask = 16'hF388;
defparam \Mux62~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y37_N13
dffeas \registerArray[2][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][1] .is_wysiwyg = "true";
defparam \registerArray[2][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N10
cycloneive_lcell_comb \Mux62~4 (
// Equation(s):
// \Mux62~4_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][1]~q )) # (!cuifregT_1 & ((\registerArray[1][1]~q )))))

	.dataa(\registerArray[3][1]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[1][1]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux62~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~4 .lut_mask = 16'h88C0;
defparam \Mux62~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N12
cycloneive_lcell_comb \Mux62~5 (
// Equation(s):
// \Mux62~5_combout  = (\Mux62~4_combout ) # ((cuifregT_1 & (!cuifregT_01 & \registerArray[2][1]~q )))

	.dataa(cuifregT_1),
	.datab(cuifregT_0),
	.datac(\registerArray[2][1]~q ),
	.datad(\Mux62~4_combout ),
	.cin(gnd),
	.combout(\Mux62~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~5 .lut_mask = 16'hFF20;
defparam \Mux62~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N2
cycloneive_lcell_comb \Mux62~6 (
// Equation(s):
// \Mux62~6_combout  = (cuifregT_2 & (cuifregT_3)) # (!cuifregT_2 & ((cuifregT_3 & (\Mux62~3_combout )) # (!cuifregT_3 & ((\Mux62~5_combout )))))

	.dataa(cuifregT_2),
	.datab(cuifregT_3),
	.datac(\Mux62~3_combout ),
	.datad(\Mux62~5_combout ),
	.cin(gnd),
	.combout(\Mux62~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~6 .lut_mask = 16'hD9C8;
defparam \Mux62~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N9
dffeas \registerArray[23][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][1] .is_wysiwyg = "true";
defparam \registerArray[23][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N7
dffeas \registerArray[19][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][1] .is_wysiwyg = "true";
defparam \registerArray[19][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N6
cycloneive_lcell_comb \Mux62~17 (
// Equation(s):
// \Mux62~17_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[27][1]~q )) # (!cuifregT_3 & ((\registerArray[19][1]~q )))))

	.dataa(cuifregT_2),
	.datab(\registerArray[27][1]~q ),
	.datac(\registerArray[19][1]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux62~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~17 .lut_mask = 16'hEE50;
defparam \Mux62~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N4
cycloneive_lcell_comb \Mux62~18 (
// Equation(s):
// \Mux62~18_combout  = (cuifregT_2 & ((\Mux62~17_combout  & ((\registerArray[31][1]~q ))) # (!\Mux62~17_combout  & (\registerArray[23][1]~q )))) # (!cuifregT_2 & (((\Mux62~17_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[23][1]~q ),
	.datac(\registerArray[31][1]~q ),
	.datad(\Mux62~17_combout ),
	.cin(gnd),
	.combout(\Mux62~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~18 .lut_mask = 16'hF588;
defparam \Mux62~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N0
cycloneive_lcell_comb \Mux62~14 (
// Equation(s):
// \Mux62~14_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[20][1]~q )) # (!cuifregT_2 & ((\registerArray[16][1]~q )))))

	.dataa(\registerArray[20][1]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[16][1]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux62~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~14 .lut_mask = 16'hEE30;
defparam \Mux62~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N26
cycloneive_lcell_comb \Mux62~15 (
// Equation(s):
// \Mux62~15_combout  = (cuifregT_3 & ((\Mux62~14_combout  & ((\registerArray[28][1]~q ))) # (!\Mux62~14_combout  & (\registerArray[24][1]~q )))) # (!cuifregT_3 & (((\Mux62~14_combout ))))

	.dataa(\registerArray[24][1]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[28][1]~q ),
	.datad(\Mux62~14_combout ),
	.cin(gnd),
	.combout(\Mux62~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~15 .lut_mask = 16'hF388;
defparam \Mux62~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N0
cycloneive_lcell_comb \Mux62~12 (
// Equation(s):
// \Mux62~12_combout  = (cuifregT_2 & (((\registerArray[22][1]~q ) # (cuifregT_3)))) # (!cuifregT_2 & (\registerArray[18][1]~q  & ((!cuifregT_3))))

	.dataa(\registerArray[18][1]~q ),
	.datab(\registerArray[22][1]~q ),
	.datac(cuifregT_2),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux62~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~12 .lut_mask = 16'hF0CA;
defparam \Mux62~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N18
cycloneive_lcell_comb \Mux62~13 (
// Equation(s):
// \Mux62~13_combout  = (cuifregT_3 & ((\Mux62~12_combout  & ((\registerArray[30][1]~q ))) # (!\Mux62~12_combout  & (\registerArray[26][1]~q )))) # (!cuifregT_3 & (((\Mux62~12_combout ))))

	.dataa(\registerArray[26][1]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[30][1]~q ),
	.datad(\Mux62~12_combout ),
	.cin(gnd),
	.combout(\Mux62~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~13 .lut_mask = 16'hF388;
defparam \Mux62~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N4
cycloneive_lcell_comb \Mux62~16 (
// Equation(s):
// \Mux62~16_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & ((\Mux62~13_combout ))) # (!cuifregT_1 & (\Mux62~15_combout ))))

	.dataa(\Mux62~15_combout ),
	.datab(cuifregT_0),
	.datac(cuifregT_1),
	.datad(\Mux62~13_combout ),
	.cin(gnd),
	.combout(\Mux62~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~16 .lut_mask = 16'hF2C2;
defparam \Mux62~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N4
cycloneive_lcell_comb \registerArray[29][1]~feeder (
// Equation(s):
// \registerArray[29][1]~feeder_combout  = \Mux67~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux67),
	.cin(gnd),
	.combout(\registerArray[29][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[29][1]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[29][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N5
dffeas \registerArray[29][1] (
	.clk(clk),
	.d(\registerArray[29][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][1] .is_wysiwyg = "true";
defparam \registerArray[29][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y31_N9
dffeas \registerArray[17][1] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux67),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][1] .is_wysiwyg = "true";
defparam \registerArray[17][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N8
cycloneive_lcell_comb \Mux62~10 (
// Equation(s):
// \Mux62~10_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[25][1]~q )) # (!cuifregT_3 & ((\registerArray[17][1]~q )))))

	.dataa(cuifregT_2),
	.datab(\registerArray[25][1]~q ),
	.datac(\registerArray[17][1]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux62~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~10 .lut_mask = 16'hEE50;
defparam \Mux62~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N14
cycloneive_lcell_comb \Mux62~11 (
// Equation(s):
// \Mux62~11_combout  = (cuifregT_2 & ((\Mux62~10_combout  & ((\registerArray[29][1]~q ))) # (!\Mux62~10_combout  & (\registerArray[21][1]~q )))) # (!cuifregT_2 & (((\Mux62~10_combout ))))

	.dataa(\registerArray[21][1]~q ),
	.datab(\registerArray[29][1]~q ),
	.datac(cuifregT_2),
	.datad(\Mux62~10_combout ),
	.cin(gnd),
	.combout(\Mux62~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~11 .lut_mask = 16'hCFA0;
defparam \Mux62~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y39_N1
dffeas \registerArray[7][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][4] .is_wysiwyg = "true";
defparam \registerArray[7][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y39_N11
dffeas \registerArray[6][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][4] .is_wysiwyg = "true";
defparam \registerArray[6][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N9
dffeas \registerArray[5][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][4] .is_wysiwyg = "true";
defparam \registerArray[5][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N8
cycloneive_lcell_comb \Mux27~10 (
// Equation(s):
// \Mux27~10_combout  = (cuifregS_0 & (((\registerArray[5][4]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[4][4]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[4][4]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[5][4]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux27~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~10 .lut_mask = 16'hCCE2;
defparam \Mux27~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N10
cycloneive_lcell_comb \Mux27~11 (
// Equation(s):
// \Mux27~11_combout  = (cuifregS_1 & ((\Mux27~10_combout  & (\registerArray[7][4]~q )) # (!\Mux27~10_combout  & ((\registerArray[6][4]~q ))))) # (!cuifregS_1 & (((\Mux27~10_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[7][4]~q ),
	.datac(\registerArray[6][4]~q ),
	.datad(\Mux27~10_combout ),
	.cin(gnd),
	.combout(\Mux27~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~11 .lut_mask = 16'hDDA0;
defparam \Mux27~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N25
dffeas \registerArray[9][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][4] .is_wysiwyg = "true";
defparam \registerArray[9][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N3
dffeas \registerArray[11][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][4] .is_wysiwyg = "true";
defparam \registerArray[11][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y35_N11
dffeas \registerArray[8][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][4] .is_wysiwyg = "true";
defparam \registerArray[8][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N10
cycloneive_lcell_comb \Mux27~12 (
// Equation(s):
// \Mux27~12_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\registerArray[10][4]~q )) # (!cuifregS_1 & ((\registerArray[8][4]~q )))))

	.dataa(\registerArray[10][4]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[8][4]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux27~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~12 .lut_mask = 16'hEE30;
defparam \Mux27~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N2
cycloneive_lcell_comb \Mux27~13 (
// Equation(s):
// \Mux27~13_combout  = (cuifregS_0 & ((\Mux27~12_combout  & ((\registerArray[11][4]~q ))) # (!\Mux27~12_combout  & (\registerArray[9][4]~q )))) # (!cuifregS_0 & (((\Mux27~12_combout ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[9][4]~q ),
	.datac(\registerArray[11][4]~q ),
	.datad(\Mux27~12_combout ),
	.cin(gnd),
	.combout(\Mux27~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~13 .lut_mask = 16'hF588;
defparam \Mux27~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N7
dffeas \registerArray[2][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][4] .is_wysiwyg = "true";
defparam \registerArray[2][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N2
cycloneive_lcell_comb \registerArray[3][4]~feeder (
// Equation(s):
// \registerArray[3][4]~feeder_combout  = \Mux64~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux64),
	.cin(gnd),
	.combout(\registerArray[3][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[3][4]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[3][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y42_N3
dffeas \registerArray[3][4] (
	.clk(clk),
	.d(\registerArray[3][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][4] .is_wysiwyg = "true";
defparam \registerArray[3][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N10
cycloneive_lcell_comb \Mux27~14 (
// Equation(s):
// \Mux27~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][4]~q ))) # (!cuifregS_1 & (\registerArray[1][4]~q ))))

	.dataa(\registerArray[1][4]~q ),
	.datab(\registerArray[3][4]~q ),
	.datac(cuifregS_1),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux27~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~14 .lut_mask = 16'hCA00;
defparam \Mux27~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N6
cycloneive_lcell_comb \Mux27~15 (
// Equation(s):
// \Mux27~15_combout  = (\Mux27~14_combout ) # ((cuifregS_1 & (!cuifregS_0 & \registerArray[2][4]~q )))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\registerArray[2][4]~q ),
	.datad(\Mux27~14_combout ),
	.cin(gnd),
	.combout(\Mux27~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~15 .lut_mask = 16'hFF20;
defparam \Mux27~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N14
cycloneive_lcell_comb \Mux27~16 (
// Equation(s):
// \Mux27~16_combout  = (cuifregS_3 & ((cuifregS_2) # ((\Mux27~13_combout )))) # (!cuifregS_3 & (!cuifregS_2 & ((\Mux27~15_combout ))))

	.dataa(cuifregS_3),
	.datab(cuifregS_2),
	.datac(\Mux27~13_combout ),
	.datad(\Mux27~15_combout ),
	.cin(gnd),
	.combout(\Mux27~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~16 .lut_mask = 16'hB9A8;
defparam \Mux27~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N6
cycloneive_lcell_comb \registerArray[15][4]~feeder (
// Equation(s):
// \registerArray[15][4]~feeder_combout  = \Mux64~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux64),
	.cin(gnd),
	.combout(\registerArray[15][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[15][4]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[15][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y32_N7
dffeas \registerArray[15][4] (
	.clk(clk),
	.d(\registerArray[15][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][4] .is_wysiwyg = "true";
defparam \registerArray[15][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N23
dffeas \registerArray[13][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][4] .is_wysiwyg = "true";
defparam \registerArray[13][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N0
cycloneive_lcell_comb \Mux27~17 (
// Equation(s):
// \Mux27~17_combout  = (cuifregS_0 & (((\registerArray[13][4]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[12][4]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[12][4]~q ),
	.datab(\registerArray[13][4]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux27~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~17 .lut_mask = 16'hF0CA;
defparam \Mux27~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N8
cycloneive_lcell_comb \Mux27~18 (
// Equation(s):
// \Mux27~18_combout  = (\Mux27~17_combout  & (((\registerArray[15][4]~q ) # (!cuifregS_1)))) # (!\Mux27~17_combout  & (\registerArray[14][4]~q  & ((cuifregS_1))))

	.dataa(\registerArray[14][4]~q ),
	.datab(\registerArray[15][4]~q ),
	.datac(\Mux27~17_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux27~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~18 .lut_mask = 16'hCAF0;
defparam \Mux27~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N4
cycloneive_lcell_comb \Mux27~19 (
// Equation(s):
// \Mux27~19_combout  = (cuifregS_2 & ((\Mux27~16_combout  & ((\Mux27~18_combout ))) # (!\Mux27~16_combout  & (\Mux27~11_combout )))) # (!cuifregS_2 & (((\Mux27~16_combout ))))

	.dataa(\Mux27~11_combout ),
	.datab(cuifregS_2),
	.datac(\Mux27~16_combout ),
	.datad(\Mux27~18_combout ),
	.cin(gnd),
	.combout(\Mux27~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~19 .lut_mask = 16'hF838;
defparam \Mux27~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N24
cycloneive_lcell_comb \registerArray[21][4]~feeder (
// Equation(s):
// \registerArray[21][4]~feeder_combout  = \Mux64~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux64),
	.cin(gnd),
	.combout(\registerArray[21][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[21][4]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[21][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N25
dffeas \registerArray[21][4] (
	.clk(clk),
	.d(\registerArray[21][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][4] .is_wysiwyg = "true";
defparam \registerArray[21][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N23
dffeas \registerArray[17][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][4] .is_wysiwyg = "true";
defparam \registerArray[17][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N0
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (cuifregS_3 & ((\registerArray[25][4]~q ) # ((cuifregS_2)))) # (!cuifregS_3 & (((\registerArray[17][4]~q  & !cuifregS_2))))

	.dataa(\registerArray[25][4]~q ),
	.datab(\registerArray[17][4]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'hF0AC;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N18
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// \Mux27~1_combout  = (cuifregS_2 & ((\Mux27~0_combout  & (\registerArray[29][4]~q )) # (!\Mux27~0_combout  & ((\registerArray[21][4]~q ))))) # (!cuifregS_2 & (((\Mux27~0_combout ))))

	.dataa(\registerArray[29][4]~q ),
	.datab(\registerArray[21][4]~q ),
	.datac(cuifregS_2),
	.datad(\Mux27~0_combout ),
	.cin(gnd),
	.combout(\Mux27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hAFC0;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y31_N21
dffeas \registerArray[30][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][4] .is_wysiwyg = "true";
defparam \registerArray[30][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N17
dffeas \registerArray[26][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][4] .is_wysiwyg = "true";
defparam \registerArray[26][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N11
dffeas \registerArray[18][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][4] .is_wysiwyg = "true";
defparam \registerArray[18][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N11
dffeas \registerArray[22][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][4] .is_wysiwyg = "true";
defparam \registerArray[22][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N10
cycloneive_lcell_comb \Mux27~2 (
// Equation(s):
// \Mux27~2_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[22][4]~q ))) # (!cuifregS_2 & (\registerArray[18][4]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[18][4]~q ),
	.datac(\registerArray[22][4]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux27~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~2 .lut_mask = 16'hFA44;
defparam \Mux27~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N16
cycloneive_lcell_comb \Mux27~3 (
// Equation(s):
// \Mux27~3_combout  = (cuifregS_3 & ((\Mux27~2_combout  & (\registerArray[30][4]~q )) # (!\Mux27~2_combout  & ((\registerArray[26][4]~q ))))) # (!cuifregS_3 & (((\Mux27~2_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[30][4]~q ),
	.datac(\registerArray[26][4]~q ),
	.datad(\Mux27~2_combout ),
	.cin(gnd),
	.combout(\Mux27~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~3 .lut_mask = 16'hDDA0;
defparam \Mux27~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y34_N15
dffeas \registerArray[28][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][4] .is_wysiwyg = "true";
defparam \registerArray[28][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N25
dffeas \registerArray[24][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][4] .is_wysiwyg = "true";
defparam \registerArray[24][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N1
dffeas \registerArray[16][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][4] .is_wysiwyg = "true";
defparam \registerArray[16][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N11
dffeas \registerArray[20][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][4] .is_wysiwyg = "true";
defparam \registerArray[20][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N10
cycloneive_lcell_comb \Mux27~4 (
// Equation(s):
// \Mux27~4_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[20][4]~q ))) # (!cuifregS_2 & (\registerArray[16][4]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[16][4]~q ),
	.datac(\registerArray[20][4]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux27~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~4 .lut_mask = 16'hFA44;
defparam \Mux27~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N24
cycloneive_lcell_comb \Mux27~5 (
// Equation(s):
// \Mux27~5_combout  = (cuifregS_3 & ((\Mux27~4_combout  & (\registerArray[28][4]~q )) # (!\Mux27~4_combout  & ((\registerArray[24][4]~q ))))) # (!cuifregS_3 & (((\Mux27~4_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[28][4]~q ),
	.datac(\registerArray[24][4]~q ),
	.datad(\Mux27~4_combout ),
	.cin(gnd),
	.combout(\Mux27~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~5 .lut_mask = 16'hDDA0;
defparam \Mux27~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N30
cycloneive_lcell_comb \Mux27~6 (
// Equation(s):
// \Mux27~6_combout  = (cuifregS_0 & (cuifregS_1)) # (!cuifregS_0 & ((cuifregS_1 & (\Mux27~3_combout )) # (!cuifregS_1 & ((\Mux27~5_combout )))))

	.dataa(cuifregS_0),
	.datab(cuifregS_1),
	.datac(\Mux27~3_combout ),
	.datad(\Mux27~5_combout ),
	.cin(gnd),
	.combout(\Mux27~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~6 .lut_mask = 16'hD9C8;
defparam \Mux27~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N4
cycloneive_lcell_comb \registerArray[23][4]~feeder (
// Equation(s):
// \registerArray[23][4]~feeder_combout  = \Mux64~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux64),
	.cin(gnd),
	.combout(\registerArray[23][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[23][4]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[23][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y40_N5
dffeas \registerArray[23][4] (
	.clk(clk),
	.d(\registerArray[23][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][4] .is_wysiwyg = "true";
defparam \registerArray[23][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N31
dffeas \registerArray[19][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][4] .is_wysiwyg = "true";
defparam \registerArray[19][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N21
dffeas \registerArray[27][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][4] .is_wysiwyg = "true";
defparam \registerArray[27][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N20
cycloneive_lcell_comb \Mux27~7 (
// Equation(s):
// \Mux27~7_combout  = (cuifregS_3 & (((\registerArray[27][4]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[19][4]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[19][4]~q ),
	.datac(\registerArray[27][4]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux27~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~7 .lut_mask = 16'hAAE4;
defparam \Mux27~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y37_N2
cycloneive_lcell_comb \Mux27~8 (
// Equation(s):
// \Mux27~8_combout  = (cuifregS_2 & ((\Mux27~7_combout  & (\registerArray[31][4]~q )) # (!\Mux27~7_combout  & ((\registerArray[23][4]~q ))))) # (!cuifregS_2 & (((\Mux27~7_combout ))))

	.dataa(\registerArray[31][4]~q ),
	.datab(\registerArray[23][4]~q ),
	.datac(cuifregS_2),
	.datad(\Mux27~7_combout ),
	.cin(gnd),
	.combout(\Mux27~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~8 .lut_mask = 16'hAFC0;
defparam \Mux27~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N24
cycloneive_lcell_comb \Mux27~9 (
// Equation(s):
// \Mux27~9_combout  = (cuifregS_0 & ((\Mux27~6_combout  & ((\Mux27~8_combout ))) # (!\Mux27~6_combout  & (\Mux27~1_combout )))) # (!cuifregS_0 & (((\Mux27~6_combout ))))

	.dataa(cuifregS_0),
	.datab(\Mux27~1_combout ),
	.datac(\Mux27~6_combout ),
	.datad(\Mux27~8_combout ),
	.cin(gnd),
	.combout(\Mux27~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~9 .lut_mask = 16'hF858;
defparam \Mux27~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y31_N3
dffeas \registerArray[29][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][3] .is_wysiwyg = "true";
defparam \registerArray[29][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y31_N29
dffeas \registerArray[21][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][3] .is_wysiwyg = "true";
defparam \registerArray[21][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N28
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (cuifregS_2 & (((\registerArray[21][3]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[17][3]~q  & ((!cuifregS_3))))

	.dataa(\registerArray[17][3]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[21][3]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'hCCE2;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N8
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// \Mux28~1_combout  = (cuifregS_3 & ((\Mux28~0_combout  & ((\registerArray[29][3]~q ))) # (!\Mux28~0_combout  & (\registerArray[25][3]~q )))) # (!cuifregS_3 & (((\Mux28~0_combout ))))

	.dataa(\registerArray[25][3]~q ),
	.datab(\registerArray[29][3]~q ),
	.datac(cuifregS_3),
	.datad(\Mux28~0_combout ),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hCFA0;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y31_N9
dffeas \registerArray[30][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~65_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[30][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[30][3] .is_wysiwyg = "true";
defparam \registerArray[30][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N5
dffeas \registerArray[22][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][3] .is_wysiwyg = "true";
defparam \registerArray[22][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N4
cycloneive_lcell_comb \Mux28~3 (
// Equation(s):
// \Mux28~3_combout  = (\Mux28~2_combout  & ((\registerArray[30][3]~q ) # ((!cuifregS_2)))) # (!\Mux28~2_combout  & (((\registerArray[22][3]~q  & cuifregS_2))))

	.dataa(\Mux28~2_combout ),
	.datab(\registerArray[30][3]~q ),
	.datac(\registerArray[22][3]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux28~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~3 .lut_mask = 16'hD8AA;
defparam \Mux28~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N25
dffeas \registerArray[16][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][3] .is_wysiwyg = "true";
defparam \registerArray[16][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N15
dffeas \registerArray[24][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][3] .is_wysiwyg = "true";
defparam \registerArray[24][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N14
cycloneive_lcell_comb \Mux28~4 (
// Equation(s):
// \Mux28~4_combout  = (cuifregS_3 & (((\registerArray[24][3]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[16][3]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[16][3]~q ),
	.datac(\registerArray[24][3]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux28~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~4 .lut_mask = 16'hAAE4;
defparam \Mux28~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N17
dffeas \registerArray[20][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][3] .is_wysiwyg = "true";
defparam \registerArray[20][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N16
cycloneive_lcell_comb \Mux28~5 (
// Equation(s):
// \Mux28~5_combout  = (\Mux28~4_combout  & ((\registerArray[28][3]~q ) # ((!cuifregS_2)))) # (!\Mux28~4_combout  & (((\registerArray[20][3]~q  & cuifregS_2))))

	.dataa(\registerArray[28][3]~q ),
	.datab(\Mux28~4_combout ),
	.datac(\registerArray[20][3]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux28~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~5 .lut_mask = 16'hB8CC;
defparam \Mux28~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N8
cycloneive_lcell_comb \Mux28~6 (
// Equation(s):
// \Mux28~6_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\Mux28~3_combout )) # (!cuifregS_1 & ((\Mux28~5_combout )))))

	.dataa(cuifregS_0),
	.datab(\Mux28~3_combout ),
	.datac(cuifregS_1),
	.datad(\Mux28~5_combout ),
	.cin(gnd),
	.combout(\Mux28~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~6 .lut_mask = 16'hE5E0;
defparam \Mux28~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N22
cycloneive_lcell_comb \registerArray[27][3]~feeder (
// Equation(s):
// \registerArray[27][3]~feeder_combout  = \Mux65~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux65),
	.cin(gnd),
	.combout(\registerArray[27][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[27][3]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[27][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N23
dffeas \registerArray[27][3] (
	.clk(clk),
	.d(\registerArray[27][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][3] .is_wysiwyg = "true";
defparam \registerArray[27][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N1
dffeas \registerArray[23][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][3] .is_wysiwyg = "true";
defparam \registerArray[23][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N0
cycloneive_lcell_comb \Mux28~7 (
// Equation(s):
// \Mux28~7_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[23][3]~q ))) # (!cuifregS_2 & (\registerArray[19][3]~q ))))

	.dataa(\registerArray[19][3]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[23][3]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux28~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~7 .lut_mask = 16'hFC22;
defparam \Mux28~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N2
cycloneive_lcell_comb \Mux28~8 (
// Equation(s):
// \Mux28~8_combout  = (cuifregS_3 & ((\Mux28~7_combout  & (\registerArray[31][3]~q )) # (!\Mux28~7_combout  & ((\registerArray[27][3]~q ))))) # (!cuifregS_3 & (((\Mux28~7_combout ))))

	.dataa(\registerArray[31][3]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[27][3]~q ),
	.datad(\Mux28~7_combout ),
	.cin(gnd),
	.combout(\Mux28~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~8 .lut_mask = 16'hBBC0;
defparam \Mux28~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N26
cycloneive_lcell_comb \Mux28~9 (
// Equation(s):
// \Mux28~9_combout  = (cuifregS_0 & ((\Mux28~6_combout  & ((\Mux28~8_combout ))) # (!\Mux28~6_combout  & (\Mux28~1_combout )))) # (!cuifregS_0 & (((\Mux28~6_combout ))))

	.dataa(cuifregS_0),
	.datab(\Mux28~1_combout ),
	.datac(\Mux28~6_combout ),
	.datad(\Mux28~8_combout ),
	.cin(gnd),
	.combout(\Mux28~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~9 .lut_mask = 16'hF858;
defparam \Mux28~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N15
dffeas \registerArray[10][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][3] .is_wysiwyg = "true";
defparam \registerArray[10][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N0
cycloneive_lcell_comb \registerArray[8][3]~feeder (
// Equation(s):
// \registerArray[8][3]~feeder_combout  = \Mux65~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux65),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[8][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[8][3]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[8][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N1
dffeas \registerArray[8][3] (
	.clk(clk),
	.d(\registerArray[8][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][3] .is_wysiwyg = "true";
defparam \registerArray[8][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N14
cycloneive_lcell_comb \Mux28~10 (
// Equation(s):
// \Mux28~10_combout  = (cuifregS_1 & ((cuifregS_0) # ((\registerArray[10][3]~q )))) # (!cuifregS_1 & (!cuifregS_0 & ((\registerArray[8][3]~q ))))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\registerArray[10][3]~q ),
	.datad(\registerArray[8][3]~q ),
	.cin(gnd),
	.combout(\Mux28~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~10 .lut_mask = 16'hB9A8;
defparam \Mux28~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N21
dffeas \registerArray[9][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][3] .is_wysiwyg = "true";
defparam \registerArray[9][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N20
cycloneive_lcell_comb \Mux28~11 (
// Equation(s):
// \Mux28~11_combout  = (\Mux28~10_combout  & ((\registerArray[11][3]~q ) # ((!cuifregS_0)))) # (!\Mux28~10_combout  & (((\registerArray[9][3]~q  & cuifregS_0))))

	.dataa(\registerArray[11][3]~q ),
	.datab(\Mux28~10_combout ),
	.datac(\registerArray[9][3]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux28~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~11 .lut_mask = 16'hB8CC;
defparam \Mux28~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N26
cycloneive_lcell_comb \registerArray[15][3]~feeder (
// Equation(s):
// \registerArray[15][3]~feeder_combout  = \Mux65~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux65),
	.cin(gnd),
	.combout(\registerArray[15][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[15][3]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[15][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N27
dffeas \registerArray[15][3] (
	.clk(clk),
	.d(\registerArray[15][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][3] .is_wysiwyg = "true";
defparam \registerArray[15][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y36_N7
dffeas \registerArray[13][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][3] .is_wysiwyg = "true";
defparam \registerArray[13][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N12
cycloneive_lcell_comb \Mux28~17 (
// Equation(s):
// \Mux28~17_combout  = (cuifregS_0 & (((\registerArray[13][3]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[12][3]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[12][3]~q ),
	.datab(\registerArray[13][3]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux28~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~17 .lut_mask = 16'hF0CA;
defparam \Mux28~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N22
cycloneive_lcell_comb \Mux28~18 (
// Equation(s):
// \Mux28~18_combout  = (cuifregS_1 & ((\Mux28~17_combout  & ((\registerArray[15][3]~q ))) # (!\Mux28~17_combout  & (\registerArray[14][3]~q )))) # (!cuifregS_1 & (((\Mux28~17_combout ))))

	.dataa(\registerArray[14][3]~q ),
	.datab(\registerArray[15][3]~q ),
	.datac(cuifregS_1),
	.datad(\Mux28~17_combout ),
	.cin(gnd),
	.combout(\Mux28~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~18 .lut_mask = 16'hCFA0;
defparam \Mux28~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N9
dffeas \registerArray[6][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][3] .is_wysiwyg = "true";
defparam \registerArray[6][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N3
dffeas \registerArray[7][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][3] .is_wysiwyg = "true";
defparam \registerArray[7][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y35_N23
dffeas \registerArray[4][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][3] .is_wysiwyg = "true";
defparam \registerArray[4][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N22
cycloneive_lcell_comb \Mux28~12 (
// Equation(s):
// \Mux28~12_combout  = (cuifregS_0 & ((\registerArray[5][3]~q ) # ((cuifregS_1)))) # (!cuifregS_0 & (((\registerArray[4][3]~q  & !cuifregS_1))))

	.dataa(\registerArray[5][3]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[4][3]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux28~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~12 .lut_mask = 16'hCCB8;
defparam \Mux28~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N2
cycloneive_lcell_comb \Mux28~13 (
// Equation(s):
// \Mux28~13_combout  = (cuifregS_1 & ((\Mux28~12_combout  & ((\registerArray[7][3]~q ))) # (!\Mux28~12_combout  & (\registerArray[6][3]~q )))) # (!cuifregS_1 & (((\Mux28~12_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[6][3]~q ),
	.datac(\registerArray[7][3]~q ),
	.datad(\Mux28~12_combout ),
	.cin(gnd),
	.combout(\Mux28~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~13 .lut_mask = 16'hF588;
defparam \Mux28~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y43_N1
dffeas \registerArray[1][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][3] .is_wysiwyg = "true";
defparam \registerArray[1][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y43_N31
dffeas \registerArray[3][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][3] .is_wysiwyg = "true";
defparam \registerArray[3][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N0
cycloneive_lcell_comb \Mux28~14 (
// Equation(s):
// \Mux28~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][3]~q ))) # (!cuifregS_1 & (\registerArray[1][3]~q ))))

	.dataa(cuifregS_0),
	.datab(cuifregS_1),
	.datac(\registerArray[1][3]~q ),
	.datad(\registerArray[3][3]~q ),
	.cin(gnd),
	.combout(\Mux28~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~14 .lut_mask = 16'hA820;
defparam \Mux28~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N12
cycloneive_lcell_comb \Mux28~15 (
// Equation(s):
// \Mux28~15_combout  = (\Mux28~14_combout ) # ((\registerArray[2][3]~q  & (!cuifregS_0 & cuifregS_1)))

	.dataa(\registerArray[2][3]~q ),
	.datab(cuifregS_0),
	.datac(\Mux28~14_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux28~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~15 .lut_mask = 16'hF2F0;
defparam \Mux28~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N2
cycloneive_lcell_comb \Mux28~16 (
// Equation(s):
// \Mux28~16_combout  = (cuifregS_2 & ((cuifregS_3) # ((\Mux28~13_combout )))) # (!cuifregS_2 & (!cuifregS_3 & ((\Mux28~15_combout ))))

	.dataa(cuifregS_2),
	.datab(cuifregS_3),
	.datac(\Mux28~13_combout ),
	.datad(\Mux28~15_combout ),
	.cin(gnd),
	.combout(\Mux28~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~16 .lut_mask = 16'hB9A8;
defparam \Mux28~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N28
cycloneive_lcell_comb \Mux28~19 (
// Equation(s):
// \Mux28~19_combout  = (cuifregS_3 & ((\Mux28~16_combout  & ((\Mux28~18_combout ))) # (!\Mux28~16_combout  & (\Mux28~11_combout )))) # (!cuifregS_3 & (((\Mux28~16_combout ))))

	.dataa(\Mux28~11_combout ),
	.datab(cuifregS_3),
	.datac(\Mux28~18_combout ),
	.datad(\Mux28~16_combout ),
	.cin(gnd),
	.combout(\Mux28~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~19 .lut_mask = 16'hF388;
defparam \Mux28~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N12
cycloneive_lcell_comb \Mux61~4 (
// Equation(s):
// \Mux61~4_combout  = (cuifregT_3 & ((\registerArray[24][2]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[16][2]~q  & !cuifregT_2))))

	.dataa(cuifregT_3),
	.datab(\registerArray[24][2]~q ),
	.datac(\registerArray[16][2]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux61~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~4 .lut_mask = 16'hAAD8;
defparam \Mux61~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N14
cycloneive_lcell_comb \Mux61~5 (
// Equation(s):
// \Mux61~5_combout  = (cuifregT_2 & ((\Mux61~4_combout  & ((\registerArray[28][2]~q ))) # (!\Mux61~4_combout  & (\registerArray[20][2]~q )))) # (!cuifregT_2 & (((\Mux61~4_combout ))))

	.dataa(\registerArray[20][2]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[28][2]~q ),
	.datad(\Mux61~4_combout ),
	.cin(gnd),
	.combout(\Mux61~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~5 .lut_mask = 16'hF388;
defparam \Mux61~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y31_N29
dffeas \registerArray[18][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][2] .is_wysiwyg = "true";
defparam \registerArray[18][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N28
cycloneive_lcell_comb \Mux61~2 (
// Equation(s):
// \Mux61~2_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[26][2]~q )) # (!cuifregT_3 & ((\registerArray[18][2]~q )))))

	.dataa(\registerArray[26][2]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[18][2]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux61~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~2 .lut_mask = 16'hEE30;
defparam \Mux61~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N2
cycloneive_lcell_comb \Mux61~3 (
// Equation(s):
// \Mux61~3_combout  = (cuifregT_2 & ((\Mux61~2_combout  & ((\registerArray[30][2]~q ))) # (!\Mux61~2_combout  & (\registerArray[22][2]~q )))) # (!cuifregT_2 & (((\Mux61~2_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[22][2]~q ),
	.datac(\registerArray[30][2]~q ),
	.datad(\Mux61~2_combout ),
	.cin(gnd),
	.combout(\Mux61~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~3 .lut_mask = 16'hF588;
defparam \Mux61~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N4
cycloneive_lcell_comb \Mux61~6 (
// Equation(s):
// \Mux61~6_combout  = (cuifregT_01 & (cuifregT_1)) # (!cuifregT_01 & ((cuifregT_1 & ((\Mux61~3_combout ))) # (!cuifregT_1 & (\Mux61~5_combout ))))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\Mux61~5_combout ),
	.datad(\Mux61~3_combout ),
	.cin(gnd),
	.combout(\Mux61~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~6 .lut_mask = 16'hDC98;
defparam \Mux61~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N24
cycloneive_lcell_comb \registerArray[23][2]~feeder (
// Equation(s):
// \registerArray[23][2]~feeder_combout  = \Mux66~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux66),
	.cin(gnd),
	.combout(\registerArray[23][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[23][2]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[23][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N25
dffeas \registerArray[23][2] (
	.clk(clk),
	.d(\registerArray[23][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][2] .is_wysiwyg = "true";
defparam \registerArray[23][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N24
cycloneive_lcell_comb \Mux61~7 (
// Equation(s):
// \Mux61~7_combout  = (cuifregT_2 & ((\registerArray[23][2]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[19][2]~q  & !cuifregT_3))))

	.dataa(cuifregT_2),
	.datab(\registerArray[23][2]~q ),
	.datac(\registerArray[19][2]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux61~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~7 .lut_mask = 16'hAAD8;
defparam \Mux61~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N28
cycloneive_lcell_comb \Mux61~8 (
// Equation(s):
// \Mux61~8_combout  = (cuifregT_3 & ((\Mux61~7_combout  & ((\registerArray[31][2]~q ))) # (!\Mux61~7_combout  & (\registerArray[27][2]~q )))) # (!cuifregT_3 & (((\Mux61~7_combout ))))

	.dataa(\registerArray[27][2]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[31][2]~q ),
	.datad(\Mux61~7_combout ),
	.cin(gnd),
	.combout(\Mux61~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~8 .lut_mask = 16'hF388;
defparam \Mux61~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N10
cycloneive_lcell_comb \registerArray[29][2]~feeder (
// Equation(s):
// \registerArray[29][2]~feeder_combout  = \Mux66~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux66),
	.cin(gnd),
	.combout(\registerArray[29][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[29][2]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[29][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N11
dffeas \registerArray[29][2] (
	.clk(clk),
	.d(\registerArray[29][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][2] .is_wysiwyg = "true";
defparam \registerArray[29][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N14
cycloneive_lcell_comb \registerArray[25][2]~feeder (
// Equation(s):
// \registerArray[25][2]~feeder_combout  = \Mux66~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux66),
	.cin(gnd),
	.combout(\registerArray[25][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[25][2]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[25][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N15
dffeas \registerArray[25][2] (
	.clk(clk),
	.d(\registerArray[25][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][2] .is_wysiwyg = "true";
defparam \registerArray[25][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N8
cycloneive_lcell_comb \Mux61~0 (
// Equation(s):
// \Mux61~0_combout  = (cuifregT_2 & ((\registerArray[21][2]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[17][2]~q  & !cuifregT_3))))

	.dataa(cuifregT_2),
	.datab(\registerArray[21][2]~q ),
	.datac(\registerArray[17][2]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux61~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~0 .lut_mask = 16'hAAD8;
defparam \Mux61~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N12
cycloneive_lcell_comb \Mux61~1 (
// Equation(s):
// \Mux61~1_combout  = (cuifregT_3 & ((\Mux61~0_combout  & (\registerArray[29][2]~q )) # (!\Mux61~0_combout  & ((\registerArray[25][2]~q ))))) # (!cuifregT_3 & (((\Mux61~0_combout ))))

	.dataa(\registerArray[29][2]~q ),
	.datab(\registerArray[25][2]~q ),
	.datac(cuifregT_3),
	.datad(\Mux61~0_combout ),
	.cin(gnd),
	.combout(\Mux61~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~1 .lut_mask = 16'hAFC0;
defparam \Mux61~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N28
cycloneive_lcell_comb \registerArray[10][2]~feeder (
// Equation(s):
// \registerArray[10][2]~feeder_combout  = \Mux66~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux66),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[10][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[10][2]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[10][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N29
dffeas \registerArray[10][2] (
	.clk(clk),
	.d(\registerArray[10][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][2] .is_wysiwyg = "true";
defparam \registerArray[10][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N12
cycloneive_lcell_comb \Mux61~10 (
// Equation(s):
// \Mux61~10_combout  = (cuifregT_1 & (((\registerArray[10][2]~q ) # (cuifregT_01)))) # (!cuifregT_1 & (\registerArray[8][2]~q  & ((!cuifregT_01))))

	.dataa(\registerArray[8][2]~q ),
	.datab(\registerArray[10][2]~q ),
	.datac(cuifregT_1),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux61~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~10 .lut_mask = 16'hF0CA;
defparam \Mux61~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N8
cycloneive_lcell_comb \Mux61~11 (
// Equation(s):
// \Mux61~11_combout  = (cuifregT_01 & ((\Mux61~10_combout  & (\registerArray[11][2]~q )) # (!\Mux61~10_combout  & ((\registerArray[9][2]~q ))))) # (!cuifregT_01 & (((\Mux61~10_combout ))))

	.dataa(cuifregT_0),
	.datab(\registerArray[11][2]~q ),
	.datac(\registerArray[9][2]~q ),
	.datad(\Mux61~10_combout ),
	.cin(gnd),
	.combout(\Mux61~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~11 .lut_mask = 16'hDDA0;
defparam \Mux61~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N3
dffeas \registerArray[15][2] (
	.clk(clk),
	.d(Mux66),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~84_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[15][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[15][2] .is_wysiwyg = "true";
defparam \registerArray[15][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N14
cycloneive_lcell_comb \Mux61~17 (
// Equation(s):
// \Mux61~17_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & ((\registerArray[13][2]~q ))) # (!cuifregT_01 & (\registerArray[12][2]~q ))))

	.dataa(\registerArray[12][2]~q ),
	.datab(\registerArray[13][2]~q ),
	.datac(cuifregT_1),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux61~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~17 .lut_mask = 16'hFC0A;
defparam \Mux61~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N26
cycloneive_lcell_comb \Mux61~18 (
// Equation(s):
// \Mux61~18_combout  = (cuifregT_1 & ((\Mux61~17_combout  & ((\registerArray[15][2]~q ))) # (!\Mux61~17_combout  & (\registerArray[14][2]~q )))) # (!cuifregT_1 & (((\Mux61~17_combout ))))

	.dataa(\registerArray[14][2]~q ),
	.datab(\registerArray[15][2]~q ),
	.datac(cuifregT_1),
	.datad(\Mux61~17_combout ),
	.cin(gnd),
	.combout(\Mux61~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~18 .lut_mask = 16'hCFA0;
defparam \Mux61~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N11
dffeas \registerArray[4][2] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux66),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][2] .is_wysiwyg = "true";
defparam \registerArray[4][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N10
cycloneive_lcell_comb \Mux61~12 (
// Equation(s):
// \Mux61~12_combout  = (cuifregT_01 & ((\registerArray[5][2]~q ) # ((cuifregT_1)))) # (!cuifregT_01 & (((\registerArray[4][2]~q  & !cuifregT_1))))

	.dataa(cuifregT_0),
	.datab(\registerArray[5][2]~q ),
	.datac(\registerArray[4][2]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux61~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~12 .lut_mask = 16'hAAD8;
defparam \Mux61~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N16
cycloneive_lcell_comb \Mux61~13 (
// Equation(s):
// \Mux61~13_combout  = (cuifregT_1 & ((\Mux61~12_combout  & (\registerArray[7][2]~q )) # (!\Mux61~12_combout  & ((\registerArray[6][2]~q ))))) # (!cuifregT_1 & (((\Mux61~12_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[7][2]~q ),
	.datac(\registerArray[6][2]~q ),
	.datad(\Mux61~12_combout ),
	.cin(gnd),
	.combout(\Mux61~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~13 .lut_mask = 16'hDDA0;
defparam \Mux61~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N8
cycloneive_lcell_comb \registerArray[3][2]~feeder (
// Equation(s):
// \registerArray[3][2]~feeder_combout  = \Mux66~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux66),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[3][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[3][2]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[3][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y42_N9
dffeas \registerArray[3][2] (
	.clk(clk),
	.d(\registerArray[3][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][2] .is_wysiwyg = "true";
defparam \registerArray[3][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N4
cycloneive_lcell_comb \Mux61~14 (
// Equation(s):
// \Mux61~14_combout  = (cuifregT_01 & ((cuifregT_1 & ((\registerArray[3][2]~q ))) # (!cuifregT_1 & (\registerArray[1][2]~q ))))

	.dataa(\registerArray[1][2]~q ),
	.datab(\registerArray[3][2]~q ),
	.datac(cuifregT_1),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux61~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~14 .lut_mask = 16'hCA00;
defparam \Mux61~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N18
cycloneive_lcell_comb \Mux61~15 (
// Equation(s):
// \Mux61~15_combout  = (\Mux61~14_combout ) # ((!cuifregT_01 & (cuifregT_1 & \registerArray[2][2]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\Mux61~14_combout ),
	.datad(\registerArray[2][2]~q ),
	.cin(gnd),
	.combout(\Mux61~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~15 .lut_mask = 16'hF4F0;
defparam \Mux61~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N16
cycloneive_lcell_comb \Mux61~16 (
// Equation(s):
// \Mux61~16_combout  = (cuifregT_3 & (cuifregT_2)) # (!cuifregT_3 & ((cuifregT_2 & (\Mux61~13_combout )) # (!cuifregT_2 & ((\Mux61~15_combout )))))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\Mux61~13_combout ),
	.datad(\Mux61~15_combout ),
	.cin(gnd),
	.combout(\Mux61~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~16 .lut_mask = 16'hD9C8;
defparam \Mux61~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N0
cycloneive_lcell_comb \registerArray[21][8]~feeder (
// Equation(s):
// \registerArray[21][8]~feeder_combout  = \Mux60~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux602),
	.cin(gnd),
	.combout(\registerArray[21][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[21][8]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[21][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y37_N1
dffeas \registerArray[21][8] (
	.clk(clk),
	.d(\registerArray[21][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][8] .is_wysiwyg = "true";
defparam \registerArray[21][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N30
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// \Mux23~0_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & (\registerArray[25][8]~q )) # (!cuifregS_3 & ((\registerArray[17][8]~q )))))

	.dataa(\registerArray[25][8]~q ),
	.datab(\registerArray[17][8]~q ),
	.datac(cuifregS_2),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hFA0C;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N20
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// \Mux23~1_combout  = (cuifregS_2 & ((\Mux23~0_combout  & (\registerArray[29][8]~q )) # (!\Mux23~0_combout  & ((\registerArray[21][8]~q ))))) # (!cuifregS_2 & (((\Mux23~0_combout ))))

	.dataa(\registerArray[29][8]~q ),
	.datab(\registerArray[21][8]~q ),
	.datac(cuifregS_2),
	.datad(\Mux23~0_combout ),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'hAFC0;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y35_N27
dffeas \registerArray[16][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][8] .is_wysiwyg = "true";
defparam \registerArray[16][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N8
cycloneive_lcell_comb \Mux23~4 (
// Equation(s):
// \Mux23~4_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[20][8]~q ))) # (!cuifregS_2 & (\registerArray[16][8]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[16][8]~q ),
	.datac(\registerArray[20][8]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux23~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~4 .lut_mask = 16'hFA44;
defparam \Mux23~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N28
cycloneive_lcell_comb \Mux23~5 (
// Equation(s):
// \Mux23~5_combout  = (cuifregS_3 & ((\Mux23~4_combout  & ((\registerArray[28][8]~q ))) # (!\Mux23~4_combout  & (\registerArray[24][8]~q )))) # (!cuifregS_3 & (((\Mux23~4_combout ))))

	.dataa(\registerArray[24][8]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[28][8]~q ),
	.datad(\Mux23~4_combout ),
	.cin(gnd),
	.combout(\Mux23~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~5 .lut_mask = 16'hF388;
defparam \Mux23~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N14
cycloneive_lcell_comb \Mux23~6 (
// Equation(s):
// \Mux23~6_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\Mux23~3_combout )) # (!cuifregS_1 & ((\Mux23~5_combout )))))

	.dataa(\Mux23~3_combout ),
	.datab(cuifregS_0),
	.datac(cuifregS_1),
	.datad(\Mux23~5_combout ),
	.cin(gnd),
	.combout(\Mux23~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~6 .lut_mask = 16'hE3E0;
defparam \Mux23~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N0
cycloneive_lcell_comb \Mux23~7 (
// Equation(s):
// \Mux23~7_combout  = (cuifregS_3 & (((\registerArray[27][8]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[19][8]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[19][8]~q ),
	.datac(\registerArray[27][8]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux23~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~7 .lut_mask = 16'hAAE4;
defparam \Mux23~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N18
cycloneive_lcell_comb \Mux23~8 (
// Equation(s):
// \Mux23~8_combout  = (cuifregS_2 & ((\Mux23~7_combout  & ((\registerArray[31][8]~q ))) # (!\Mux23~7_combout  & (\registerArray[23][8]~q )))) # (!cuifregS_2 & (((\Mux23~7_combout ))))

	.dataa(\registerArray[23][8]~q ),
	.datab(\registerArray[31][8]~q ),
	.datac(cuifregS_2),
	.datad(\Mux23~7_combout ),
	.cin(gnd),
	.combout(\Mux23~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~8 .lut_mask = 16'hCFA0;
defparam \Mux23~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N4
cycloneive_lcell_comb \Mux23~9 (
// Equation(s):
// \Mux23~9_combout  = (cuifregS_0 & ((\Mux23~6_combout  & ((\Mux23~8_combout ))) # (!\Mux23~6_combout  & (\Mux23~1_combout )))) # (!cuifregS_0 & (((\Mux23~6_combout ))))

	.dataa(\Mux23~1_combout ),
	.datab(cuifregS_0),
	.datac(\Mux23~6_combout ),
	.datad(\Mux23~8_combout ),
	.cin(gnd),
	.combout(\Mux23~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~9 .lut_mask = 16'hF838;
defparam \Mux23~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N29
dffeas \registerArray[3][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][8] .is_wysiwyg = "true";
defparam \registerArray[3][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N28
cycloneive_lcell_comb \Mux23~14 (
// Equation(s):
// \Mux23~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][8]~q ))) # (!cuifregS_1 & (\registerArray[1][8]~q ))))

	.dataa(\registerArray[1][8]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[3][8]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux23~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~14 .lut_mask = 16'hC088;
defparam \Mux23~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N22
cycloneive_lcell_comb \Mux23~15 (
// Equation(s):
// \Mux23~15_combout  = (\Mux23~14_combout ) # ((\registerArray[2][8]~q  & (cuifregS_1 & !cuifregS_0)))

	.dataa(\registerArray[2][8]~q ),
	.datab(cuifregS_1),
	.datac(\Mux23~14_combout ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux23~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~15 .lut_mask = 16'hF0F8;
defparam \Mux23~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N19
dffeas \registerArray[10][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][8] .is_wysiwyg = "true";
defparam \registerArray[10][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N18
cycloneive_lcell_comb \Mux23~12 (
// Equation(s):
// \Mux23~12_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][8]~q ))) # (!cuifregS_1 & (\registerArray[8][8]~q ))))

	.dataa(\registerArray[8][8]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[10][8]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux23~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~12 .lut_mask = 16'hFC22;
defparam \Mux23~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N8
cycloneive_lcell_comb \Mux23~13 (
// Equation(s):
// \Mux23~13_combout  = (cuifregS_0 & ((\Mux23~12_combout  & (\registerArray[11][8]~q )) # (!\Mux23~12_combout  & ((\registerArray[9][8]~q ))))) # (!cuifregS_0 & (((\Mux23~12_combout ))))

	.dataa(\registerArray[11][8]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[9][8]~q ),
	.datad(\Mux23~12_combout ),
	.cin(gnd),
	.combout(\Mux23~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~13 .lut_mask = 16'hBBC0;
defparam \Mux23~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N0
cycloneive_lcell_comb \Mux23~16 (
// Equation(s):
// \Mux23~16_combout  = (cuifregS_2 & (cuifregS_3)) # (!cuifregS_2 & ((cuifregS_3 & ((\Mux23~13_combout ))) # (!cuifregS_3 & (\Mux23~15_combout ))))

	.dataa(cuifregS_2),
	.datab(cuifregS_3),
	.datac(\Mux23~15_combout ),
	.datad(\Mux23~13_combout ),
	.cin(gnd),
	.combout(\Mux23~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~16 .lut_mask = 16'hDC98;
defparam \Mux23~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y33_N5
dffeas \registerArray[13][8] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux602),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][8] .is_wysiwyg = "true";
defparam \registerArray[13][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N8
cycloneive_lcell_comb \Mux23~17 (
// Equation(s):
// \Mux23~17_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & (\registerArray[13][8]~q )) # (!cuifregS_0 & ((\registerArray[12][8]~q )))))

	.dataa(cuifregS_1),
	.datab(\registerArray[13][8]~q ),
	.datac(\registerArray[12][8]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux23~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~17 .lut_mask = 16'hEE50;
defparam \Mux23~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N2
cycloneive_lcell_comb \Mux23~18 (
// Equation(s):
// \Mux23~18_combout  = (\Mux23~17_combout  & (((\registerArray[15][8]~q ) # (!cuifregS_1)))) # (!\Mux23~17_combout  & (\registerArray[14][8]~q  & ((cuifregS_1))))

	.dataa(\registerArray[14][8]~q ),
	.datab(\registerArray[15][8]~q ),
	.datac(\Mux23~17_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux23~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~18 .lut_mask = 16'hCAF0;
defparam \Mux23~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N22
cycloneive_lcell_comb \Mux23~10 (
// Equation(s):
// \Mux23~10_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & (\registerArray[5][8]~q )) # (!cuifregS_0 & ((\registerArray[4][8]~q )))))

	.dataa(\registerArray[5][8]~q ),
	.datab(cuifregS_1),
	.datac(\registerArray[4][8]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux23~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~10 .lut_mask = 16'hEE30;
defparam \Mux23~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N8
cycloneive_lcell_comb \Mux23~11 (
// Equation(s):
// \Mux23~11_combout  = (\Mux23~10_combout  & ((\registerArray[7][8]~q ) # ((!cuifregS_1)))) # (!\Mux23~10_combout  & (((\registerArray[6][8]~q  & cuifregS_1))))

	.dataa(\registerArray[7][8]~q ),
	.datab(\registerArray[6][8]~q ),
	.datac(\Mux23~10_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux23~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~11 .lut_mask = 16'hACF0;
defparam \Mux23~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N2
cycloneive_lcell_comb \Mux23~19 (
// Equation(s):
// \Mux23~19_combout  = (cuifregS_2 & ((\Mux23~16_combout  & (\Mux23~18_combout )) # (!\Mux23~16_combout  & ((\Mux23~11_combout ))))) # (!cuifregS_2 & (\Mux23~16_combout ))

	.dataa(cuifregS_2),
	.datab(\Mux23~16_combout ),
	.datac(\Mux23~18_combout ),
	.datad(\Mux23~11_combout ),
	.cin(gnd),
	.combout(\Mux23~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~19 .lut_mask = 16'hE6C4;
defparam \Mux23~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N0
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[21][7]~q ))) # (!cuifregS_2 & (\registerArray[17][7]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[17][7]~q ),
	.datac(\registerArray[21][7]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'hFA44;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N18
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// \Mux24~1_combout  = (cuifregS_3 & ((\Mux24~0_combout  & ((\registerArray[29][7]~q ))) # (!\Mux24~0_combout  & (\registerArray[25][7]~q )))) # (!cuifregS_3 & (\Mux24~0_combout ))

	.dataa(cuifregS_3),
	.datab(\Mux24~0_combout ),
	.datac(\registerArray[25][7]~q ),
	.datad(\registerArray[29][7]~q ),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'hEC64;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N27
dffeas \registerArray[27][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][7] .is_wysiwyg = "true";
defparam \registerArray[27][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N16
cycloneive_lcell_comb \Mux24~7 (
// Equation(s):
// \Mux24~7_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[23][7]~q ))) # (!cuifregS_2 & (\registerArray[19][7]~q ))))

	.dataa(\registerArray[19][7]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[23][7]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux24~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~7 .lut_mask = 16'hFC22;
defparam \Mux24~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N26
cycloneive_lcell_comb \Mux24~8 (
// Equation(s):
// \Mux24~8_combout  = (cuifregS_3 & ((\Mux24~7_combout  & (\registerArray[31][7]~q )) # (!\Mux24~7_combout  & ((\registerArray[27][7]~q ))))) # (!cuifregS_3 & (((\Mux24~7_combout ))))

	.dataa(\registerArray[31][7]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[27][7]~q ),
	.datad(\Mux24~7_combout ),
	.cin(gnd),
	.combout(\Mux24~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~8 .lut_mask = 16'hBBC0;
defparam \Mux24~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N24
cycloneive_lcell_comb \registerArray[26][7]~feeder (
// Equation(s):
// \registerArray[26][7]~feeder_combout  = \Mux61~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux612),
	.cin(gnd),
	.combout(\registerArray[26][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[26][7]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[26][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N25
dffeas \registerArray[26][7] (
	.clk(clk),
	.d(\registerArray[26][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][7] .is_wysiwyg = "true";
defparam \registerArray[26][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N30
cycloneive_lcell_comb \Mux24~2 (
// Equation(s):
// \Mux24~2_combout  = (cuifregS_3 & (((\registerArray[26][7]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[18][7]~q  & ((!cuifregS_2))))

	.dataa(\registerArray[18][7]~q ),
	.datab(\registerArray[26][7]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux24~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~2 .lut_mask = 16'hF0CA;
defparam \Mux24~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N8
cycloneive_lcell_comb \Mux24~3 (
// Equation(s):
// \Mux24~3_combout  = (\Mux24~2_combout  & (((\registerArray[30][7]~q ) # (!cuifregS_2)))) # (!\Mux24~2_combout  & (\registerArray[22][7]~q  & ((cuifregS_2))))

	.dataa(\registerArray[22][7]~q ),
	.datab(\registerArray[30][7]~q ),
	.datac(\Mux24~2_combout ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux24~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~3 .lut_mask = 16'hCAF0;
defparam \Mux24~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y33_N27
dffeas \registerArray[20][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][7] .is_wysiwyg = "true";
defparam \registerArray[20][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N13
dffeas \registerArray[24][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][7] .is_wysiwyg = "true";
defparam \registerArray[24][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N12
cycloneive_lcell_comb \Mux24~4 (
// Equation(s):
// \Mux24~4_combout  = (cuifregS_3 & (((\registerArray[24][7]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[16][7]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[16][7]~q ),
	.datac(\registerArray[24][7]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux24~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~4 .lut_mask = 16'hAAE4;
defparam \Mux24~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N26
cycloneive_lcell_comb \Mux24~5 (
// Equation(s):
// \Mux24~5_combout  = (cuifregS_2 & ((\Mux24~4_combout  & (\registerArray[28][7]~q )) # (!\Mux24~4_combout  & ((\registerArray[20][7]~q ))))) # (!cuifregS_2 & (((\Mux24~4_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[28][7]~q ),
	.datac(\registerArray[20][7]~q ),
	.datad(\Mux24~4_combout ),
	.cin(gnd),
	.combout(\Mux24~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~5 .lut_mask = 16'hDDA0;
defparam \Mux24~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N28
cycloneive_lcell_comb \Mux24~6 (
// Equation(s):
// \Mux24~6_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\Mux24~3_combout )) # (!cuifregS_1 & ((\Mux24~5_combout )))))

	.dataa(cuifregS_0),
	.datab(\Mux24~3_combout ),
	.datac(cuifregS_1),
	.datad(\Mux24~5_combout ),
	.cin(gnd),
	.combout(\Mux24~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~6 .lut_mask = 16'hE5E0;
defparam \Mux24~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N30
cycloneive_lcell_comb \Mux24~9 (
// Equation(s):
// \Mux24~9_combout  = (cuifregS_0 & ((\Mux24~6_combout  & ((\Mux24~8_combout ))) # (!\Mux24~6_combout  & (\Mux24~1_combout )))) # (!cuifregS_0 & (((\Mux24~6_combout ))))

	.dataa(\Mux24~1_combout ),
	.datab(cuifregS_0),
	.datac(\Mux24~8_combout ),
	.datad(\Mux24~6_combout ),
	.cin(gnd),
	.combout(\Mux24~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~9 .lut_mask = 16'hF388;
defparam \Mux24~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N4
cycloneive_lcell_comb \Mux24~17 (
// Equation(s):
// \Mux24~17_combout  = (cuifregS_0 & (((\registerArray[13][7]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[12][7]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[12][7]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[13][7]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux24~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~17 .lut_mask = 16'hCCE2;
defparam \Mux24~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N6
cycloneive_lcell_comb \Mux24~18 (
// Equation(s):
// \Mux24~18_combout  = (cuifregS_1 & ((\Mux24~17_combout  & ((\registerArray[15][7]~q ))) # (!\Mux24~17_combout  & (\registerArray[14][7]~q )))) # (!cuifregS_1 & (((\Mux24~17_combout ))))

	.dataa(\registerArray[14][7]~q ),
	.datab(\registerArray[15][7]~q ),
	.datac(cuifregS_1),
	.datad(\Mux24~17_combout ),
	.cin(gnd),
	.combout(\Mux24~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~18 .lut_mask = 16'hCFA0;
defparam \Mux24~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N13
dffeas \registerArray[9][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][7] .is_wysiwyg = "true";
defparam \registerArray[9][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N12
cycloneive_lcell_comb \Mux24~11 (
// Equation(s):
// \Mux24~11_combout  = (\Mux24~10_combout  & (((\registerArray[11][7]~q )) # (!cuifregS_0))) # (!\Mux24~10_combout  & (cuifregS_0 & (\registerArray[9][7]~q )))

	.dataa(\Mux24~10_combout ),
	.datab(cuifregS_0),
	.datac(\registerArray[9][7]~q ),
	.datad(\registerArray[11][7]~q ),
	.cin(gnd),
	.combout(\Mux24~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~11 .lut_mask = 16'hEA62;
defparam \Mux24~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N25
dffeas \registerArray[5][7] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux612),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][7] .is_wysiwyg = "true";
defparam \registerArray[5][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N24
cycloneive_lcell_comb \Mux24~12 (
// Equation(s):
// \Mux24~12_combout  = (cuifregS_0 & (((\registerArray[5][7]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[4][7]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[4][7]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[5][7]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux24~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~12 .lut_mask = 16'hCCE2;
defparam \Mux24~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N20
cycloneive_lcell_comb \Mux24~13 (
// Equation(s):
// \Mux24~13_combout  = (cuifregS_1 & ((\Mux24~12_combout  & (\registerArray[7][7]~q )) # (!\Mux24~12_combout  & ((\registerArray[6][7]~q ))))) # (!cuifregS_1 & (((\Mux24~12_combout ))))

	.dataa(\registerArray[7][7]~q ),
	.datab(cuifregS_1),
	.datac(\registerArray[6][7]~q ),
	.datad(\Mux24~12_combout ),
	.cin(gnd),
	.combout(\Mux24~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~13 .lut_mask = 16'hBBC0;
defparam \Mux24~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N12
cycloneive_lcell_comb \Mux24~16 (
// Equation(s):
// \Mux24~16_combout  = (cuifregS_2 & (((cuifregS_3) # (\Mux24~13_combout )))) # (!cuifregS_2 & (\Mux24~15_combout  & (!cuifregS_3)))

	.dataa(\Mux24~15_combout ),
	.datab(cuifregS_2),
	.datac(cuifregS_3),
	.datad(\Mux24~13_combout ),
	.cin(gnd),
	.combout(\Mux24~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~16 .lut_mask = 16'hCEC2;
defparam \Mux24~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N16
cycloneive_lcell_comb \Mux24~19 (
// Equation(s):
// \Mux24~19_combout  = (cuifregS_3 & ((\Mux24~16_combout  & (\Mux24~18_combout )) # (!\Mux24~16_combout  & ((\Mux24~11_combout ))))) # (!cuifregS_3 & (((\Mux24~16_combout ))))

	.dataa(\Mux24~18_combout ),
	.datab(\Mux24~11_combout ),
	.datac(cuifregS_3),
	.datad(\Mux24~16_combout ),
	.cin(gnd),
	.combout(\Mux24~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~19 .lut_mask = 16'hAFC0;
defparam \Mux24~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N4
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (cuifregS_3 & (((\registerArray[25][6]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[17][6]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[17][6]~q ),
	.datac(\registerArray[25][6]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hAAE4;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N30
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// \Mux25~1_combout  = (\Mux25~0_combout  & ((\registerArray[29][6]~q ) # ((!cuifregS_2)))) # (!\Mux25~0_combout  & (((\registerArray[21][6]~q  & cuifregS_2))))

	.dataa(\registerArray[29][6]~q ),
	.datab(\Mux25~0_combout ),
	.datac(\registerArray[21][6]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hB8CC;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y31_N9
dffeas \registerArray[19][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][6] .is_wysiwyg = "true";
defparam \registerArray[19][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N8
cycloneive_lcell_comb \Mux25~7 (
// Equation(s):
// \Mux25~7_combout  = (cuifregS_3 & ((\registerArray[27][6]~q ) # ((cuifregS_2)))) # (!cuifregS_3 & (((\registerArray[19][6]~q  & !cuifregS_2))))

	.dataa(\registerArray[27][6]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[19][6]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux25~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~7 .lut_mask = 16'hCCB8;
defparam \Mux25~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N4
cycloneive_lcell_comb \Mux25~8 (
// Equation(s):
// \Mux25~8_combout  = (cuifregS_2 & ((\Mux25~7_combout  & (\registerArray[31][6]~q )) # (!\Mux25~7_combout  & ((\registerArray[23][6]~q ))))) # (!cuifregS_2 & (((\Mux25~7_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[31][6]~q ),
	.datac(\registerArray[23][6]~q ),
	.datad(\Mux25~7_combout ),
	.cin(gnd),
	.combout(\Mux25~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~8 .lut_mask = 16'hDDA0;
defparam \Mux25~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y41_N10
cycloneive_lcell_comb \registerArray[16][6]~feeder (
// Equation(s):
// \registerArray[16][6]~feeder_combout  = \Mux62~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux622),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[16][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[16][6]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[16][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y41_N11
dffeas \registerArray[16][6] (
	.clk(clk),
	.d(\registerArray[16][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][6] .is_wysiwyg = "true";
defparam \registerArray[16][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N21
dffeas \registerArray[20][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][6] .is_wysiwyg = "true";
defparam \registerArray[20][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N20
cycloneive_lcell_comb \Mux25~4 (
// Equation(s):
// \Mux25~4_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[20][6]~q ))) # (!cuifregS_2 & (\registerArray[16][6]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[16][6]~q ),
	.datac(\registerArray[20][6]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux25~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~4 .lut_mask = 16'hFA44;
defparam \Mux25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N6
cycloneive_lcell_comb \Mux25~5 (
// Equation(s):
// \Mux25~5_combout  = (cuifregS_3 & ((\Mux25~4_combout  & (\registerArray[28][6]~q )) # (!\Mux25~4_combout  & ((\registerArray[24][6]~q ))))) # (!cuifregS_3 & (((\Mux25~4_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[28][6]~q ),
	.datac(\registerArray[24][6]~q ),
	.datad(\Mux25~4_combout ),
	.cin(gnd),
	.combout(\Mux25~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~5 .lut_mask = 16'hDDA0;
defparam \Mux25~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y32_N19
dffeas \registerArray[26][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][6] .is_wysiwyg = "true";
defparam \registerArray[26][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N0
cycloneive_lcell_comb \Mux25~2 (
// Equation(s):
// \Mux25~2_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[22][6]~q ))) # (!cuifregS_2 & (\registerArray[18][6]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[18][6]~q ),
	.datac(\registerArray[22][6]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux25~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~2 .lut_mask = 16'hFA44;
defparam \Mux25~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N18
cycloneive_lcell_comb \Mux25~3 (
// Equation(s):
// \Mux25~3_combout  = (cuifregS_3 & ((\Mux25~2_combout  & (\registerArray[30][6]~q )) # (!\Mux25~2_combout  & ((\registerArray[26][6]~q ))))) # (!cuifregS_3 & (((\Mux25~2_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[30][6]~q ),
	.datac(\registerArray[26][6]~q ),
	.datad(\Mux25~2_combout ),
	.cin(gnd),
	.combout(\Mux25~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~3 .lut_mask = 16'hDDA0;
defparam \Mux25~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N2
cycloneive_lcell_comb \Mux25~6 (
// Equation(s):
// \Mux25~6_combout  = (cuifregS_1 & ((cuifregS_0) # ((\Mux25~3_combout )))) # (!cuifregS_1 & (!cuifregS_0 & (\Mux25~5_combout )))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\Mux25~5_combout ),
	.datad(\Mux25~3_combout ),
	.cin(gnd),
	.combout(\Mux25~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~6 .lut_mask = 16'hBA98;
defparam \Mux25~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N8
cycloneive_lcell_comb \Mux25~9 (
// Equation(s):
// \Mux25~9_combout  = (cuifregS_0 & ((\Mux25~6_combout  & ((\Mux25~8_combout ))) # (!\Mux25~6_combout  & (\Mux25~1_combout )))) # (!cuifregS_0 & (((\Mux25~6_combout ))))

	.dataa(\Mux25~1_combout ),
	.datab(cuifregS_0),
	.datac(\Mux25~8_combout ),
	.datad(\Mux25~6_combout ),
	.cin(gnd),
	.combout(\Mux25~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~9 .lut_mask = 16'hF388;
defparam \Mux25~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N26
cycloneive_lcell_comb \Mux25~10 (
// Equation(s):
// \Mux25~10_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & ((\registerArray[5][6]~q ))) # (!cuifregS_0 & (\registerArray[4][6]~q ))))

	.dataa(\registerArray[4][6]~q ),
	.datab(cuifregS_1),
	.datac(\registerArray[5][6]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux25~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~10 .lut_mask = 16'hFC22;
defparam \Mux25~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N20
cycloneive_lcell_comb \Mux25~11 (
// Equation(s):
// \Mux25~11_combout  = (\Mux25~10_combout  & (((\registerArray[7][6]~q ) # (!cuifregS_1)))) # (!\Mux25~10_combout  & (\registerArray[6][6]~q  & ((cuifregS_1))))

	.dataa(\registerArray[6][6]~q ),
	.datab(\registerArray[7][6]~q ),
	.datac(\Mux25~10_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux25~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~11 .lut_mask = 16'hCAF0;
defparam \Mux25~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N18
cycloneive_lcell_comb \Mux25~17 (
// Equation(s):
// \Mux25~17_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & ((\registerArray[13][6]~q ))) # (!cuifregS_0 & (\registerArray[12][6]~q ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[12][6]~q ),
	.datac(\registerArray[13][6]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux25~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~17 .lut_mask = 16'hFA44;
defparam \Mux25~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N8
cycloneive_lcell_comb \Mux25~18 (
// Equation(s):
// \Mux25~18_combout  = (cuifregS_1 & ((\Mux25~17_combout  & ((\registerArray[15][6]~q ))) # (!\Mux25~17_combout  & (\registerArray[14][6]~q )))) # (!cuifregS_1 & (((\Mux25~17_combout ))))

	.dataa(\registerArray[14][6]~q ),
	.datab(\registerArray[15][6]~q ),
	.datac(cuifregS_1),
	.datad(\Mux25~17_combout ),
	.cin(gnd),
	.combout(\Mux25~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~18 .lut_mask = 16'hCFA0;
defparam \Mux25~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N3
dffeas \registerArray[10][6] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux622),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][6] .is_wysiwyg = "true";
defparam \registerArray[10][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N2
cycloneive_lcell_comb \Mux25~12 (
// Equation(s):
// \Mux25~12_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][6]~q ))) # (!cuifregS_1 & (\registerArray[8][6]~q ))))

	.dataa(\registerArray[8][6]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[10][6]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux25~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~12 .lut_mask = 16'hFC22;
defparam \Mux25~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N24
cycloneive_lcell_comb \Mux25~13 (
// Equation(s):
// \Mux25~13_combout  = (cuifregS_0 & ((\Mux25~12_combout  & (\registerArray[11][6]~q )) # (!\Mux25~12_combout  & ((\registerArray[9][6]~q ))))) # (!cuifregS_0 & (((\Mux25~12_combout ))))

	.dataa(\registerArray[11][6]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[9][6]~q ),
	.datad(\Mux25~12_combout ),
	.cin(gnd),
	.combout(\Mux25~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~13 .lut_mask = 16'hBBC0;
defparam \Mux25~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N18
cycloneive_lcell_comb \Mux25~14 (
// Equation(s):
// \Mux25~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][6]~q ))) # (!cuifregS_1 & (\registerArray[1][6]~q ))))

	.dataa(\registerArray[1][6]~q ),
	.datab(\registerArray[3][6]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux25~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~14 .lut_mask = 16'hC0A0;
defparam \Mux25~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N6
cycloneive_lcell_comb \Mux25~15 (
// Equation(s):
// \Mux25~15_combout  = (\Mux25~14_combout ) # ((\registerArray[2][6]~q  & (!cuifregS_0 & cuifregS_1)))

	.dataa(\registerArray[2][6]~q ),
	.datab(cuifregS_0),
	.datac(\Mux25~14_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux25~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~15 .lut_mask = 16'hF2F0;
defparam \Mux25~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N28
cycloneive_lcell_comb \Mux25~16 (
// Equation(s):
// \Mux25~16_combout  = (cuifregS_3 & ((cuifregS_2) # ((\Mux25~13_combout )))) # (!cuifregS_3 & (!cuifregS_2 & ((\Mux25~15_combout ))))

	.dataa(cuifregS_3),
	.datab(cuifregS_2),
	.datac(\Mux25~13_combout ),
	.datad(\Mux25~15_combout ),
	.cin(gnd),
	.combout(\Mux25~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~16 .lut_mask = 16'hB9A8;
defparam \Mux25~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N10
cycloneive_lcell_comb \Mux25~19 (
// Equation(s):
// \Mux25~19_combout  = (cuifregS_2 & ((\Mux25~16_combout  & ((\Mux25~18_combout ))) # (!\Mux25~16_combout  & (\Mux25~11_combout )))) # (!cuifregS_2 & (((\Mux25~16_combout ))))

	.dataa(\Mux25~11_combout ),
	.datab(\Mux25~18_combout ),
	.datac(cuifregS_2),
	.datad(\Mux25~16_combout ),
	.cin(gnd),
	.combout(\Mux25~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~19 .lut_mask = 16'hCFA0;
defparam \Mux25~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N20
cycloneive_lcell_comb \Mux26~7 (
// Equation(s):
// \Mux26~7_combout  = (cuifregS_2 & (((\registerArray[23][5]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[19][5]~q  & ((!cuifregS_3))))

	.dataa(\registerArray[19][5]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[23][5]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux26~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~7 .lut_mask = 16'hCCE2;
defparam \Mux26~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N10
cycloneive_lcell_comb \Mux26~8 (
// Equation(s):
// \Mux26~8_combout  = (cuifregS_3 & ((\Mux26~7_combout  & (\registerArray[31][5]~q )) # (!\Mux26~7_combout  & ((\registerArray[27][5]~q ))))) # (!cuifregS_3 & (((\Mux26~7_combout ))))

	.dataa(\registerArray[31][5]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[27][5]~q ),
	.datad(\Mux26~7_combout ),
	.cin(gnd),
	.combout(\Mux26~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~8 .lut_mask = 16'hBBC0;
defparam \Mux26~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N9
dffeas \registerArray[24][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][5] .is_wysiwyg = "true";
defparam \registerArray[24][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N8
cycloneive_lcell_comb \Mux26~4 (
// Equation(s):
// \Mux26~4_combout  = (cuifregS_3 & (((\registerArray[24][5]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[16][5]~q  & ((!cuifregS_2))))

	.dataa(\registerArray[16][5]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[24][5]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux26~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~4 .lut_mask = 16'hCCE2;
defparam \Mux26~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N10
cycloneive_lcell_comb \Mux26~5 (
// Equation(s):
// \Mux26~5_combout  = (\Mux26~4_combout  & ((\registerArray[28][5]~q ) # ((!cuifregS_2)))) # (!\Mux26~4_combout  & (((\registerArray[20][5]~q  & cuifregS_2))))

	.dataa(\registerArray[28][5]~q ),
	.datab(\Mux26~4_combout ),
	.datac(\registerArray[20][5]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux26~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~5 .lut_mask = 16'hB8CC;
defparam \Mux26~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y32_N15
dffeas \registerArray[22][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][5] .is_wysiwyg = "true";
defparam \registerArray[22][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N29
dffeas \registerArray[26][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][5] .is_wysiwyg = "true";
defparam \registerArray[26][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N28
cycloneive_lcell_comb \Mux26~2 (
// Equation(s):
// \Mux26~2_combout  = (cuifregS_3 & (((\registerArray[26][5]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[18][5]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[18][5]~q ),
	.datac(\registerArray[26][5]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux26~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~2 .lut_mask = 16'hAAE4;
defparam \Mux26~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N14
cycloneive_lcell_comb \Mux26~3 (
// Equation(s):
// \Mux26~3_combout  = (cuifregS_2 & ((\Mux26~2_combout  & (\registerArray[30][5]~q )) # (!\Mux26~2_combout  & ((\registerArray[22][5]~q ))))) # (!cuifregS_2 & (((\Mux26~2_combout ))))

	.dataa(\registerArray[30][5]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[22][5]~q ),
	.datad(\Mux26~2_combout ),
	.cin(gnd),
	.combout(\Mux26~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~3 .lut_mask = 16'hBBC0;
defparam \Mux26~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N26
cycloneive_lcell_comb \Mux26~6 (
// Equation(s):
// \Mux26~6_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\Mux26~3_combout ))) # (!cuifregS_1 & (\Mux26~5_combout ))))

	.dataa(cuifregS_0),
	.datab(\Mux26~5_combout ),
	.datac(cuifregS_1),
	.datad(\Mux26~3_combout ),
	.cin(gnd),
	.combout(\Mux26~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~6 .lut_mask = 16'hF4A4;
defparam \Mux26~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y41_N3
dffeas \registerArray[25][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][5] .is_wysiwyg = "true";
defparam \registerArray[25][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N0
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[21][5]~q ))) # (!cuifregS_2 & (\registerArray[17][5]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[17][5]~q ),
	.datac(\registerArray[21][5]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hFA44;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N2
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// \Mux26~1_combout  = (cuifregS_3 & ((\Mux26~0_combout  & (\registerArray[29][5]~q )) # (!\Mux26~0_combout  & ((\registerArray[25][5]~q ))))) # (!cuifregS_3 & (((\Mux26~0_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[29][5]~q ),
	.datac(\registerArray[25][5]~q ),
	.datad(\Mux26~0_combout ),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hDDA0;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N4
cycloneive_lcell_comb \Mux26~9 (
// Equation(s):
// \Mux26~9_combout  = (cuifregS_0 & ((\Mux26~6_combout  & (\Mux26~8_combout )) # (!\Mux26~6_combout  & ((\Mux26~1_combout ))))) # (!cuifregS_0 & (((\Mux26~6_combout ))))

	.dataa(cuifregS_0),
	.datab(\Mux26~8_combout ),
	.datac(\Mux26~6_combout ),
	.datad(\Mux26~1_combout ),
	.cin(gnd),
	.combout(\Mux26~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~9 .lut_mask = 16'hDAD0;
defparam \Mux26~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N7
dffeas \registerArray[10][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][5] .is_wysiwyg = "true";
defparam \registerArray[10][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N6
cycloneive_lcell_comb \Mux26~10 (
// Equation(s):
// \Mux26~10_combout  = (cuifregS_1 & ((cuifregS_0) # ((\registerArray[10][5]~q )))) # (!cuifregS_1 & (!cuifregS_0 & ((\registerArray[8][5]~q ))))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\registerArray[10][5]~q ),
	.datad(\registerArray[8][5]~q ),
	.cin(gnd),
	.combout(\Mux26~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~10 .lut_mask = 16'hB9A8;
defparam \Mux26~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N4
cycloneive_lcell_comb \Mux26~11 (
// Equation(s):
// \Mux26~11_combout  = (cuifregS_0 & ((\Mux26~10_combout  & (\registerArray[11][5]~q )) # (!\Mux26~10_combout  & ((\registerArray[9][5]~q ))))) # (!cuifregS_0 & (((\Mux26~10_combout ))))

	.dataa(\registerArray[11][5]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[9][5]~q ),
	.datad(\Mux26~10_combout ),
	.cin(gnd),
	.combout(\Mux26~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~11 .lut_mask = 16'hBBC0;
defparam \Mux26~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N26
cycloneive_lcell_comb \registerArray[13][5]~feeder (
// Equation(s):
// \registerArray[13][5]~feeder_combout  = \Mux63~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux632),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[13][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[13][5]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[13][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y44_N27
dffeas \registerArray[13][5] (
	.clk(clk),
	.d(\registerArray[13][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][5] .is_wysiwyg = "true";
defparam \registerArray[13][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N18
cycloneive_lcell_comb \Mux26~17 (
// Equation(s):
// \Mux26~17_combout  = (cuifregS_0 & (((\registerArray[13][5]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[12][5]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[12][5]~q ),
	.datab(\registerArray[13][5]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux26~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~17 .lut_mask = 16'hF0CA;
defparam \Mux26~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N0
cycloneive_lcell_comb \Mux26~18 (
// Equation(s):
// \Mux26~18_combout  = (cuifregS_1 & ((\Mux26~17_combout  & (\registerArray[15][5]~q )) # (!\Mux26~17_combout  & ((\registerArray[14][5]~q ))))) # (!cuifregS_1 & (((\Mux26~17_combout ))))

	.dataa(\registerArray[15][5]~q ),
	.datab(\registerArray[14][5]~q ),
	.datac(cuifregS_1),
	.datad(\Mux26~17_combout ),
	.cin(gnd),
	.combout(\Mux26~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~18 .lut_mask = 16'hAFC0;
defparam \Mux26~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y43_N23
dffeas \registerArray[1][5] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux632),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][5] .is_wysiwyg = "true";
defparam \registerArray[1][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N8
cycloneive_lcell_comb \Mux26~14 (
// Equation(s):
// \Mux26~14_combout  = (cuifregS_0 & ((cuifregS_1 & (\registerArray[3][5]~q )) # (!cuifregS_1 & ((\registerArray[1][5]~q )))))

	.dataa(cuifregS_0),
	.datab(cuifregS_1),
	.datac(\registerArray[3][5]~q ),
	.datad(\registerArray[1][5]~q ),
	.cin(gnd),
	.combout(\Mux26~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~14 .lut_mask = 16'hA280;
defparam \Mux26~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N0
cycloneive_lcell_comb \registerArray[2][5]~feeder (
// Equation(s):
// \registerArray[2][5]~feeder_combout  = \Mux63~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux632),
	.cin(gnd),
	.combout(\registerArray[2][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[2][5]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[2][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y42_N1
dffeas \registerArray[2][5] (
	.clk(clk),
	.d(\registerArray[2][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][5] .is_wysiwyg = "true";
defparam \registerArray[2][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N18
cycloneive_lcell_comb \Mux26~15 (
// Equation(s):
// \Mux26~15_combout  = (\Mux26~14_combout ) # ((!cuifregS_0 & (cuifregS_1 & \registerArray[2][5]~q )))

	.dataa(cuifregS_0),
	.datab(cuifregS_1),
	.datac(\Mux26~14_combout ),
	.datad(\registerArray[2][5]~q ),
	.cin(gnd),
	.combout(\Mux26~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~15 .lut_mask = 16'hF4F0;
defparam \Mux26~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N28
cycloneive_lcell_comb \Mux26~16 (
// Equation(s):
// \Mux26~16_combout  = (cuifregS_2 & ((\Mux26~13_combout ) # ((cuifregS_3)))) # (!cuifregS_2 & (((!cuifregS_3 & \Mux26~15_combout ))))

	.dataa(\Mux26~13_combout ),
	.datab(cuifregS_2),
	.datac(cuifregS_3),
	.datad(\Mux26~15_combout ),
	.cin(gnd),
	.combout(\Mux26~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~16 .lut_mask = 16'hCBC8;
defparam \Mux26~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N2
cycloneive_lcell_comb \Mux26~19 (
// Equation(s):
// \Mux26~19_combout  = (cuifregS_3 & ((\Mux26~16_combout  & ((\Mux26~18_combout ))) # (!\Mux26~16_combout  & (\Mux26~11_combout )))) # (!cuifregS_3 & (((\Mux26~16_combout ))))

	.dataa(cuifregS_3),
	.datab(\Mux26~11_combout ),
	.datac(\Mux26~18_combout ),
	.datad(\Mux26~16_combout ),
	.cin(gnd),
	.combout(\Mux26~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~19 .lut_mask = 16'hF588;
defparam \Mux26~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y34_N31
dffeas \registerArray[28][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][3] .is_wysiwyg = "true";
defparam \registerArray[28][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N24
cycloneive_lcell_comb \Mux60~4 (
// Equation(s):
// \Mux60~4_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[20][3]~q )) # (!cuifregT_2 & ((\registerArray[16][3]~q )))))

	.dataa(cuifregT_3),
	.datab(\registerArray[20][3]~q ),
	.datac(\registerArray[16][3]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux60~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~4 .lut_mask = 16'hEE50;
defparam \Mux60~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N30
cycloneive_lcell_comb \Mux60~5 (
// Equation(s):
// \Mux60~5_combout  = (cuifregT_3 & ((\Mux60~4_combout  & ((\registerArray[28][3]~q ))) # (!\Mux60~4_combout  & (\registerArray[24][3]~q )))) # (!cuifregT_3 & (((\Mux60~4_combout ))))

	.dataa(cuifregT_3),
	.datab(\registerArray[24][3]~q ),
	.datac(\registerArray[28][3]~q ),
	.datad(\Mux60~4_combout ),
	.cin(gnd),
	.combout(\Mux60~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~5 .lut_mask = 16'hF588;
defparam \Mux60~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y31_N15
dffeas \registerArray[18][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~64_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[18][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[18][3] .is_wysiwyg = "true";
defparam \registerArray[18][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N14
cycloneive_lcell_comb \Mux60~2 (
// Equation(s):
// \Mux60~2_combout  = (cuifregT_2 & ((\registerArray[22][3]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[18][3]~q  & !cuifregT_3))))

	.dataa(\registerArray[22][3]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[18][3]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux60~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~2 .lut_mask = 16'hCCB8;
defparam \Mux60~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N8
cycloneive_lcell_comb \Mux60~3 (
// Equation(s):
// \Mux60~3_combout  = (\Mux60~2_combout  & (((\registerArray[30][3]~q ) # (!cuifregT_3)))) # (!\Mux60~2_combout  & (\registerArray[26][3]~q  & ((cuifregT_3))))

	.dataa(\registerArray[26][3]~q ),
	.datab(\Mux60~2_combout ),
	.datac(\registerArray[30][3]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux60~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~3 .lut_mask = 16'hE2CC;
defparam \Mux60~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N8
cycloneive_lcell_comb \Mux60~6 (
// Equation(s):
// \Mux60~6_combout  = (cuifregT_1 & (((cuifregT_01) # (\Mux60~3_combout )))) # (!cuifregT_1 & (\Mux60~5_combout  & (!cuifregT_01)))

	.dataa(\Mux60~5_combout ),
	.datab(cuifregT_1),
	.datac(cuifregT_0),
	.datad(\Mux60~3_combout ),
	.cin(gnd),
	.combout(\Mux60~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~6 .lut_mask = 16'hCEC2;
defparam \Mux60~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N0
cycloneive_lcell_comb \registerArray[25][3]~feeder (
// Equation(s):
// \registerArray[25][3]~feeder_combout  = \Mux65~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux65),
	.cin(gnd),
	.combout(\registerArray[25][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[25][3]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[25][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N1
dffeas \registerArray[25][3] (
	.clk(clk),
	.d(\registerArray[25][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][3] .is_wysiwyg = "true";
defparam \registerArray[25][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N6
cycloneive_lcell_comb \Mux60~0 (
// Equation(s):
// \Mux60~0_combout  = (cuifregT_3 & (((\registerArray[25][3]~q ) # (cuifregT_2)))) # (!cuifregT_3 & (\registerArray[17][3]~q  & ((!cuifregT_2))))

	.dataa(\registerArray[17][3]~q ),
	.datab(\registerArray[25][3]~q ),
	.datac(cuifregT_3),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux60~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~0 .lut_mask = 16'hF0CA;
defparam \Mux60~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N2
cycloneive_lcell_comb \Mux60~1 (
// Equation(s):
// \Mux60~1_combout  = (cuifregT_2 & ((\Mux60~0_combout  & ((\registerArray[29][3]~q ))) # (!\Mux60~0_combout  & (\registerArray[21][3]~q )))) # (!cuifregT_2 & (((\Mux60~0_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[21][3]~q ),
	.datac(\registerArray[29][3]~q ),
	.datad(\Mux60~0_combout ),
	.cin(gnd),
	.combout(\Mux60~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~1 .lut_mask = 16'hF588;
defparam \Mux60~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N9
dffeas \registerArray[19][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~70_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[19][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[19][3] .is_wysiwyg = "true";
defparam \registerArray[19][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N8
cycloneive_lcell_comb \Mux60~7 (
// Equation(s):
// \Mux60~7_combout  = (cuifregT_3 & ((\registerArray[27][3]~q ) # ((cuifregT_2)))) # (!cuifregT_3 & (((\registerArray[19][3]~q  & !cuifregT_2))))

	.dataa(\registerArray[27][3]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[19][3]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux60~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~7 .lut_mask = 16'hCCB8;
defparam \Mux60~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y39_N19
dffeas \registerArray[31][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][3] .is_wysiwyg = "true";
defparam \registerArray[31][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y39_N18
cycloneive_lcell_comb \Mux60~8 (
// Equation(s):
// \Mux60~8_combout  = (\Mux60~7_combout  & (((\registerArray[31][3]~q ) # (!cuifregT_2)))) # (!\Mux60~7_combout  & (\registerArray[23][3]~q  & ((cuifregT_2))))

	.dataa(\registerArray[23][3]~q ),
	.datab(\Mux60~7_combout ),
	.datac(\registerArray[31][3]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux60~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~8 .lut_mask = 16'hE2CC;
defparam \Mux60~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N5
dffeas \registerArray[14][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][3] .is_wysiwyg = "true";
defparam \registerArray[14][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N0
cycloneive_lcell_comb \registerArray[12][3]~feeder (
// Equation(s):
// \registerArray[12][3]~feeder_combout  = \Mux65~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux65),
	.cin(gnd),
	.combout(\registerArray[12][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[12][3]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[12][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y30_N1
dffeas \registerArray[12][3] (
	.clk(clk),
	.d(\registerArray[12][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][3] .is_wysiwyg = "true";
defparam \registerArray[12][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N6
cycloneive_lcell_comb \Mux60~17 (
// Equation(s):
// \Mux60~17_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & ((\registerArray[13][3]~q ))) # (!cuifregT_01 & (\registerArray[12][3]~q ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[12][3]~q ),
	.datac(\registerArray[13][3]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux60~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~17 .lut_mask = 16'hFA44;
defparam \Mux60~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N4
cycloneive_lcell_comb \Mux60~18 (
// Equation(s):
// \Mux60~18_combout  = (cuifregT_1 & ((\Mux60~17_combout  & (\registerArray[15][3]~q )) # (!\Mux60~17_combout  & ((\registerArray[14][3]~q ))))) # (!cuifregT_1 & (((\Mux60~17_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[15][3]~q ),
	.datac(\registerArray[14][3]~q ),
	.datad(\Mux60~17_combout ),
	.cin(gnd),
	.combout(\Mux60~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~18 .lut_mask = 16'hDDA0;
defparam \Mux60~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N5
dffeas \registerArray[5][3] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux65),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][3] .is_wysiwyg = "true";
defparam \registerArray[5][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N4
cycloneive_lcell_comb \Mux60~10 (
// Equation(s):
// \Mux60~10_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & ((\registerArray[5][3]~q ))) # (!cuifregT_01 & (\registerArray[4][3]~q ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[4][3]~q ),
	.datac(\registerArray[5][3]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux60~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~10 .lut_mask = 16'hFA44;
defparam \Mux60~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N8
cycloneive_lcell_comb \Mux60~11 (
// Equation(s):
// \Mux60~11_combout  = (cuifregT_1 & ((\Mux60~10_combout  & (\registerArray[7][3]~q )) # (!\Mux60~10_combout  & ((\registerArray[6][3]~q ))))) # (!cuifregT_1 & (((\Mux60~10_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[7][3]~q ),
	.datac(\registerArray[6][3]~q ),
	.datad(\Mux60~10_combout ),
	.cin(gnd),
	.combout(\Mux60~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~11 .lut_mask = 16'hDDA0;
defparam \Mux60~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N26
cycloneive_lcell_comb \registerArray[2][3]~feeder (
// Equation(s):
// \registerArray[2][3]~feeder_combout  = \Mux65~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux65),
	.cin(gnd),
	.combout(\registerArray[2][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[2][3]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[2][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y44_N27
dffeas \registerArray[2][3] (
	.clk(clk),
	.d(\registerArray[2][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~80_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[2][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[2][3] .is_wysiwyg = "true";
defparam \registerArray[2][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N30
cycloneive_lcell_comb \Mux60~14 (
// Equation(s):
// \Mux60~14_combout  = (cuifregT_01 & ((cuifregT_1 & ((\registerArray[3][3]~q ))) # (!cuifregT_1 & (\registerArray[1][3]~q ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[1][3]~q ),
	.datac(\registerArray[3][3]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux60~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~14 .lut_mask = 16'hE400;
defparam \Mux60~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N14
cycloneive_lcell_comb \Mux60~15 (
// Equation(s):
// \Mux60~15_combout  = (\Mux60~14_combout ) # ((!cuifregT_01 & (cuifregT_1 & \registerArray[2][3]~q )))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\registerArray[2][3]~q ),
	.datad(\Mux60~14_combout ),
	.cin(gnd),
	.combout(\Mux60~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~15 .lut_mask = 16'hFF40;
defparam \Mux60~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N10
cycloneive_lcell_comb \registerArray[11][3]~feeder (
// Equation(s):
// \registerArray[11][3]~feeder_combout  = \Mux65~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux65),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[11][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[11][3]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[11][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N11
dffeas \registerArray[11][3] (
	.clk(clk),
	.d(\registerArray[11][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][3] .is_wysiwyg = "true";
defparam \registerArray[11][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N14
cycloneive_lcell_comb \Mux60~12 (
// Equation(s):
// \Mux60~12_combout  = (cuifregT_01 & (((cuifregT_1)))) # (!cuifregT_01 & ((cuifregT_1 & ((\registerArray[10][3]~q ))) # (!cuifregT_1 & (\registerArray[8][3]~q ))))

	.dataa(\registerArray[8][3]~q ),
	.datab(cuifregT_0),
	.datac(\registerArray[10][3]~q ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux60~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~12 .lut_mask = 16'hFC22;
defparam \Mux60~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N16
cycloneive_lcell_comb \Mux60~13 (
// Equation(s):
// \Mux60~13_combout  = (\Mux60~12_combout  & (((\registerArray[11][3]~q ) # (!cuifregT_01)))) # (!\Mux60~12_combout  & (\registerArray[9][3]~q  & ((cuifregT_01))))

	.dataa(\registerArray[9][3]~q ),
	.datab(\registerArray[11][3]~q ),
	.datac(\Mux60~12_combout ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux60~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~13 .lut_mask = 16'hCAF0;
defparam \Mux60~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y34_N12
cycloneive_lcell_comb \Mux60~16 (
// Equation(s):
// \Mux60~16_combout  = (cuifregT_3 & ((cuifregT_2) # ((\Mux60~13_combout )))) # (!cuifregT_3 & (!cuifregT_2 & (\Mux60~15_combout )))

	.dataa(cuifregT_3),
	.datab(cuifregT_2),
	.datac(\Mux60~15_combout ),
	.datad(\Mux60~13_combout ),
	.cin(gnd),
	.combout(\Mux60~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~16 .lut_mask = 16'hBA98;
defparam \Mux60~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y37_N10
cycloneive_lcell_comb \registerArray[7][16]~feeder (
// Equation(s):
// \registerArray[7][16]~feeder_combout  = \Mux52~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux522),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[7][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[7][16]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[7][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y37_N11
dffeas \registerArray[7][16] (
	.clk(clk),
	.d(\registerArray[7][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][16] .is_wysiwyg = "true";
defparam \registerArray[7][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N20
cycloneive_lcell_comb \Mux15~10 (
// Equation(s):
// \Mux15~10_combout  = (cuifregS_0 & ((\registerArray[5][16]~q ) # ((cuifregS_1)))) # (!cuifregS_0 & (((\registerArray[4][16]~q  & !cuifregS_1))))

	.dataa(\registerArray[5][16]~q ),
	.datab(\registerArray[4][16]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux15~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~10 .lut_mask = 16'hF0AC;
defparam \Mux15~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N16
cycloneive_lcell_comb \Mux15~11 (
// Equation(s):
// \Mux15~11_combout  = (cuifregS_1 & ((\Mux15~10_combout  & (\registerArray[7][16]~q )) # (!\Mux15~10_combout  & ((\registerArray[6][16]~q ))))) # (!cuifregS_1 & (((\Mux15~10_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[7][16]~q ),
	.datac(\registerArray[6][16]~q ),
	.datad(\Mux15~10_combout ),
	.cin(gnd),
	.combout(\Mux15~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~11 .lut_mask = 16'hDDA0;
defparam \Mux15~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N0
cycloneive_lcell_comb \Mux15~14 (
// Equation(s):
// \Mux15~14_combout  = (cuifregS_0 & ((cuifregS_1 & (\registerArray[3][16]~q )) # (!cuifregS_1 & ((\registerArray[1][16]~q )))))

	.dataa(\registerArray[3][16]~q ),
	.datab(\registerArray[1][16]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux15~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~14 .lut_mask = 16'hA0C0;
defparam \Mux15~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N26
cycloneive_lcell_comb \Mux15~15 (
// Equation(s):
// \Mux15~15_combout  = (\Mux15~14_combout ) # ((\registerArray[2][16]~q  & (!cuifregS_0 & cuifregS_1)))

	.dataa(\registerArray[2][16]~q ),
	.datab(cuifregS_0),
	.datac(cuifregS_1),
	.datad(\Mux15~14_combout ),
	.cin(gnd),
	.combout(\Mux15~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~15 .lut_mask = 16'hFF20;
defparam \Mux15~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N11
dffeas \registerArray[10][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][16] .is_wysiwyg = "true";
defparam \registerArray[10][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N10
cycloneive_lcell_comb \Mux15~12 (
// Equation(s):
// \Mux15~12_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][16]~q ))) # (!cuifregS_1 & (\registerArray[8][16]~q ))))

	.dataa(\registerArray[8][16]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[10][16]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux15~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~12 .lut_mask = 16'hFC22;
defparam \Mux15~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N0
cycloneive_lcell_comb \Mux15~13 (
// Equation(s):
// \Mux15~13_combout  = (cuifregS_0 & ((\Mux15~12_combout  & (\registerArray[11][16]~q )) # (!\Mux15~12_combout  & ((\registerArray[9][16]~q ))))) # (!cuifregS_0 & (((\Mux15~12_combout ))))

	.dataa(\registerArray[11][16]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[9][16]~q ),
	.datad(\Mux15~12_combout ),
	.cin(gnd),
	.combout(\Mux15~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~13 .lut_mask = 16'hBBC0;
defparam \Mux15~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N8
cycloneive_lcell_comb \Mux15~16 (
// Equation(s):
// \Mux15~16_combout  = (cuifregS_3 & ((cuifregS_2) # ((\Mux15~13_combout )))) # (!cuifregS_3 & (!cuifregS_2 & (\Mux15~15_combout )))

	.dataa(cuifregS_3),
	.datab(cuifregS_2),
	.datac(\Mux15~15_combout ),
	.datad(\Mux15~13_combout ),
	.cin(gnd),
	.combout(\Mux15~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~16 .lut_mask = 16'hBA98;
defparam \Mux15~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N20
cycloneive_lcell_comb \registerArray[13][16]~feeder (
// Equation(s):
// \registerArray[13][16]~feeder_combout  = \Mux52~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux522),
	.cin(gnd),
	.combout(\registerArray[13][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[13][16]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[13][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y37_N21
dffeas \registerArray[13][16] (
	.clk(clk),
	.d(\registerArray[13][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][16] .is_wysiwyg = "true";
defparam \registerArray[13][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N28
cycloneive_lcell_comb \Mux15~17 (
// Equation(s):
// \Mux15~17_combout  = (cuifregS_0 & (((\registerArray[13][16]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[12][16]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[12][16]~q ),
	.datab(\registerArray[13][16]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux15~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~17 .lut_mask = 16'hF0CA;
defparam \Mux15~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y40_N18
cycloneive_lcell_comb \Mux15~18 (
// Equation(s):
// \Mux15~18_combout  = (cuifregS_1 & ((\Mux15~17_combout  & (\registerArray[15][16]~q )) # (!\Mux15~17_combout  & ((\registerArray[14][16]~q ))))) # (!cuifregS_1 & (((\Mux15~17_combout ))))

	.dataa(\registerArray[15][16]~q ),
	.datab(\registerArray[14][16]~q ),
	.datac(cuifregS_1),
	.datad(\Mux15~17_combout ),
	.cin(gnd),
	.combout(\Mux15~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~18 .lut_mask = 16'hAFC0;
defparam \Mux15~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N14
cycloneive_lcell_comb \Mux15~19 (
// Equation(s):
// \Mux15~19_combout  = (cuifregS_2 & ((\Mux15~16_combout  & ((\Mux15~18_combout ))) # (!\Mux15~16_combout  & (\Mux15~11_combout )))) # (!cuifregS_2 & (((\Mux15~16_combout ))))

	.dataa(\Mux15~11_combout ),
	.datab(cuifregS_2),
	.datac(\Mux15~16_combout ),
	.datad(\Mux15~18_combout ),
	.cin(gnd),
	.combout(\Mux15~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~19 .lut_mask = 16'hF838;
defparam \Mux15~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N21
dffeas \registerArray[22][16] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux522),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][16] .is_wysiwyg = "true";
defparam \registerArray[22][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N20
cycloneive_lcell_comb \Mux15~2 (
// Equation(s):
// \Mux15~2_combout  = (cuifregS_2 & (((\registerArray[22][16]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[18][16]~q  & ((!cuifregS_3))))

	.dataa(\registerArray[18][16]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[22][16]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux15~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~2 .lut_mask = 16'hCCE2;
defparam \Mux15~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N2
cycloneive_lcell_comb \Mux15~3 (
// Equation(s):
// \Mux15~3_combout  = (cuifregS_3 & ((\Mux15~2_combout  & (\registerArray[30][16]~q )) # (!\Mux15~2_combout  & ((\registerArray[26][16]~q ))))) # (!cuifregS_3 & (((\Mux15~2_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[30][16]~q ),
	.datac(\registerArray[26][16]~q ),
	.datad(\Mux15~2_combout ),
	.cin(gnd),
	.combout(\Mux15~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~3 .lut_mask = 16'hDDA0;
defparam \Mux15~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N10
cycloneive_lcell_comb \Mux15~6 (
// Equation(s):
// \Mux15~6_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\Mux15~3_combout ))) # (!cuifregS_1 & (\Mux15~5_combout ))))

	.dataa(\Mux15~5_combout ),
	.datab(cuifregS_0),
	.datac(cuifregS_1),
	.datad(\Mux15~3_combout ),
	.cin(gnd),
	.combout(\Mux15~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~6 .lut_mask = 16'hF2C2;
defparam \Mux15~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N2
cycloneive_lcell_comb \Mux15~7 (
// Equation(s):
// \Mux15~7_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & ((\registerArray[27][16]~q ))) # (!cuifregS_3 & (\registerArray[19][16]~q ))))

	.dataa(\registerArray[19][16]~q ),
	.datab(\registerArray[27][16]~q ),
	.datac(cuifregS_2),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux15~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~7 .lut_mask = 16'hFC0A;
defparam \Mux15~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y40_N0
cycloneive_lcell_comb \Mux15~8 (
// Equation(s):
// \Mux15~8_combout  = (cuifregS_2 & ((\Mux15~7_combout  & ((\registerArray[31][16]~q ))) # (!\Mux15~7_combout  & (\registerArray[23][16]~q )))) # (!cuifregS_2 & (((\Mux15~7_combout ))))

	.dataa(\registerArray[23][16]~q ),
	.datab(\registerArray[31][16]~q ),
	.datac(cuifregS_2),
	.datad(\Mux15~7_combout ),
	.cin(gnd),
	.combout(\Mux15~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~8 .lut_mask = 16'hCFA0;
defparam \Mux15~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N14
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// \Mux15~0_combout  = (cuifregS_3 & (((\registerArray[25][16]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[17][16]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[17][16]~q ),
	.datac(\registerArray[25][16]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hAAE4;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N0
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// \Mux15~1_combout  = (cuifregS_2 & ((\Mux15~0_combout  & ((\registerArray[29][16]~q ))) # (!\Mux15~0_combout  & (\registerArray[21][16]~q )))) # (!cuifregS_2 & (((\Mux15~0_combout ))))

	.dataa(\registerArray[21][16]~q ),
	.datab(cuifregS_2),
	.datac(\Mux15~0_combout ),
	.datad(\registerArray[29][16]~q ),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'hF838;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N24
cycloneive_lcell_comb \Mux15~9 (
// Equation(s):
// \Mux15~9_combout  = (\Mux15~6_combout  & (((\Mux15~8_combout )) # (!cuifregS_0))) # (!\Mux15~6_combout  & (cuifregS_0 & ((\Mux15~1_combout ))))

	.dataa(\Mux15~6_combout ),
	.datab(cuifregS_0),
	.datac(\Mux15~8_combout ),
	.datad(\Mux15~1_combout ),
	.cin(gnd),
	.combout(\Mux15~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~9 .lut_mask = 16'hE6A2;
defparam \Mux15~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N16
cycloneive_lcell_comb \Mux16~2 (
// Equation(s):
// \Mux16~2_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & (\registerArray[26][15]~q )) # (!cuifregS_3 & ((\registerArray[18][15]~q )))))

	.dataa(\registerArray[26][15]~q ),
	.datab(\registerArray[18][15]~q ),
	.datac(cuifregS_2),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux16~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~2 .lut_mask = 16'hFA0C;
defparam \Mux16~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N30
cycloneive_lcell_comb \Mux16~3 (
// Equation(s):
// \Mux16~3_combout  = (cuifregS_2 & ((\Mux16~2_combout  & (\registerArray[30][15]~q )) # (!\Mux16~2_combout  & ((\registerArray[22][15]~q ))))) # (!cuifregS_2 & (((\Mux16~2_combout ))))

	.dataa(\registerArray[30][15]~q ),
	.datab(\registerArray[22][15]~q ),
	.datac(cuifregS_2),
	.datad(\Mux16~2_combout ),
	.cin(gnd),
	.combout(\Mux16~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~3 .lut_mask = 16'hAFC0;
defparam \Mux16~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N3
dffeas \registerArray[20][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][15] .is_wysiwyg = "true";
defparam \registerArray[20][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y43_N1
dffeas \registerArray[24][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][15] .is_wysiwyg = "true";
defparam \registerArray[24][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N0
cycloneive_lcell_comb \Mux16~4 (
// Equation(s):
// \Mux16~4_combout  = (cuifregS_3 & (((\registerArray[24][15]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[16][15]~q  & ((!cuifregS_2))))

	.dataa(\registerArray[16][15]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[24][15]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux16~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~4 .lut_mask = 16'hCCE2;
defparam \Mux16~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N2
cycloneive_lcell_comb \Mux16~5 (
// Equation(s):
// \Mux16~5_combout  = (cuifregS_2 & ((\Mux16~4_combout  & (\registerArray[28][15]~q )) # (!\Mux16~4_combout  & ((\registerArray[20][15]~q ))))) # (!cuifregS_2 & (((\Mux16~4_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[28][15]~q ),
	.datac(\registerArray[20][15]~q ),
	.datad(\Mux16~4_combout ),
	.cin(gnd),
	.combout(\Mux16~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~5 .lut_mask = 16'hDDA0;
defparam \Mux16~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N24
cycloneive_lcell_comb \Mux16~6 (
// Equation(s):
// \Mux16~6_combout  = (cuifregS_0 & (cuifregS_1)) # (!cuifregS_0 & ((cuifregS_1 & (\Mux16~3_combout )) # (!cuifregS_1 & ((\Mux16~5_combout )))))

	.dataa(cuifregS_0),
	.datab(cuifregS_1),
	.datac(\Mux16~3_combout ),
	.datad(\Mux16~5_combout ),
	.cin(gnd),
	.combout(\Mux16~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~6 .lut_mask = 16'hD9C8;
defparam \Mux16~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N18
cycloneive_lcell_comb \Mux16~7 (
// Equation(s):
// \Mux16~7_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[23][15]~q ))) # (!cuifregS_2 & (\registerArray[19][15]~q ))))

	.dataa(\registerArray[19][15]~q ),
	.datab(\registerArray[23][15]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux16~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~7 .lut_mask = 16'hFC0A;
defparam \Mux16~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N24
cycloneive_lcell_comb \Mux16~8 (
// Equation(s):
// \Mux16~8_combout  = (cuifregS_3 & ((\Mux16~7_combout  & ((\registerArray[31][15]~q ))) # (!\Mux16~7_combout  & (\registerArray[27][15]~q )))) # (!cuifregS_3 & (((\Mux16~7_combout ))))

	.dataa(\registerArray[27][15]~q ),
	.datab(\registerArray[31][15]~q ),
	.datac(cuifregS_3),
	.datad(\Mux16~7_combout ),
	.cin(gnd),
	.combout(\Mux16~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~8 .lut_mask = 16'hCFA0;
defparam \Mux16~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y30_N3
dffeas \registerArray[25][15] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux532),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][15] .is_wysiwyg = "true";
defparam \registerArray[25][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N20
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// \Mux16~0_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[21][15]~q ))) # (!cuifregS_2 & (\registerArray[17][15]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[17][15]~q ),
	.datac(\registerArray[21][15]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'hFA44;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N2
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// \Mux16~1_combout  = (cuifregS_3 & ((\Mux16~0_combout  & (\registerArray[29][15]~q )) # (!\Mux16~0_combout  & ((\registerArray[25][15]~q ))))) # (!cuifregS_3 & (((\Mux16~0_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[29][15]~q ),
	.datac(\registerArray[25][15]~q ),
	.datad(\Mux16~0_combout ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hDDA0;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N14
cycloneive_lcell_comb \Mux16~9 (
// Equation(s):
// \Mux16~9_combout  = (\Mux16~6_combout  & (((\Mux16~8_combout )) # (!cuifregS_0))) # (!\Mux16~6_combout  & (cuifregS_0 & ((\Mux16~1_combout ))))

	.dataa(\Mux16~6_combout ),
	.datab(cuifregS_0),
	.datac(\Mux16~8_combout ),
	.datad(\Mux16~1_combout ),
	.cin(gnd),
	.combout(\Mux16~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~9 .lut_mask = 16'hE6A2;
defparam \Mux16~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N16
cycloneive_lcell_comb \registerArray[5][15]~feeder (
// Equation(s):
// \registerArray[5][15]~feeder_combout  = \Mux53~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux532),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[5][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[5][15]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[5][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y31_N17
dffeas \registerArray[5][15] (
	.clk(clk),
	.d(\registerArray[5][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][15] .is_wysiwyg = "true";
defparam \registerArray[5][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N22
cycloneive_lcell_comb \Mux16~12 (
// Equation(s):
// \Mux16~12_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & (\registerArray[5][15]~q )) # (!cuifregS_0 & ((\registerArray[4][15]~q )))))

	.dataa(cuifregS_1),
	.datab(\registerArray[5][15]~q ),
	.datac(cuifregS_0),
	.datad(\registerArray[4][15]~q ),
	.cin(gnd),
	.combout(\Mux16~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~12 .lut_mask = 16'hE5E0;
defparam \Mux16~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N12
cycloneive_lcell_comb \Mux16~13 (
// Equation(s):
// \Mux16~13_combout  = (\Mux16~12_combout  & ((\registerArray[7][15]~q ) # ((!cuifregS_1)))) # (!\Mux16~12_combout  & (((\registerArray[6][15]~q  & cuifregS_1))))

	.dataa(\registerArray[7][15]~q ),
	.datab(\registerArray[6][15]~q ),
	.datac(\Mux16~12_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux16~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~13 .lut_mask = 16'hACF0;
defparam \Mux16~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N22
cycloneive_lcell_comb \Mux16~16 (
// Equation(s):
// \Mux16~16_combout  = (cuifregS_2 & (((cuifregS_3) # (\Mux16~13_combout )))) # (!cuifregS_2 & (\Mux16~15_combout  & (!cuifregS_3)))

	.dataa(\Mux16~15_combout ),
	.datab(cuifregS_2),
	.datac(cuifregS_3),
	.datad(\Mux16~13_combout ),
	.cin(gnd),
	.combout(\Mux16~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~16 .lut_mask = 16'hCEC2;
defparam \Mux16~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N28
cycloneive_lcell_comb \registerArray[13][15]~feeder (
// Equation(s):
// \registerArray[13][15]~feeder_combout  = \Mux53~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux532),
	.cin(gnd),
	.combout(\registerArray[13][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[13][15]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[13][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N29
dffeas \registerArray[13][15] (
	.clk(clk),
	.d(\registerArray[13][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][15] .is_wysiwyg = "true";
defparam \registerArray[13][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N0
cycloneive_lcell_comb \Mux16~17 (
// Equation(s):
// \Mux16~17_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & (\registerArray[13][15]~q )) # (!cuifregS_0 & ((\registerArray[12][15]~q )))))

	.dataa(cuifregS_1),
	.datab(\registerArray[13][15]~q ),
	.datac(\registerArray[12][15]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux16~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~17 .lut_mask = 16'hEE50;
defparam \Mux16~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N26
cycloneive_lcell_comb \Mux16~18 (
// Equation(s):
// \Mux16~18_combout  = (cuifregS_1 & ((\Mux16~17_combout  & (\registerArray[15][15]~q )) # (!\Mux16~17_combout  & ((\registerArray[14][15]~q ))))) # (!cuifregS_1 & (((\Mux16~17_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[15][15]~q ),
	.datac(\registerArray[14][15]~q ),
	.datad(\Mux16~17_combout ),
	.cin(gnd),
	.combout(\Mux16~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~18 .lut_mask = 16'hDDA0;
defparam \Mux16~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N10
cycloneive_lcell_comb \Mux16~10 (
// Equation(s):
// \Mux16~10_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\registerArray[10][15]~q )) # (!cuifregS_1 & ((\registerArray[8][15]~q )))))

	.dataa(\registerArray[10][15]~q ),
	.datab(\registerArray[8][15]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux16~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~10 .lut_mask = 16'hFA0C;
defparam \Mux16~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y37_N18
cycloneive_lcell_comb \Mux16~11 (
// Equation(s):
// \Mux16~11_combout  = (\Mux16~10_combout  & (((\registerArray[11][15]~q ) # (!cuifregS_0)))) # (!\Mux16~10_combout  & (\registerArray[9][15]~q  & ((cuifregS_0))))

	.dataa(\registerArray[9][15]~q ),
	.datab(\registerArray[11][15]~q ),
	.datac(\Mux16~10_combout ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux16~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~11 .lut_mask = 16'hCAF0;
defparam \Mux16~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N16
cycloneive_lcell_comb \Mux16~19 (
// Equation(s):
// \Mux16~19_combout  = (\Mux16~16_combout  & (((\Mux16~18_combout )) # (!cuifregS_3))) # (!\Mux16~16_combout  & (cuifregS_3 & ((\Mux16~11_combout ))))

	.dataa(\Mux16~16_combout ),
	.datab(cuifregS_3),
	.datac(\Mux16~18_combout ),
	.datad(\Mux16~11_combout ),
	.cin(gnd),
	.combout(\Mux16~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~19 .lut_mask = 16'hE6A2;
defparam \Mux16~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N26
cycloneive_lcell_comb \Mux17~14 (
// Equation(s):
// \Mux17~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][14]~q ))) # (!cuifregS_1 & (\registerArray[1][14]~q ))))

	.dataa(\registerArray[1][14]~q ),
	.datab(\registerArray[3][14]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux17~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~14 .lut_mask = 16'hC0A0;
defparam \Mux17~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N4
cycloneive_lcell_comb \Mux17~15 (
// Equation(s):
// \Mux17~15_combout  = (\Mux17~14_combout ) # ((\registerArray[2][14]~q  & (cuifregS_1 & !cuifregS_0)))

	.dataa(\registerArray[2][14]~q ),
	.datab(\Mux17~14_combout ),
	.datac(cuifregS_1),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux17~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~15 .lut_mask = 16'hCCEC;
defparam \Mux17~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N28
cycloneive_lcell_comb \Mux17~13 (
// Equation(s):
// \Mux17~13_combout  = (\Mux17~12_combout  & (((\registerArray[11][14]~q )) # (!cuifregS_0))) # (!\Mux17~12_combout  & (cuifregS_0 & (\registerArray[9][14]~q )))

	.dataa(\Mux17~12_combout ),
	.datab(cuifregS_0),
	.datac(\registerArray[9][14]~q ),
	.datad(\registerArray[11][14]~q ),
	.cin(gnd),
	.combout(\Mux17~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~13 .lut_mask = 16'hEA62;
defparam \Mux17~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N18
cycloneive_lcell_comb \Mux17~16 (
// Equation(s):
// \Mux17~16_combout  = (cuifregS_2 & (cuifregS_3)) # (!cuifregS_2 & ((cuifregS_3 & ((\Mux17~13_combout ))) # (!cuifregS_3 & (\Mux17~15_combout ))))

	.dataa(cuifregS_2),
	.datab(cuifregS_3),
	.datac(\Mux17~15_combout ),
	.datad(\Mux17~13_combout ),
	.cin(gnd),
	.combout(\Mux17~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~16 .lut_mask = 16'hDC98;
defparam \Mux17~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y39_N17
dffeas \registerArray[13][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][14] .is_wysiwyg = "true";
defparam \registerArray[13][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N16
cycloneive_lcell_comb \Mux17~17 (
// Equation(s):
// \Mux17~17_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & ((\registerArray[13][14]~q ))) # (!cuifregS_0 & (\registerArray[12][14]~q ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[12][14]~q ),
	.datac(\registerArray[13][14]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux17~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~17 .lut_mask = 16'hFA44;
defparam \Mux17~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N4
cycloneive_lcell_comb \Mux17~18 (
// Equation(s):
// \Mux17~18_combout  = (cuifregS_1 & ((\Mux17~17_combout  & (\registerArray[15][14]~q )) # (!\Mux17~17_combout  & ((\registerArray[14][14]~q ))))) # (!cuifregS_1 & (((\Mux17~17_combout ))))

	.dataa(\registerArray[15][14]~q ),
	.datab(\registerArray[14][14]~q ),
	.datac(cuifregS_1),
	.datad(\Mux17~17_combout ),
	.cin(gnd),
	.combout(\Mux17~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~18 .lut_mask = 16'hAFC0;
defparam \Mux17~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N8
cycloneive_lcell_comb \registerArray[6][14]~feeder (
// Equation(s):
// \registerArray[6][14]~feeder_combout  = \Mux54~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux542),
	.cin(gnd),
	.combout(\registerArray[6][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[6][14]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[6][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N9
dffeas \registerArray[6][14] (
	.clk(clk),
	.d(\registerArray[6][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][14] .is_wysiwyg = "true";
defparam \registerArray[6][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N30
cycloneive_lcell_comb \Mux17~10 (
// Equation(s):
// \Mux17~10_combout  = (cuifregS_0 & ((\registerArray[5][14]~q ) # ((cuifregS_1)))) # (!cuifregS_0 & (((\registerArray[4][14]~q  & !cuifregS_1))))

	.dataa(\registerArray[5][14]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[4][14]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux17~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~10 .lut_mask = 16'hCCB8;
defparam \Mux17~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N28
cycloneive_lcell_comb \Mux17~11 (
// Equation(s):
// \Mux17~11_combout  = (\Mux17~10_combout  & ((\registerArray[7][14]~q ) # ((!cuifregS_1)))) # (!\Mux17~10_combout  & (((\registerArray[6][14]~q  & cuifregS_1))))

	.dataa(\registerArray[7][14]~q ),
	.datab(\registerArray[6][14]~q ),
	.datac(\Mux17~10_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux17~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~11 .lut_mask = 16'hACF0;
defparam \Mux17~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N8
cycloneive_lcell_comb \Mux17~19 (
// Equation(s):
// \Mux17~19_combout  = (cuifregS_2 & ((\Mux17~16_combout  & (\Mux17~18_combout )) # (!\Mux17~16_combout  & ((\Mux17~11_combout ))))) # (!cuifregS_2 & (\Mux17~16_combout ))

	.dataa(cuifregS_2),
	.datab(\Mux17~16_combout ),
	.datac(\Mux17~18_combout ),
	.datad(\Mux17~11_combout ),
	.cin(gnd),
	.combout(\Mux17~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~19 .lut_mask = 16'hE6C4;
defparam \Mux17~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y41_N27
dffeas \registerArray[21][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][14] .is_wysiwyg = "true";
defparam \registerArray[21][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N12
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// \Mux17~0_combout  = (cuifregS_3 & (((\registerArray[25][14]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[17][14]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[17][14]~q ),
	.datac(\registerArray[25][14]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'hAAE4;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N26
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// \Mux17~1_combout  = (cuifregS_2 & ((\Mux17~0_combout  & (\registerArray[29][14]~q )) # (!\Mux17~0_combout  & ((\registerArray[21][14]~q ))))) # (!cuifregS_2 & (((\Mux17~0_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[29][14]~q ),
	.datac(\registerArray[21][14]~q ),
	.datad(\Mux17~0_combout ),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hDDA0;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N16
cycloneive_lcell_comb \registerArray[23][14]~feeder (
// Equation(s):
// \registerArray[23][14]~feeder_combout  = \Mux54~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux542),
	.cin(gnd),
	.combout(\registerArray[23][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[23][14]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[23][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y44_N17
dffeas \registerArray[23][14] (
	.clk(clk),
	.d(\registerArray[23][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][14] .is_wysiwyg = "true";
defparam \registerArray[23][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N26
cycloneive_lcell_comb \Mux17~7 (
// Equation(s):
// \Mux17~7_combout  = (cuifregS_3 & ((\registerArray[27][14]~q ) # ((cuifregS_2)))) # (!cuifregS_3 & (((\registerArray[19][14]~q  & !cuifregS_2))))

	.dataa(\registerArray[27][14]~q ),
	.datab(\registerArray[19][14]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux17~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~7 .lut_mask = 16'hF0AC;
defparam \Mux17~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N4
cycloneive_lcell_comb \Mux17~8 (
// Equation(s):
// \Mux17~8_combout  = (\Mux17~7_combout  & ((\registerArray[31][14]~q ) # ((!cuifregS_2)))) # (!\Mux17~7_combout  & (((\registerArray[23][14]~q  & cuifregS_2))))

	.dataa(\registerArray[31][14]~q ),
	.datab(\registerArray[23][14]~q ),
	.datac(\Mux17~7_combout ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux17~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~8 .lut_mask = 16'hACF0;
defparam \Mux17~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N28
cycloneive_lcell_comb \Mux17~4 (
// Equation(s):
// \Mux17~4_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[20][14]~q ))) # (!cuifregS_2 & (\registerArray[16][14]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[16][14]~q ),
	.datac(\registerArray[20][14]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux17~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~4 .lut_mask = 16'hFA44;
defparam \Mux17~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N30
cycloneive_lcell_comb \Mux17~5 (
// Equation(s):
// \Mux17~5_combout  = (cuifregS_3 & ((\Mux17~4_combout  & (\registerArray[28][14]~q )) # (!\Mux17~4_combout  & ((\registerArray[24][14]~q ))))) # (!cuifregS_3 & (((\Mux17~4_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[28][14]~q ),
	.datac(\registerArray[24][14]~q ),
	.datad(\Mux17~4_combout ),
	.cin(gnd),
	.combout(\Mux17~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~5 .lut_mask = 16'hDDA0;
defparam \Mux17~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y32_N9
dffeas \registerArray[22][14] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux542),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][14] .is_wysiwyg = "true";
defparam \registerArray[22][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N8
cycloneive_lcell_comb \Mux17~2 (
// Equation(s):
// \Mux17~2_combout  = (cuifregS_2 & (((\registerArray[22][14]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[18][14]~q  & ((!cuifregS_3))))

	.dataa(\registerArray[18][14]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[22][14]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux17~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~2 .lut_mask = 16'hCCE2;
defparam \Mux17~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N22
cycloneive_lcell_comb \Mux17~3 (
// Equation(s):
// \Mux17~3_combout  = (\Mux17~2_combout  & ((\registerArray[30][14]~q ) # ((!cuifregS_3)))) # (!\Mux17~2_combout  & (((\registerArray[26][14]~q  & cuifregS_3))))

	.dataa(\registerArray[30][14]~q ),
	.datab(\Mux17~2_combout ),
	.datac(\registerArray[26][14]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux17~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~3 .lut_mask = 16'hB8CC;
defparam \Mux17~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N16
cycloneive_lcell_comb \Mux17~6 (
// Equation(s):
// \Mux17~6_combout  = (cuifregS_0 & (cuifregS_1)) # (!cuifregS_0 & ((cuifregS_1 & ((\Mux17~3_combout ))) # (!cuifregS_1 & (\Mux17~5_combout ))))

	.dataa(cuifregS_0),
	.datab(cuifregS_1),
	.datac(\Mux17~5_combout ),
	.datad(\Mux17~3_combout ),
	.cin(gnd),
	.combout(\Mux17~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~6 .lut_mask = 16'hDC98;
defparam \Mux17~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N10
cycloneive_lcell_comb \Mux17~9 (
// Equation(s):
// \Mux17~9_combout  = (cuifregS_0 & ((\Mux17~6_combout  & ((\Mux17~8_combout ))) # (!\Mux17~6_combout  & (\Mux17~1_combout )))) # (!cuifregS_0 & (((\Mux17~6_combout ))))

	.dataa(cuifregS_0),
	.datab(\Mux17~1_combout ),
	.datac(\Mux17~8_combout ),
	.datad(\Mux17~6_combout ),
	.cin(gnd),
	.combout(\Mux17~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~9 .lut_mask = 16'hF588;
defparam \Mux17~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N12
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// \Mux18~0_combout  = (cuifregS_2 & (((\registerArray[21][13]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[17][13]~q  & ((!cuifregS_3))))

	.dataa(\registerArray[17][13]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[21][13]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'hCCE2;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N20
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// \Mux18~1_combout  = (cuifregS_3 & ((\Mux18~0_combout  & (\registerArray[29][13]~q )) # (!\Mux18~0_combout  & ((\registerArray[25][13]~q ))))) # (!cuifregS_3 & (((\Mux18~0_combout ))))

	.dataa(\registerArray[29][13]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[25][13]~q ),
	.datad(\Mux18~0_combout ),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'hBBC0;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N28
cycloneive_lcell_comb \Mux18~7 (
// Equation(s):
// \Mux18~7_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[23][13]~q ))) # (!cuifregS_2 & (\registerArray[19][13]~q ))))

	.dataa(\registerArray[19][13]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[23][13]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux18~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~7 .lut_mask = 16'hFC22;
defparam \Mux18~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N30
cycloneive_lcell_comb \Mux18~8 (
// Equation(s):
// \Mux18~8_combout  = (cuifregS_3 & ((\Mux18~7_combout  & (\registerArray[31][13]~q )) # (!\Mux18~7_combout  & ((\registerArray[27][13]~q ))))) # (!cuifregS_3 & (((\Mux18~7_combout ))))

	.dataa(\registerArray[31][13]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[27][13]~q ),
	.datad(\Mux18~7_combout ),
	.cin(gnd),
	.combout(\Mux18~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~8 .lut_mask = 16'hBBC0;
defparam \Mux18~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N24
cycloneive_lcell_comb \Mux18~2 (
// Equation(s):
// \Mux18~2_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & ((\registerArray[26][13]~q ))) # (!cuifregS_3 & (\registerArray[18][13]~q ))))

	.dataa(\registerArray[18][13]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[26][13]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux18~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~2 .lut_mask = 16'hFC22;
defparam \Mux18~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N6
cycloneive_lcell_comb \Mux18~3 (
// Equation(s):
// \Mux18~3_combout  = (cuifregS_2 & ((\Mux18~2_combout  & (\registerArray[30][13]~q )) # (!\Mux18~2_combout  & ((\registerArray[22][13]~q ))))) # (!cuifregS_2 & (((\Mux18~2_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[30][13]~q ),
	.datac(\registerArray[22][13]~q ),
	.datad(\Mux18~2_combout ),
	.cin(gnd),
	.combout(\Mux18~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~3 .lut_mask = 16'hDDA0;
defparam \Mux18~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N6
cycloneive_lcell_comb \Mux18~4 (
// Equation(s):
// \Mux18~4_combout  = (cuifregS_3 & ((\registerArray[24][13]~q ) # ((cuifregS_2)))) # (!cuifregS_3 & (((\registerArray[16][13]~q  & !cuifregS_2))))

	.dataa(\registerArray[24][13]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[16][13]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux18~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~4 .lut_mask = 16'hCCB8;
defparam \Mux18~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y39_N28
cycloneive_lcell_comb \Mux18~5 (
// Equation(s):
// \Mux18~5_combout  = (cuifregS_2 & ((\Mux18~4_combout  & ((\registerArray[28][13]~q ))) # (!\Mux18~4_combout  & (\registerArray[20][13]~q )))) # (!cuifregS_2 & (((\Mux18~4_combout ))))

	.dataa(\registerArray[20][13]~q ),
	.datab(\registerArray[28][13]~q ),
	.datac(cuifregS_2),
	.datad(\Mux18~4_combout ),
	.cin(gnd),
	.combout(\Mux18~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~5 .lut_mask = 16'hCFA0;
defparam \Mux18~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N28
cycloneive_lcell_comb \Mux18~6 (
// Equation(s):
// \Mux18~6_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\Mux18~3_combout )) # (!cuifregS_1 & ((\Mux18~5_combout )))))

	.dataa(cuifregS_0),
	.datab(\Mux18~3_combout ),
	.datac(cuifregS_1),
	.datad(\Mux18~5_combout ),
	.cin(gnd),
	.combout(\Mux18~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~6 .lut_mask = 16'hE5E0;
defparam \Mux18~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N14
cycloneive_lcell_comb \Mux18~9 (
// Equation(s):
// \Mux18~9_combout  = (cuifregS_0 & ((\Mux18~6_combout  & ((\Mux18~8_combout ))) # (!\Mux18~6_combout  & (\Mux18~1_combout )))) # (!cuifregS_0 & (((\Mux18~6_combout ))))

	.dataa(cuifregS_0),
	.datab(\Mux18~1_combout ),
	.datac(\Mux18~8_combout ),
	.datad(\Mux18~6_combout ),
	.cin(gnd),
	.combout(\Mux18~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~9 .lut_mask = 16'hF588;
defparam \Mux18~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N9
dffeas \registerArray[9][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][13] .is_wysiwyg = "true";
defparam \registerArray[9][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N19
dffeas \registerArray[10][13] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux552),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][13] .is_wysiwyg = "true";
defparam \registerArray[10][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N18
cycloneive_lcell_comb \Mux18~10 (
// Equation(s):
// \Mux18~10_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][13]~q ))) # (!cuifregS_1 & (\registerArray[8][13]~q ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[8][13]~q ),
	.datac(\registerArray[10][13]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux18~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~10 .lut_mask = 16'hFA44;
defparam \Mux18~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N8
cycloneive_lcell_comb \Mux18~11 (
// Equation(s):
// \Mux18~11_combout  = (cuifregS_0 & ((\Mux18~10_combout  & (\registerArray[11][13]~q )) # (!\Mux18~10_combout  & ((\registerArray[9][13]~q ))))) # (!cuifregS_0 & (((\Mux18~10_combout ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[11][13]~q ),
	.datac(\registerArray[9][13]~q ),
	.datad(\Mux18~10_combout ),
	.cin(gnd),
	.combout(\Mux18~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~11 .lut_mask = 16'hDDA0;
defparam \Mux18~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N10
cycloneive_lcell_comb \Mux18~17 (
// Equation(s):
// \Mux18~17_combout  = (cuifregS_0 & (((\registerArray[13][13]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[12][13]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[12][13]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[13][13]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux18~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~17 .lut_mask = 16'hCCE2;
defparam \Mux18~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N0
cycloneive_lcell_comb \Mux18~18 (
// Equation(s):
// \Mux18~18_combout  = (\Mux18~17_combout  & ((\registerArray[15][13]~q ) # ((!cuifregS_1)))) # (!\Mux18~17_combout  & (((\registerArray[14][13]~q  & cuifregS_1))))

	.dataa(\registerArray[15][13]~q ),
	.datab(\registerArray[14][13]~q ),
	.datac(\Mux18~17_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux18~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~18 .lut_mask = 16'hACF0;
defparam \Mux18~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N20
cycloneive_lcell_comb \Mux18~14 (
// Equation(s):
// \Mux18~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][13]~q ))) # (!cuifregS_1 & (\registerArray[1][13]~q ))))

	.dataa(\registerArray[1][13]~q ),
	.datab(\registerArray[3][13]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux18~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~14 .lut_mask = 16'hC0A0;
defparam \Mux18~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N0
cycloneive_lcell_comb \Mux18~15 (
// Equation(s):
// \Mux18~15_combout  = (\Mux18~14_combout ) # ((!cuifregS_0 & (\registerArray[2][13]~q  & cuifregS_1)))

	.dataa(cuifregS_0),
	.datab(\registerArray[2][13]~q ),
	.datac(cuifregS_1),
	.datad(\Mux18~14_combout ),
	.cin(gnd),
	.combout(\Mux18~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~15 .lut_mask = 16'hFF40;
defparam \Mux18~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N2
cycloneive_lcell_comb \Mux18~12 (
// Equation(s):
// \Mux18~12_combout  = (cuifregS_0 & ((\registerArray[5][13]~q ) # ((cuifregS_1)))) # (!cuifregS_0 & (((\registerArray[4][13]~q  & !cuifregS_1))))

	.dataa(\registerArray[5][13]~q ),
	.datab(\registerArray[4][13]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux18~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~12 .lut_mask = 16'hF0AC;
defparam \Mux18~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N6
cycloneive_lcell_comb \Mux18~13 (
// Equation(s):
// \Mux18~13_combout  = (cuifregS_1 & ((\Mux18~12_combout  & (\registerArray[7][13]~q )) # (!\Mux18~12_combout  & ((\registerArray[6][13]~q ))))) # (!cuifregS_1 & (((\Mux18~12_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[7][13]~q ),
	.datac(\registerArray[6][13]~q ),
	.datad(\Mux18~12_combout ),
	.cin(gnd),
	.combout(\Mux18~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~13 .lut_mask = 16'hDDA0;
defparam \Mux18~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N6
cycloneive_lcell_comb \Mux18~16 (
// Equation(s):
// \Mux18~16_combout  = (cuifregS_2 & ((cuifregS_3) # ((\Mux18~13_combout )))) # (!cuifregS_2 & (!cuifregS_3 & (\Mux18~15_combout )))

	.dataa(cuifregS_2),
	.datab(cuifregS_3),
	.datac(\Mux18~15_combout ),
	.datad(\Mux18~13_combout ),
	.cin(gnd),
	.combout(\Mux18~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~16 .lut_mask = 16'hBA98;
defparam \Mux18~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y43_N12
cycloneive_lcell_comb \Mux18~19 (
// Equation(s):
// \Mux18~19_combout  = (cuifregS_3 & ((\Mux18~16_combout  & ((\Mux18~18_combout ))) # (!\Mux18~16_combout  & (\Mux18~11_combout )))) # (!cuifregS_3 & (((\Mux18~16_combout ))))

	.dataa(\Mux18~11_combout ),
	.datab(cuifregS_3),
	.datac(\Mux18~18_combout ),
	.datad(\Mux18~16_combout ),
	.cin(gnd),
	.combout(\Mux18~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~19 .lut_mask = 16'hF388;
defparam \Mux18~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N18
cycloneive_lcell_comb \Mux19~7 (
// Equation(s):
// \Mux19~7_combout  = (cuifregS_3 & ((\registerArray[27][12]~q ) # ((cuifregS_2)))) # (!cuifregS_3 & (((\registerArray[19][12]~q  & !cuifregS_2))))

	.dataa(\registerArray[27][12]~q ),
	.datab(\registerArray[19][12]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux19~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~7 .lut_mask = 16'hF0AC;
defparam \Mux19~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N0
cycloneive_lcell_comb \Mux19~8 (
// Equation(s):
// \Mux19~8_combout  = (cuifregS_2 & ((\Mux19~7_combout  & (\registerArray[31][12]~q )) # (!\Mux19~7_combout  & ((\registerArray[23][12]~q ))))) # (!cuifregS_2 & (((\Mux19~7_combout ))))

	.dataa(\registerArray[31][12]~q ),
	.datab(\registerArray[23][12]~q ),
	.datac(cuifregS_2),
	.datad(\Mux19~7_combout ),
	.cin(gnd),
	.combout(\Mux19~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~8 .lut_mask = 16'hAFC0;
defparam \Mux19~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N10
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (cuifregS_3 & ((\registerArray[25][12]~q ) # ((cuifregS_2)))) # (!cuifregS_3 & (((\registerArray[17][12]~q  & !cuifregS_2))))

	.dataa(\registerArray[25][12]~q ),
	.datab(\registerArray[17][12]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'hF0AC;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N16
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// \Mux19~1_combout  = (cuifregS_2 & ((\Mux19~0_combout  & ((\registerArray[29][12]~q ))) # (!\Mux19~0_combout  & (\registerArray[21][12]~q )))) # (!cuifregS_2 & (((\Mux19~0_combout ))))

	.dataa(\registerArray[21][12]~q ),
	.datab(\registerArray[29][12]~q ),
	.datac(cuifregS_2),
	.datad(\Mux19~0_combout ),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'hCFA0;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N31
dffeas \registerArray[24][12] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux562),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][12] .is_wysiwyg = "true";
defparam \registerArray[24][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N20
cycloneive_lcell_comb \Mux19~4 (
// Equation(s):
// \Mux19~4_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[20][12]~q ))) # (!cuifregS_2 & (\registerArray[16][12]~q ))))

	.dataa(\registerArray[16][12]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[20][12]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux19~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~4 .lut_mask = 16'hFC22;
defparam \Mux19~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N30
cycloneive_lcell_comb \Mux19~5 (
// Equation(s):
// \Mux19~5_combout  = (cuifregS_3 & ((\Mux19~4_combout  & (\registerArray[28][12]~q )) # (!\Mux19~4_combout  & ((\registerArray[24][12]~q ))))) # (!cuifregS_3 & (((\Mux19~4_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[28][12]~q ),
	.datac(\registerArray[24][12]~q ),
	.datad(\Mux19~4_combout ),
	.cin(gnd),
	.combout(\Mux19~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~5 .lut_mask = 16'hDDA0;
defparam \Mux19~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N6
cycloneive_lcell_comb \Mux19~2 (
// Equation(s):
// \Mux19~2_combout  = (cuifregS_2 & ((\registerArray[22][12]~q ) # ((cuifregS_3)))) # (!cuifregS_2 & (((\registerArray[18][12]~q  & !cuifregS_3))))

	.dataa(\registerArray[22][12]~q ),
	.datab(\registerArray[18][12]~q ),
	.datac(cuifregS_2),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~2 .lut_mask = 16'hF0AC;
defparam \Mux19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N0
cycloneive_lcell_comb \Mux19~3 (
// Equation(s):
// \Mux19~3_combout  = (cuifregS_3 & ((\Mux19~2_combout  & (\registerArray[30][12]~q )) # (!\Mux19~2_combout  & ((\registerArray[26][12]~q ))))) # (!cuifregS_3 & (((\Mux19~2_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[30][12]~q ),
	.datac(\registerArray[26][12]~q ),
	.datad(\Mux19~2_combout ),
	.cin(gnd),
	.combout(\Mux19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~3 .lut_mask = 16'hDDA0;
defparam \Mux19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N6
cycloneive_lcell_comb \Mux19~6 (
// Equation(s):
// \Mux19~6_combout  = (cuifregS_0 & (cuifregS_1)) # (!cuifregS_0 & ((cuifregS_1 & ((\Mux19~3_combout ))) # (!cuifregS_1 & (\Mux19~5_combout ))))

	.dataa(cuifregS_0),
	.datab(cuifregS_1),
	.datac(\Mux19~5_combout ),
	.datad(\Mux19~3_combout ),
	.cin(gnd),
	.combout(\Mux19~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~6 .lut_mask = 16'hDC98;
defparam \Mux19~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N14
cycloneive_lcell_comb \Mux19~9 (
// Equation(s):
// \Mux19~9_combout  = (cuifregS_0 & ((\Mux19~6_combout  & (\Mux19~8_combout )) # (!\Mux19~6_combout  & ((\Mux19~1_combout ))))) # (!cuifregS_0 & (((\Mux19~6_combout ))))

	.dataa(cuifregS_0),
	.datab(\Mux19~8_combout ),
	.datac(\Mux19~1_combout ),
	.datad(\Mux19~6_combout ),
	.cin(gnd),
	.combout(\Mux19~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~9 .lut_mask = 16'hDDA0;
defparam \Mux19~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N20
cycloneive_lcell_comb \Mux19~10 (
// Equation(s):
// \Mux19~10_combout  = (cuifregS_0 & (((\registerArray[5][12]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[4][12]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[4][12]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[5][12]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux19~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~10 .lut_mask = 16'hCCE2;
defparam \Mux19~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N8
cycloneive_lcell_comb \Mux19~11 (
// Equation(s):
// \Mux19~11_combout  = (cuifregS_1 & ((\Mux19~10_combout  & (\registerArray[7][12]~q )) # (!\Mux19~10_combout  & ((\registerArray[6][12]~q ))))) # (!cuifregS_1 & (((\Mux19~10_combout ))))

	.dataa(\registerArray[7][12]~q ),
	.datab(cuifregS_1),
	.datac(\registerArray[6][12]~q ),
	.datad(\Mux19~10_combout ),
	.cin(gnd),
	.combout(\Mux19~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~11 .lut_mask = 16'hBBC0;
defparam \Mux19~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N18
cycloneive_lcell_comb \registerArray[13][12]~feeder (
// Equation(s):
// \registerArray[13][12]~feeder_combout  = \Mux56~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux562),
	.cin(gnd),
	.combout(\registerArray[13][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[13][12]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[13][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y36_N19
dffeas \registerArray[13][12] (
	.clk(clk),
	.d(\registerArray[13][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][12] .is_wysiwyg = "true";
defparam \registerArray[13][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N0
cycloneive_lcell_comb \Mux19~17 (
// Equation(s):
// \Mux19~17_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & ((\registerArray[13][12]~q ))) # (!cuifregS_0 & (\registerArray[12][12]~q ))))

	.dataa(\registerArray[12][12]~q ),
	.datab(\registerArray[13][12]~q ),
	.datac(cuifregS_1),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux19~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~17 .lut_mask = 16'hFC0A;
defparam \Mux19~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y36_N26
cycloneive_lcell_comb \Mux19~18 (
// Equation(s):
// \Mux19~18_combout  = (cuifregS_1 & ((\Mux19~17_combout  & ((\registerArray[15][12]~q ))) # (!\Mux19~17_combout  & (\registerArray[14][12]~q )))) # (!cuifregS_1 & (((\Mux19~17_combout ))))

	.dataa(\registerArray[14][12]~q ),
	.datab(\registerArray[15][12]~q ),
	.datac(cuifregS_1),
	.datad(\Mux19~17_combout ),
	.cin(gnd),
	.combout(\Mux19~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~18 .lut_mask = 16'hCFA0;
defparam \Mux19~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N8
cycloneive_lcell_comb \Mux19~15 (
// Equation(s):
// \Mux19~15_combout  = (\Mux19~14_combout ) # ((\registerArray[2][12]~q  & (!cuifregS_0 & cuifregS_1)))

	.dataa(\Mux19~14_combout ),
	.datab(\registerArray[2][12]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux19~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~15 .lut_mask = 16'hAEAA;
defparam \Mux19~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N16
cycloneive_lcell_comb \Mux19~12 (
// Equation(s):
// \Mux19~12_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][12]~q ))) # (!cuifregS_1 & (\registerArray[8][12]~q ))))

	.dataa(\registerArray[8][12]~q ),
	.datab(\registerArray[10][12]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux19~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~12 .lut_mask = 16'hFC0A;
defparam \Mux19~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N18
cycloneive_lcell_comb \Mux19~13 (
// Equation(s):
// \Mux19~13_combout  = (cuifregS_0 & ((\Mux19~12_combout  & (\registerArray[11][12]~q )) # (!\Mux19~12_combout  & ((\registerArray[9][12]~q ))))) # (!cuifregS_0 & (((\Mux19~12_combout ))))

	.dataa(\registerArray[11][12]~q ),
	.datab(\registerArray[9][12]~q ),
	.datac(cuifregS_0),
	.datad(\Mux19~12_combout ),
	.cin(gnd),
	.combout(\Mux19~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~13 .lut_mask = 16'hAFC0;
defparam \Mux19~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N18
cycloneive_lcell_comb \Mux19~16 (
// Equation(s):
// \Mux19~16_combout  = (cuifregS_3 & ((cuifregS_2) # ((\Mux19~13_combout )))) # (!cuifregS_3 & (!cuifregS_2 & (\Mux19~15_combout )))

	.dataa(cuifregS_3),
	.datab(cuifregS_2),
	.datac(\Mux19~15_combout ),
	.datad(\Mux19~13_combout ),
	.cin(gnd),
	.combout(\Mux19~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~16 .lut_mask = 16'hBA98;
defparam \Mux19~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N24
cycloneive_lcell_comb \Mux19~19 (
// Equation(s):
// \Mux19~19_combout  = (cuifregS_2 & ((\Mux19~16_combout  & ((\Mux19~18_combout ))) # (!\Mux19~16_combout  & (\Mux19~11_combout )))) # (!cuifregS_2 & (((\Mux19~16_combout ))))

	.dataa(\Mux19~11_combout ),
	.datab(cuifregS_2),
	.datac(\Mux19~18_combout ),
	.datad(\Mux19~16_combout ),
	.cin(gnd),
	.combout(\Mux19~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~19 .lut_mask = 16'hF388;
defparam \Mux19~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N4
cycloneive_lcell_comb \Mux20~2 (
// Equation(s):
// \Mux20~2_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & ((\registerArray[26][11]~q ))) # (!cuifregS_3 & (\registerArray[18][11]~q ))))

	.dataa(\registerArray[18][11]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[26][11]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux20~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~2 .lut_mask = 16'hFC22;
defparam \Mux20~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N22
cycloneive_lcell_comb \Mux20~3 (
// Equation(s):
// \Mux20~3_combout  = (\Mux20~2_combout  & ((\registerArray[30][11]~q ) # ((!cuifregS_2)))) # (!\Mux20~2_combout  & (((\registerArray[22][11]~q  & cuifregS_2))))

	.dataa(\registerArray[30][11]~q ),
	.datab(\Mux20~2_combout ),
	.datac(\registerArray[22][11]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux20~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~3 .lut_mask = 16'hB8CC;
defparam \Mux20~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N5
dffeas \registerArray[24][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][11] .is_wysiwyg = "true";
defparam \registerArray[24][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N4
cycloneive_lcell_comb \Mux20~4 (
// Equation(s):
// \Mux20~4_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & ((\registerArray[24][11]~q ))) # (!cuifregS_3 & (\registerArray[16][11]~q ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[16][11]~q ),
	.datac(\registerArray[24][11]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux20~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~4 .lut_mask = 16'hFA44;
defparam \Mux20~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N14
cycloneive_lcell_comb \Mux20~5 (
// Equation(s):
// \Mux20~5_combout  = (\Mux20~4_combout  & ((\registerArray[28][11]~q ) # ((!cuifregS_2)))) # (!\Mux20~4_combout  & (((\registerArray[20][11]~q  & cuifregS_2))))

	.dataa(\registerArray[28][11]~q ),
	.datab(\Mux20~4_combout ),
	.datac(\registerArray[20][11]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux20~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~5 .lut_mask = 16'hB8CC;
defparam \Mux20~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N0
cycloneive_lcell_comb \Mux20~6 (
// Equation(s):
// \Mux20~6_combout  = (cuifregS_0 & (cuifregS_1)) # (!cuifregS_0 & ((cuifregS_1 & (\Mux20~3_combout )) # (!cuifregS_1 & ((\Mux20~5_combout )))))

	.dataa(cuifregS_0),
	.datab(cuifregS_1),
	.datac(\Mux20~3_combout ),
	.datad(\Mux20~5_combout ),
	.cin(gnd),
	.combout(\Mux20~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~6 .lut_mask = 16'hD9C8;
defparam \Mux20~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N14
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// \Mux20~0_combout  = (cuifregS_2 & (((\registerArray[21][11]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[17][11]~q  & ((!cuifregS_3))))

	.dataa(\registerArray[17][11]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[21][11]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'hCCE2;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N0
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// \Mux20~1_combout  = (cuifregS_3 & ((\Mux20~0_combout  & (\registerArray[29][11]~q )) # (!\Mux20~0_combout  & ((\registerArray[25][11]~q ))))) # (!cuifregS_3 & (((\Mux20~0_combout ))))

	.dataa(\registerArray[29][11]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[25][11]~q ),
	.datad(\Mux20~0_combout ),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'hBBC0;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N10
cycloneive_lcell_comb \Mux20~7 (
// Equation(s):
// \Mux20~7_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[23][11]~q ))) # (!cuifregS_2 & (\registerArray[19][11]~q ))))

	.dataa(\registerArray[19][11]~q ),
	.datab(\registerArray[23][11]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux20~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~7 .lut_mask = 16'hFC0A;
defparam \Mux20~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y44_N20
cycloneive_lcell_comb \Mux20~8 (
// Equation(s):
// \Mux20~8_combout  = (cuifregS_3 & ((\Mux20~7_combout  & (\registerArray[31][11]~q )) # (!\Mux20~7_combout  & ((\registerArray[27][11]~q ))))) # (!cuifregS_3 & (((\Mux20~7_combout ))))

	.dataa(\registerArray[31][11]~q ),
	.datab(\registerArray[27][11]~q ),
	.datac(cuifregS_3),
	.datad(\Mux20~7_combout ),
	.cin(gnd),
	.combout(\Mux20~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~8 .lut_mask = 16'hAFC0;
defparam \Mux20~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N14
cycloneive_lcell_comb \Mux20~9 (
// Equation(s):
// \Mux20~9_combout  = (cuifregS_0 & ((\Mux20~6_combout  & ((\Mux20~8_combout ))) # (!\Mux20~6_combout  & (\Mux20~1_combout )))) # (!cuifregS_0 & (\Mux20~6_combout ))

	.dataa(cuifregS_0),
	.datab(\Mux20~6_combout ),
	.datac(\Mux20~1_combout ),
	.datad(\Mux20~8_combout ),
	.cin(gnd),
	.combout(\Mux20~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~9 .lut_mask = 16'hEC64;
defparam \Mux20~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y39_N16
cycloneive_lcell_comb \registerArray[9][11]~feeder (
// Equation(s):
// \registerArray[9][11]~feeder_combout  = \Mux57~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux572),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[9][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[9][11]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[9][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y39_N17
dffeas \registerArray[9][11] (
	.clk(clk),
	.d(\registerArray[9][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][11] .is_wysiwyg = "true";
defparam \registerArray[9][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y43_N9
dffeas \registerArray[10][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][11] .is_wysiwyg = "true";
defparam \registerArray[10][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N8
cycloneive_lcell_comb \Mux20~10 (
// Equation(s):
// \Mux20~10_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][11]~q ))) # (!cuifregS_1 & (\registerArray[8][11]~q ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[8][11]~q ),
	.datac(\registerArray[10][11]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux20~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~10 .lut_mask = 16'hFA44;
defparam \Mux20~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N18
cycloneive_lcell_comb \Mux20~11 (
// Equation(s):
// \Mux20~11_combout  = (cuifregS_0 & ((\Mux20~10_combout  & ((\registerArray[11][11]~q ))) # (!\Mux20~10_combout  & (\registerArray[9][11]~q )))) # (!cuifregS_0 & (((\Mux20~10_combout ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[9][11]~q ),
	.datac(\Mux20~10_combout ),
	.datad(\registerArray[11][11]~q ),
	.cin(gnd),
	.combout(\Mux20~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~11 .lut_mask = 16'hF858;
defparam \Mux20~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N17
dffeas \registerArray[13][11] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux572),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][11] .is_wysiwyg = "true";
defparam \registerArray[13][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N16
cycloneive_lcell_comb \Mux20~17 (
// Equation(s):
// \Mux20~17_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & ((\registerArray[13][11]~q ))) # (!cuifregS_0 & (\registerArray[12][11]~q ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[12][11]~q ),
	.datac(\registerArray[13][11]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux20~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~17 .lut_mask = 16'hFA44;
defparam \Mux20~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N18
cycloneive_lcell_comb \Mux20~18 (
// Equation(s):
// \Mux20~18_combout  = (cuifregS_1 & ((\Mux20~17_combout  & (\registerArray[15][11]~q )) # (!\Mux20~17_combout  & ((\registerArray[14][11]~q ))))) # (!cuifregS_1 & (((\Mux20~17_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[15][11]~q ),
	.datac(\registerArray[14][11]~q ),
	.datad(\Mux20~17_combout ),
	.cin(gnd),
	.combout(\Mux20~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~18 .lut_mask = 16'hDDA0;
defparam \Mux20~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N12
cycloneive_lcell_comb \Mux20~12 (
// Equation(s):
// \Mux20~12_combout  = (cuifregS_0 & (((\registerArray[5][11]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[4][11]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[4][11]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[5][11]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux20~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~12 .lut_mask = 16'hCCE2;
defparam \Mux20~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N20
cycloneive_lcell_comb \Mux20~13 (
// Equation(s):
// \Mux20~13_combout  = (cuifregS_1 & ((\Mux20~12_combout  & (\registerArray[7][11]~q )) # (!\Mux20~12_combout  & ((\registerArray[6][11]~q ))))) # (!cuifregS_1 & (((\Mux20~12_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[7][11]~q ),
	.datac(\registerArray[6][11]~q ),
	.datad(\Mux20~12_combout ),
	.cin(gnd),
	.combout(\Mux20~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~13 .lut_mask = 16'hDDA0;
defparam \Mux20~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N0
cycloneive_lcell_comb \Mux20~14 (
// Equation(s):
// \Mux20~14_combout  = (cuifregS_0 & ((cuifregS_1 & (\registerArray[3][11]~q )) # (!cuifregS_1 & ((\registerArray[1][11]~q )))))

	.dataa(cuifregS_1),
	.datab(\registerArray[3][11]~q ),
	.datac(\registerArray[1][11]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux20~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~14 .lut_mask = 16'hD800;
defparam \Mux20~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N28
cycloneive_lcell_comb \Mux20~15 (
// Equation(s):
// \Mux20~15_combout  = (\Mux20~14_combout ) # ((!cuifregS_0 & (cuifregS_1 & \registerArray[2][11]~q )))

	.dataa(cuifregS_0),
	.datab(cuifregS_1),
	.datac(\registerArray[2][11]~q ),
	.datad(\Mux20~14_combout ),
	.cin(gnd),
	.combout(\Mux20~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~15 .lut_mask = 16'hFF40;
defparam \Mux20~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N2
cycloneive_lcell_comb \Mux20~16 (
// Equation(s):
// \Mux20~16_combout  = (cuifregS_2 & ((cuifregS_3) # ((\Mux20~13_combout )))) # (!cuifregS_2 & (!cuifregS_3 & ((\Mux20~15_combout ))))

	.dataa(cuifregS_2),
	.datab(cuifregS_3),
	.datac(\Mux20~13_combout ),
	.datad(\Mux20~15_combout ),
	.cin(gnd),
	.combout(\Mux20~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~16 .lut_mask = 16'hB9A8;
defparam \Mux20~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N24
cycloneive_lcell_comb \Mux20~19 (
// Equation(s):
// \Mux20~19_combout  = (cuifregS_3 & ((\Mux20~16_combout  & ((\Mux20~18_combout ))) # (!\Mux20~16_combout  & (\Mux20~11_combout )))) # (!cuifregS_3 & (((\Mux20~16_combout ))))

	.dataa(\Mux20~11_combout ),
	.datab(cuifregS_3),
	.datac(\Mux20~18_combout ),
	.datad(\Mux20~16_combout ),
	.cin(gnd),
	.combout(\Mux20~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~19 .lut_mask = 16'hF388;
defparam \Mux20~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N8
cycloneive_lcell_comb \Mux21~7 (
// Equation(s):
// \Mux21~7_combout  = (cuifregS_3 & (((\registerArray[27][10]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[19][10]~q  & ((!cuifregS_2))))

	.dataa(\registerArray[19][10]~q ),
	.datab(\registerArray[27][10]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux21~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~7 .lut_mask = 16'hF0CA;
defparam \Mux21~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N14
cycloneive_lcell_comb \Mux21~8 (
// Equation(s):
// \Mux21~8_combout  = (\Mux21~7_combout  & (((\registerArray[31][10]~q ) # (!cuifregS_2)))) # (!\Mux21~7_combout  & (\registerArray[23][10]~q  & ((cuifregS_2))))

	.dataa(\registerArray[23][10]~q ),
	.datab(\registerArray[31][10]~q ),
	.datac(\Mux21~7_combout ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux21~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~8 .lut_mask = 16'hCAF0;
defparam \Mux21~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N16
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// \Mux21~0_combout  = (cuifregS_3 & (((\registerArray[25][10]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[17][10]~q  & ((!cuifregS_2))))

	.dataa(\registerArray[17][10]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[25][10]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hCCE2;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N30
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// \Mux21~1_combout  = (cuifregS_2 & ((\Mux21~0_combout  & ((\registerArray[29][10]~q ))) # (!\Mux21~0_combout  & (\registerArray[21][10]~q )))) # (!cuifregS_2 & (((\Mux21~0_combout ))))

	.dataa(\registerArray[21][10]~q ),
	.datab(\registerArray[29][10]~q ),
	.datac(cuifregS_2),
	.datad(\Mux21~0_combout ),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'hCFA0;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N23
dffeas \registerArray[24][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][10] .is_wysiwyg = "true";
defparam \registerArray[24][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N12
cycloneive_lcell_comb \Mux21~4 (
// Equation(s):
// \Mux21~4_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[20][10]~q ))) # (!cuifregS_2 & (\registerArray[16][10]~q ))))

	.dataa(\registerArray[16][10]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[20][10]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux21~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~4 .lut_mask = 16'hFC22;
defparam \Mux21~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N22
cycloneive_lcell_comb \Mux21~5 (
// Equation(s):
// \Mux21~5_combout  = (cuifregS_3 & ((\Mux21~4_combout  & (\registerArray[28][10]~q )) # (!\Mux21~4_combout  & ((\registerArray[24][10]~q ))))) # (!cuifregS_3 & (((\Mux21~4_combout ))))

	.dataa(\registerArray[28][10]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[24][10]~q ),
	.datad(\Mux21~4_combout ),
	.cin(gnd),
	.combout(\Mux21~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~5 .lut_mask = 16'hBBC0;
defparam \Mux21~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N17
dffeas \registerArray[22][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][10] .is_wysiwyg = "true";
defparam \registerArray[22][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N16
cycloneive_lcell_comb \Mux21~2 (
// Equation(s):
// \Mux21~2_combout  = (cuifregS_2 & (((\registerArray[22][10]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[18][10]~q  & ((!cuifregS_3))))

	.dataa(\registerArray[18][10]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[22][10]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux21~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~2 .lut_mask = 16'hCCE2;
defparam \Mux21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N26
cycloneive_lcell_comb \Mux21~3 (
// Equation(s):
// \Mux21~3_combout  = (cuifregS_3 & ((\Mux21~2_combout  & (\registerArray[30][10]~q )) # (!\Mux21~2_combout  & ((\registerArray[26][10]~q ))))) # (!cuifregS_3 & (((\Mux21~2_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[30][10]~q ),
	.datac(\registerArray[26][10]~q ),
	.datad(\Mux21~2_combout ),
	.cin(gnd),
	.combout(\Mux21~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~3 .lut_mask = 16'hDDA0;
defparam \Mux21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N0
cycloneive_lcell_comb \Mux21~6 (
// Equation(s):
// \Mux21~6_combout  = (cuifregS_1 & (((cuifregS_0) # (\Mux21~3_combout )))) # (!cuifregS_1 & (\Mux21~5_combout  & (!cuifregS_0)))

	.dataa(cuifregS_1),
	.datab(\Mux21~5_combout ),
	.datac(cuifregS_0),
	.datad(\Mux21~3_combout ),
	.cin(gnd),
	.combout(\Mux21~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~6 .lut_mask = 16'hAEA4;
defparam \Mux21~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N22
cycloneive_lcell_comb \Mux21~9 (
// Equation(s):
// \Mux21~9_combout  = (cuifregS_0 & ((\Mux21~6_combout  & (\Mux21~8_combout )) # (!\Mux21~6_combout  & ((\Mux21~1_combout ))))) # (!cuifregS_0 & (((\Mux21~6_combout ))))

	.dataa(cuifregS_0),
	.datab(\Mux21~8_combout ),
	.datac(\Mux21~1_combout ),
	.datad(\Mux21~6_combout ),
	.cin(gnd),
	.combout(\Mux21~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~9 .lut_mask = 16'hDDA0;
defparam \Mux21~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y32_N11
dffeas \registerArray[12][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][10] .is_wysiwyg = "true";
defparam \registerArray[12][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N12
cycloneive_lcell_comb \Mux21~17 (
// Equation(s):
// \Mux21~17_combout  = (cuifregS_0 & ((\registerArray[13][10]~q ) # ((cuifregS_1)))) # (!cuifregS_0 & (((\registerArray[12][10]~q  & !cuifregS_1))))

	.dataa(\registerArray[13][10]~q ),
	.datab(\registerArray[12][10]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux21~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~17 .lut_mask = 16'hF0AC;
defparam \Mux21~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y42_N2
cycloneive_lcell_comb \Mux21~18 (
// Equation(s):
// \Mux21~18_combout  = (cuifregS_1 & ((\Mux21~17_combout  & (\registerArray[15][10]~q )) # (!\Mux21~17_combout  & ((\registerArray[14][10]~q ))))) # (!cuifregS_1 & (((\Mux21~17_combout ))))

	.dataa(\registerArray[15][10]~q ),
	.datab(\registerArray[14][10]~q ),
	.datac(cuifregS_1),
	.datad(\Mux21~17_combout ),
	.cin(gnd),
	.combout(\Mux21~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~18 .lut_mask = 16'hAFC0;
defparam \Mux21~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N17
dffeas \registerArray[5][10] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux582),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][10] .is_wysiwyg = "true";
defparam \registerArray[5][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N16
cycloneive_lcell_comb \Mux21~10 (
// Equation(s):
// \Mux21~10_combout  = (cuifregS_0 & (((\registerArray[5][10]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[4][10]~q  & ((!cuifregS_1))))

	.dataa(cuifregS_0),
	.datab(\registerArray[4][10]~q ),
	.datac(\registerArray[5][10]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux21~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~10 .lut_mask = 16'hAAE4;
defparam \Mux21~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N8
cycloneive_lcell_comb \Mux21~11 (
// Equation(s):
// \Mux21~11_combout  = (\Mux21~10_combout  & (((\registerArray[7][10]~q ) # (!cuifregS_1)))) # (!\Mux21~10_combout  & (\registerArray[6][10]~q  & ((cuifregS_1))))

	.dataa(\registerArray[6][10]~q ),
	.datab(\registerArray[7][10]~q ),
	.datac(\Mux21~10_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux21~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~11 .lut_mask = 16'hCAF0;
defparam \Mux21~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N28
cycloneive_lcell_comb \Mux21~13 (
// Equation(s):
// \Mux21~13_combout  = (\Mux21~12_combout  & ((\registerArray[11][10]~q ) # ((!cuifregS_0)))) # (!\Mux21~12_combout  & (((\registerArray[9][10]~q  & cuifregS_0))))

	.dataa(\Mux21~12_combout ),
	.datab(\registerArray[11][10]~q ),
	.datac(\registerArray[9][10]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux21~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~13 .lut_mask = 16'hD8AA;
defparam \Mux21~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N2
cycloneive_lcell_comb \Mux21~16 (
// Equation(s):
// \Mux21~16_combout  = (cuifregS_3 & (((cuifregS_2) # (\Mux21~13_combout )))) # (!cuifregS_3 & (\Mux21~15_combout  & (!cuifregS_2)))

	.dataa(\Mux21~15_combout ),
	.datab(cuifregS_3),
	.datac(cuifregS_2),
	.datad(\Mux21~13_combout ),
	.cin(gnd),
	.combout(\Mux21~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~16 .lut_mask = 16'hCEC2;
defparam \Mux21~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N24
cycloneive_lcell_comb \Mux21~19 (
// Equation(s):
// \Mux21~19_combout  = (cuifregS_2 & ((\Mux21~16_combout  & (\Mux21~18_combout )) # (!\Mux21~16_combout  & ((\Mux21~11_combout ))))) # (!cuifregS_2 & (((\Mux21~16_combout ))))

	.dataa(\Mux21~18_combout ),
	.datab(cuifregS_2),
	.datac(\Mux21~11_combout ),
	.datad(\Mux21~16_combout ),
	.cin(gnd),
	.combout(\Mux21~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~19 .lut_mask = 16'hBBC0;
defparam \Mux21~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N16
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// \Mux22~0_combout  = (cuifregS_2 & (((\registerArray[21][9]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[17][9]~q  & ((!cuifregS_3))))

	.dataa(\registerArray[17][9]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[21][9]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'hCCE2;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N4
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// \Mux22~1_combout  = (cuifregS_3 & ((\Mux22~0_combout  & (\registerArray[29][9]~q )) # (!\Mux22~0_combout  & ((\registerArray[25][9]~q ))))) # (!cuifregS_3 & (((\Mux22~0_combout ))))

	.dataa(\registerArray[29][9]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[25][9]~q ),
	.datad(\Mux22~0_combout ),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'hBBC0;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N0
cycloneive_lcell_comb \Mux22~2 (
// Equation(s):
// \Mux22~2_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & ((\registerArray[26][9]~q ))) # (!cuifregS_3 & (\registerArray[18][9]~q ))))

	.dataa(\registerArray[18][9]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[26][9]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux22~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~2 .lut_mask = 16'hFC22;
defparam \Mux22~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N18
cycloneive_lcell_comb \Mux22~3 (
// Equation(s):
// \Mux22~3_combout  = (cuifregS_2 & ((\Mux22~2_combout  & (\registerArray[30][9]~q )) # (!\Mux22~2_combout  & ((\registerArray[22][9]~q ))))) # (!cuifregS_2 & (((\Mux22~2_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[30][9]~q ),
	.datac(\registerArray[22][9]~q ),
	.datad(\Mux22~2_combout ),
	.cin(gnd),
	.combout(\Mux22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~3 .lut_mask = 16'hDDA0;
defparam \Mux22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N24
cycloneive_lcell_comb \Mux22~4 (
// Equation(s):
// \Mux22~4_combout  = (cuifregS_3 & (((\registerArray[24][9]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[16][9]~q  & ((!cuifregS_2))))

	.dataa(\registerArray[16][9]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[24][9]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux22~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~4 .lut_mask = 16'hCCE2;
defparam \Mux22~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N7
dffeas \registerArray[20][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][9] .is_wysiwyg = "true";
defparam \registerArray[20][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N6
cycloneive_lcell_comb \Mux22~5 (
// Equation(s):
// \Mux22~5_combout  = (\Mux22~4_combout  & ((\registerArray[28][9]~q ) # ((!cuifregS_2)))) # (!\Mux22~4_combout  & (((\registerArray[20][9]~q  & cuifregS_2))))

	.dataa(\registerArray[28][9]~q ),
	.datab(\Mux22~4_combout ),
	.datac(\registerArray[20][9]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux22~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~5 .lut_mask = 16'hB8CC;
defparam \Mux22~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N4
cycloneive_lcell_comb \Mux22~6 (
// Equation(s):
// \Mux22~6_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\Mux22~3_combout )) # (!cuifregS_1 & ((\Mux22~5_combout )))))

	.dataa(cuifregS_0),
	.datab(\Mux22~3_combout ),
	.datac(cuifregS_1),
	.datad(\Mux22~5_combout ),
	.cin(gnd),
	.combout(\Mux22~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~6 .lut_mask = 16'hE5E0;
defparam \Mux22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N7
dffeas \registerArray[27][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][9] .is_wysiwyg = "true";
defparam \registerArray[27][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N24
cycloneive_lcell_comb \Mux22~7 (
// Equation(s):
// \Mux22~7_combout  = (cuifregS_2 & (((\registerArray[23][9]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[19][9]~q  & ((!cuifregS_3))))

	.dataa(\registerArray[19][9]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[23][9]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux22~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~7 .lut_mask = 16'hCCE2;
defparam \Mux22~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N6
cycloneive_lcell_comb \Mux22~8 (
// Equation(s):
// \Mux22~8_combout  = (cuifregS_3 & ((\Mux22~7_combout  & (\registerArray[31][9]~q )) # (!\Mux22~7_combout  & ((\registerArray[27][9]~q ))))) # (!cuifregS_3 & (((\Mux22~7_combout ))))

	.dataa(\registerArray[31][9]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[27][9]~q ),
	.datad(\Mux22~7_combout ),
	.cin(gnd),
	.combout(\Mux22~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~8 .lut_mask = 16'hBBC0;
defparam \Mux22~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N26
cycloneive_lcell_comb \Mux22~9 (
// Equation(s):
// \Mux22~9_combout  = (cuifregS_0 & ((\Mux22~6_combout  & ((\Mux22~8_combout ))) # (!\Mux22~6_combout  & (\Mux22~1_combout )))) # (!cuifregS_0 & (((\Mux22~6_combout ))))

	.dataa(\Mux22~1_combout ),
	.datab(cuifregS_0),
	.datac(\Mux22~6_combout ),
	.datad(\Mux22~8_combout ),
	.cin(gnd),
	.combout(\Mux22~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~9 .lut_mask = 16'hF838;
defparam \Mux22~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N21
dffeas \registerArray[13][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][9] .is_wysiwyg = "true";
defparam \registerArray[13][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N20
cycloneive_lcell_comb \Mux22~17 (
// Equation(s):
// \Mux22~17_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & ((\registerArray[13][9]~q ))) # (!cuifregS_0 & (\registerArray[12][9]~q ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[12][9]~q ),
	.datac(\registerArray[13][9]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux22~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~17 .lut_mask = 16'hFA44;
defparam \Mux22~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N30
cycloneive_lcell_comb \Mux22~18 (
// Equation(s):
// \Mux22~18_combout  = (\Mux22~17_combout  & ((\registerArray[15][9]~q ) # ((!cuifregS_1)))) # (!\Mux22~17_combout  & (((\registerArray[14][9]~q  & cuifregS_1))))

	.dataa(\registerArray[15][9]~q ),
	.datab(\Mux22~17_combout ),
	.datac(\registerArray[14][9]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux22~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~18 .lut_mask = 16'hB8CC;
defparam \Mux22~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N15
dffeas \registerArray[10][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][9] .is_wysiwyg = "true";
defparam \registerArray[10][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N14
cycloneive_lcell_comb \Mux22~10 (
// Equation(s):
// \Mux22~10_combout  = (cuifregS_1 & (((\registerArray[10][9]~q ) # (cuifregS_0)))) # (!cuifregS_1 & (\registerArray[8][9]~q  & ((!cuifregS_0))))

	.dataa(cuifregS_1),
	.datab(\registerArray[8][9]~q ),
	.datac(\registerArray[10][9]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux22~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~10 .lut_mask = 16'hAAE4;
defparam \Mux22~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N20
cycloneive_lcell_comb \Mux22~11 (
// Equation(s):
// \Mux22~11_combout  = (\Mux22~10_combout  & ((\registerArray[11][9]~q ) # ((!cuifregS_0)))) # (!\Mux22~10_combout  & (((\registerArray[9][9]~q  & cuifregS_0))))

	.dataa(\registerArray[11][9]~q ),
	.datab(\Mux22~10_combout ),
	.datac(\registerArray[9][9]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux22~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~11 .lut_mask = 16'hB8CC;
defparam \Mux22~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N0
cycloneive_lcell_comb \Mux22~12 (
// Equation(s):
// \Mux22~12_combout  = (cuifregS_0 & (((\registerArray[5][9]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[4][9]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[4][9]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[5][9]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux22~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~12 .lut_mask = 16'hCCE2;
defparam \Mux22~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N8
cycloneive_lcell_comb \Mux22~13 (
// Equation(s):
// \Mux22~13_combout  = (\Mux22~12_combout  & ((\registerArray[7][9]~q ) # ((!cuifregS_1)))) # (!\Mux22~12_combout  & (((\registerArray[6][9]~q  & cuifregS_1))))

	.dataa(\registerArray[7][9]~q ),
	.datab(\Mux22~12_combout ),
	.datac(\registerArray[6][9]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux22~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~13 .lut_mask = 16'hB8CC;
defparam \Mux22~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y42_N31
dffeas \registerArray[3][9] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux592),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][9] .is_wysiwyg = "true";
defparam \registerArray[3][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N30
cycloneive_lcell_comb \Mux22~14 (
// Equation(s):
// \Mux22~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][9]~q ))) # (!cuifregS_1 & (\registerArray[1][9]~q ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[1][9]~q ),
	.datac(\registerArray[3][9]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux22~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~14 .lut_mask = 16'hA088;
defparam \Mux22~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N16
cycloneive_lcell_comb \Mux22~15 (
// Equation(s):
// \Mux22~15_combout  = (\Mux22~14_combout ) # ((!cuifregS_0 & (\registerArray[2][9]~q  & cuifregS_1)))

	.dataa(cuifregS_0),
	.datab(\registerArray[2][9]~q ),
	.datac(\Mux22~14_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux22~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~15 .lut_mask = 16'hF4F0;
defparam \Mux22~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N2
cycloneive_lcell_comb \Mux22~16 (
// Equation(s):
// \Mux22~16_combout  = (cuifregS_2 & ((cuifregS_3) # ((\Mux22~13_combout )))) # (!cuifregS_2 & (!cuifregS_3 & ((\Mux22~15_combout ))))

	.dataa(cuifregS_2),
	.datab(cuifregS_3),
	.datac(\Mux22~13_combout ),
	.datad(\Mux22~15_combout ),
	.cin(gnd),
	.combout(\Mux22~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~16 .lut_mask = 16'hB9A8;
defparam \Mux22~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y42_N20
cycloneive_lcell_comb \Mux22~19 (
// Equation(s):
// \Mux22~19_combout  = (cuifregS_3 & ((\Mux22~16_combout  & (\Mux22~18_combout )) # (!\Mux22~16_combout  & ((\Mux22~11_combout ))))) # (!cuifregS_3 & (((\Mux22~16_combout ))))

	.dataa(cuifregS_3),
	.datab(\Mux22~18_combout ),
	.datac(\Mux22~11_combout ),
	.datad(\Mux22~16_combout ),
	.cin(gnd),
	.combout(\Mux22~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~19 .lut_mask = 16'hDDA0;
defparam \Mux22~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N0
cycloneive_lcell_comb \Mux59~4 (
// Equation(s):
// \Mux59~4_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[24][4]~q )) # (!cuifregT_3 & ((\registerArray[16][4]~q )))))

	.dataa(cuifregT_2),
	.datab(\registerArray[24][4]~q ),
	.datac(\registerArray[16][4]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux59~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~4 .lut_mask = 16'hEE50;
defparam \Mux59~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N14
cycloneive_lcell_comb \Mux59~5 (
// Equation(s):
// \Mux59~5_combout  = (cuifregT_2 & ((\Mux59~4_combout  & (\registerArray[28][4]~q )) # (!\Mux59~4_combout  & ((\registerArray[20][4]~q ))))) # (!cuifregT_2 & (\Mux59~4_combout ))

	.dataa(cuifregT_2),
	.datab(\Mux59~4_combout ),
	.datac(\registerArray[28][4]~q ),
	.datad(\registerArray[20][4]~q ),
	.cin(gnd),
	.combout(\Mux59~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~5 .lut_mask = 16'hE6C4;
defparam \Mux59~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N10
cycloneive_lcell_comb \Mux59~2 (
// Equation(s):
// \Mux59~2_combout  = (cuifregT_2 & (((cuifregT_3)))) # (!cuifregT_2 & ((cuifregT_3 & (\registerArray[26][4]~q )) # (!cuifregT_3 & ((\registerArray[18][4]~q )))))

	.dataa(\registerArray[26][4]~q ),
	.datab(cuifregT_2),
	.datac(\registerArray[18][4]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux59~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~2 .lut_mask = 16'hEE30;
defparam \Mux59~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N20
cycloneive_lcell_comb \Mux59~3 (
// Equation(s):
// \Mux59~3_combout  = (cuifregT_2 & ((\Mux59~2_combout  & ((\registerArray[30][4]~q ))) # (!\Mux59~2_combout  & (\registerArray[22][4]~q )))) # (!cuifregT_2 & (((\Mux59~2_combout ))))

	.dataa(cuifregT_2),
	.datab(\registerArray[22][4]~q ),
	.datac(\registerArray[30][4]~q ),
	.datad(\Mux59~2_combout ),
	.cin(gnd),
	.combout(\Mux59~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~3 .lut_mask = 16'hF588;
defparam \Mux59~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N4
cycloneive_lcell_comb \Mux59~6 (
// Equation(s):
// \Mux59~6_combout  = (cuifregT_01 & (cuifregT_1)) # (!cuifregT_01 & ((cuifregT_1 & ((\Mux59~3_combout ))) # (!cuifregT_1 & (\Mux59~5_combout ))))

	.dataa(cuifregT_0),
	.datab(cuifregT_1),
	.datac(\Mux59~5_combout ),
	.datad(\Mux59~3_combout ),
	.cin(gnd),
	.combout(\Mux59~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~6 .lut_mask = 16'hDC98;
defparam \Mux59~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N22
cycloneive_lcell_comb \Mux59~0 (
// Equation(s):
// \Mux59~0_combout  = (cuifregT_3 & (((cuifregT_2)))) # (!cuifregT_3 & ((cuifregT_2 & (\registerArray[21][4]~q )) # (!cuifregT_2 & ((\registerArray[17][4]~q )))))

	.dataa(\registerArray[21][4]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[17][4]~q ),
	.datad(cuifregT_2),
	.cin(gnd),
	.combout(\Mux59~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~0 .lut_mask = 16'hEE30;
defparam \Mux59~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N6
cycloneive_lcell_comb \registerArray[25][4]~feeder (
// Equation(s):
// \registerArray[25][4]~feeder_combout  = \Mux64~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux64),
	.cin(gnd),
	.combout(\registerArray[25][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[25][4]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[25][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N7
dffeas \registerArray[25][4] (
	.clk(clk),
	.d(\registerArray[25][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~60_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[25][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[25][4] .is_wysiwyg = "true";
defparam \registerArray[25][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y35_N17
dffeas \registerArray[29][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~61_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[29][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[29][4] .is_wysiwyg = "true";
defparam \registerArray[29][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N16
cycloneive_lcell_comb \Mux59~1 (
// Equation(s):
// \Mux59~1_combout  = (\Mux59~0_combout  & (((\registerArray[29][4]~q ) # (!cuifregT_3)))) # (!\Mux59~0_combout  & (\registerArray[25][4]~q  & ((cuifregT_3))))

	.dataa(\Mux59~0_combout ),
	.datab(\registerArray[25][4]~q ),
	.datac(\registerArray[29][4]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux59~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~1 .lut_mask = 16'hE4AA;
defparam \Mux59~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y33_N19
dffeas \registerArray[31][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~71_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[31][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[31][4] .is_wysiwyg = "true";
defparam \registerArray[31][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N30
cycloneive_lcell_comb \Mux59~7 (
// Equation(s):
// \Mux59~7_combout  = (cuifregT_2 & ((\registerArray[23][4]~q ) # ((cuifregT_3)))) # (!cuifregT_2 & (((\registerArray[19][4]~q  & !cuifregT_3))))

	.dataa(cuifregT_2),
	.datab(\registerArray[23][4]~q ),
	.datac(\registerArray[19][4]~q ),
	.datad(cuifregT_3),
	.cin(gnd),
	.combout(\Mux59~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~7 .lut_mask = 16'hAAD8;
defparam \Mux59~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N18
cycloneive_lcell_comb \Mux59~8 (
// Equation(s):
// \Mux59~8_combout  = (cuifregT_3 & ((\Mux59~7_combout  & ((\registerArray[31][4]~q ))) # (!\Mux59~7_combout  & (\registerArray[27][4]~q )))) # (!cuifregT_3 & (((\Mux59~7_combout ))))

	.dataa(\registerArray[27][4]~q ),
	.datab(cuifregT_3),
	.datac(\registerArray[31][4]~q ),
	.datad(\Mux59~7_combout ),
	.cin(gnd),
	.combout(\Mux59~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~8 .lut_mask = 16'hF388;
defparam \Mux59~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N4
cycloneive_lcell_comb \registerArray[10][4]~feeder (
// Equation(s):
// \registerArray[10][4]~feeder_combout  = \Mux64~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux64),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[10][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[10][4]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[10][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N5
dffeas \registerArray[10][4] (
	.clk(clk),
	.d(\registerArray[10][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][4] .is_wysiwyg = "true";
defparam \registerArray[10][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N2
cycloneive_lcell_comb \Mux59~10 (
// Equation(s):
// \Mux59~10_combout  = (cuifregT_1 & (((\registerArray[10][4]~q ) # (cuifregT_01)))) # (!cuifregT_1 & (\registerArray[8][4]~q  & ((!cuifregT_01))))

	.dataa(\registerArray[8][4]~q ),
	.datab(\registerArray[10][4]~q ),
	.datac(cuifregT_1),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux59~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~10 .lut_mask = 16'hF0CA;
defparam \Mux59~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N24
cycloneive_lcell_comb \Mux59~11 (
// Equation(s):
// \Mux59~11_combout  = (\Mux59~10_combout  & ((\registerArray[11][4]~q ) # ((!cuifregT_01)))) # (!\Mux59~10_combout  & (((\registerArray[9][4]~q  & cuifregT_01))))

	.dataa(\registerArray[11][4]~q ),
	.datab(\Mux59~10_combout ),
	.datac(\registerArray[9][4]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux59~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~11 .lut_mask = 16'hB8CC;
defparam \Mux59~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N12
cycloneive_lcell_comb \registerArray[14][4]~feeder (
// Equation(s):
// \registerArray[14][4]~feeder_combout  = \Mux64~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux64),
	.cin(gnd),
	.combout(\registerArray[14][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[14][4]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[14][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y32_N13
dffeas \registerArray[14][4] (
	.clk(clk),
	.d(\registerArray[14][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~81_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[14][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[14][4] .is_wysiwyg = "true";
defparam \registerArray[14][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N10
cycloneive_lcell_comb \registerArray[12][4]~feeder (
// Equation(s):
// \registerArray[12][4]~feeder_combout  = \Mux64~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux64),
	.cin(gnd),
	.combout(\registerArray[12][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[12][4]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[12][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y31_N11
dffeas \registerArray[12][4] (
	.clk(clk),
	.d(\registerArray[12][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~83_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[12][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[12][4] .is_wysiwyg = "true";
defparam \registerArray[12][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N22
cycloneive_lcell_comb \Mux59~17 (
// Equation(s):
// \Mux59~17_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & ((\registerArray[13][4]~q ))) # (!cuifregT_01 & (\registerArray[12][4]~q ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[12][4]~q ),
	.datac(\registerArray[13][4]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux59~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~17 .lut_mask = 16'hFA44;
defparam \Mux59~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N30
cycloneive_lcell_comb \Mux59~18 (
// Equation(s):
// \Mux59~18_combout  = (cuifregT_1 & ((\Mux59~17_combout  & ((\registerArray[15][4]~q ))) # (!\Mux59~17_combout  & (\registerArray[14][4]~q )))) # (!cuifregT_1 & (((\Mux59~17_combout ))))

	.dataa(\registerArray[14][4]~q ),
	.datab(cuifregT_1),
	.datac(\registerArray[15][4]~q ),
	.datad(\Mux59~17_combout ),
	.cin(gnd),
	.combout(\Mux59~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~18 .lut_mask = 16'hF388;
defparam \Mux59~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N12
cycloneive_lcell_comb \registerArray[1][4]~feeder (
// Equation(s):
// \registerArray[1][4]~feeder_combout  = \Mux64~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux64),
	.cin(gnd),
	.combout(\registerArray[1][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[1][4]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[1][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y42_N13
dffeas \registerArray[1][4] (
	.clk(clk),
	.d(\registerArray[1][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][4] .is_wysiwyg = "true";
defparam \registerArray[1][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N24
cycloneive_lcell_comb \Mux59~14 (
// Equation(s):
// \Mux59~14_combout  = (cuifregT_01 & ((cuifregT_1 & (\registerArray[3][4]~q )) # (!cuifregT_1 & ((\registerArray[1][4]~q )))))

	.dataa(\registerArray[3][4]~q ),
	.datab(\registerArray[1][4]~q ),
	.datac(cuifregT_0),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux59~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~14 .lut_mask = 16'hA0C0;
defparam \Mux59~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N26
cycloneive_lcell_comb \Mux59~15 (
// Equation(s):
// \Mux59~15_combout  = (\Mux59~14_combout ) # ((!cuifregT_01 & (\registerArray[2][4]~q  & cuifregT_1)))

	.dataa(cuifregT_0),
	.datab(\registerArray[2][4]~q ),
	.datac(\Mux59~14_combout ),
	.datad(cuifregT_1),
	.cin(gnd),
	.combout(\Mux59~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~15 .lut_mask = 16'hF4F0;
defparam \Mux59~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y35_N27
dffeas \registerArray[4][4] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux64),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][4] .is_wysiwyg = "true";
defparam \registerArray[4][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y35_N26
cycloneive_lcell_comb \Mux59~12 (
// Equation(s):
// \Mux59~12_combout  = (cuifregT_1 & (((cuifregT_01)))) # (!cuifregT_1 & ((cuifregT_01 & (\registerArray[5][4]~q )) # (!cuifregT_01 & ((\registerArray[4][4]~q )))))

	.dataa(cuifregT_1),
	.datab(\registerArray[5][4]~q ),
	.datac(\registerArray[4][4]~q ),
	.datad(cuifregT_0),
	.cin(gnd),
	.combout(\Mux59~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~12 .lut_mask = 16'hEE50;
defparam \Mux59~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y39_N0
cycloneive_lcell_comb \Mux59~13 (
// Equation(s):
// \Mux59~13_combout  = (cuifregT_1 & ((\Mux59~12_combout  & ((\registerArray[7][4]~q ))) # (!\Mux59~12_combout  & (\registerArray[6][4]~q )))) # (!cuifregT_1 & (((\Mux59~12_combout ))))

	.dataa(cuifregT_1),
	.datab(\registerArray[6][4]~q ),
	.datac(\registerArray[7][4]~q ),
	.datad(\Mux59~12_combout ),
	.cin(gnd),
	.combout(\Mux59~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~13 .lut_mask = 16'hF588;
defparam \Mux59~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N16
cycloneive_lcell_comb \Mux59~16 (
// Equation(s):
// \Mux59~16_combout  = (cuifregT_2 & ((cuifregT_3) # ((\Mux59~13_combout )))) # (!cuifregT_2 & (!cuifregT_3 & (\Mux59~15_combout )))

	.dataa(cuifregT_2),
	.datab(cuifregT_3),
	.datac(\Mux59~15_combout ),
	.datad(\Mux59~13_combout ),
	.cin(gnd),
	.combout(\Mux59~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~16 .lut_mask = 16'hBA98;
defparam \Mux59~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N1
dffeas \registerArray[10][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][31] .is_wysiwyg = "true";
defparam \registerArray[10][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N0
cycloneive_lcell_comb \Mux0~10 (
// Equation(s):
// \Mux0~10_combout  = (cuifregS_0 & (cuifregS_1)) # (!cuifregS_0 & ((cuifregS_1 & (\registerArray[10][31]~q )) # (!cuifregS_1 & ((\registerArray[8][31]~q )))))

	.dataa(cuifregS_0),
	.datab(cuifregS_1),
	.datac(\registerArray[10][31]~q ),
	.datad(\registerArray[8][31]~q ),
	.cin(gnd),
	.combout(\Mux0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~10 .lut_mask = 16'hD9C8;
defparam \Mux0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N20
cycloneive_lcell_comb \Mux0~11 (
// Equation(s):
// \Mux0~11_combout  = (cuifregS_0 & ((\Mux0~10_combout  & ((\registerArray[11][31]~q ))) # (!\Mux0~10_combout  & (\registerArray[9][31]~q )))) # (!cuifregS_0 & (((\Mux0~10_combout ))))

	.dataa(\registerArray[9][31]~q ),
	.datab(\registerArray[11][31]~q ),
	.datac(cuifregS_0),
	.datad(\Mux0~10_combout ),
	.cin(gnd),
	.combout(\Mux0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~11 .lut_mask = 16'hCFA0;
defparam \Mux0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N27
dffeas \registerArray[4][31] (
	.clk(clk),
	.d(Mux372),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][31] .is_wysiwyg = "true";
defparam \registerArray[4][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N28
cycloneive_lcell_comb \Mux0~12 (
// Equation(s):
// \Mux0~12_combout  = (cuifregS_0 & (((cuifregS_1) # (\registerArray[5][31]~q )))) # (!cuifregS_0 & (\registerArray[4][31]~q  & (!cuifregS_1)))

	.dataa(cuifregS_0),
	.datab(\registerArray[4][31]~q ),
	.datac(cuifregS_1),
	.datad(\registerArray[5][31]~q ),
	.cin(gnd),
	.combout(\Mux0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~12 .lut_mask = 16'hAEA4;
defparam \Mux0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N4
cycloneive_lcell_comb \Mux0~13 (
// Equation(s):
// \Mux0~13_combout  = (cuifregS_1 & ((\Mux0~12_combout  & ((\registerArray[7][31]~q ))) # (!\Mux0~12_combout  & (\registerArray[6][31]~q )))) # (!cuifregS_1 & (\Mux0~12_combout ))

	.dataa(cuifregS_1),
	.datab(\Mux0~12_combout ),
	.datac(\registerArray[6][31]~q ),
	.datad(\registerArray[7][31]~q ),
	.cin(gnd),
	.combout(\Mux0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~13 .lut_mask = 16'hEC64;
defparam \Mux0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N14
cycloneive_lcell_comb \Mux0~14 (
// Equation(s):
// \Mux0~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][31]~q ))) # (!cuifregS_1 & (\registerArray[1][31]~q ))))

	.dataa(\registerArray[1][31]~q ),
	.datab(\registerArray[3][31]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~14 .lut_mask = 16'hC0A0;
defparam \Mux0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N28
cycloneive_lcell_comb \Mux0~15 (
// Equation(s):
// \Mux0~15_combout  = (\Mux0~14_combout ) # ((!cuifregS_0 & (\registerArray[2][31]~q  & cuifregS_1)))

	.dataa(cuifregS_0),
	.datab(\registerArray[2][31]~q ),
	.datac(\Mux0~14_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~15 .lut_mask = 16'hF4F0;
defparam \Mux0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N30
cycloneive_lcell_comb \Mux0~16 (
// Equation(s):
// \Mux0~16_combout  = (cuifregS_2 & ((cuifregS_3) # ((\Mux0~13_combout )))) # (!cuifregS_2 & (!cuifregS_3 & ((\Mux0~15_combout ))))

	.dataa(cuifregS_2),
	.datab(cuifregS_3),
	.datac(\Mux0~13_combout ),
	.datad(\Mux0~15_combout ),
	.cin(gnd),
	.combout(\Mux0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~16 .lut_mask = 16'hB9A8;
defparam \Mux0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N0
cycloneive_lcell_comb \Mux0~17 (
// Equation(s):
// \Mux0~17_combout  = (cuifregS_0 & (((\registerArray[13][31]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[12][31]~q  & ((!cuifregS_1))))

	.dataa(cuifregS_0),
	.datab(\registerArray[12][31]~q ),
	.datac(\registerArray[13][31]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~17 .lut_mask = 16'hAAE4;
defparam \Mux0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N2
cycloneive_lcell_comb \Mux0~18 (
// Equation(s):
// \Mux0~18_combout  = (cuifregS_1 & ((\Mux0~17_combout  & (\registerArray[15][31]~q )) # (!\Mux0~17_combout  & ((\registerArray[14][31]~q ))))) # (!cuifregS_1 & (((\Mux0~17_combout ))))

	.dataa(\registerArray[15][31]~q ),
	.datab(cuifregS_1),
	.datac(\registerArray[14][31]~q ),
	.datad(\Mux0~17_combout ),
	.cin(gnd),
	.combout(\Mux0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~18 .lut_mask = 16'hBBC0;
defparam \Mux0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N8
cycloneive_lcell_comb \Mux0~19 (
// Equation(s):
// \Mux0~19_combout  = (cuifregS_3 & ((\Mux0~16_combout  & ((\Mux0~18_combout ))) # (!\Mux0~16_combout  & (\Mux0~11_combout )))) # (!cuifregS_3 & (((\Mux0~16_combout ))))

	.dataa(cuifregS_3),
	.datab(\Mux0~11_combout ),
	.datac(\Mux0~16_combout ),
	.datad(\Mux0~18_combout ),
	.cin(gnd),
	.combout(\Mux0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~19 .lut_mask = 16'hF858;
defparam \Mux0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N24
cycloneive_lcell_comb \Mux0~7 (
// Equation(s):
// \Mux0~7_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[23][31]~q ))) # (!cuifregS_2 & (\registerArray[19][31]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[19][31]~q ),
	.datac(\registerArray[23][31]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~7 .lut_mask = 16'hFA44;
defparam \Mux0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N26
cycloneive_lcell_comb \Mux0~8 (
// Equation(s):
// \Mux0~8_combout  = (\Mux0~7_combout  & ((\registerArray[31][31]~q ) # ((!cuifregS_3)))) # (!\Mux0~7_combout  & (((\registerArray[27][31]~q  & cuifregS_3))))

	.dataa(\registerArray[31][31]~q ),
	.datab(\Mux0~7_combout ),
	.datac(\registerArray[27][31]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~8 .lut_mask = 16'hB8CC;
defparam \Mux0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y43_N29
dffeas \registerArray[24][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][31] .is_wysiwyg = "true";
defparam \registerArray[24][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N28
cycloneive_lcell_comb \Mux0~4 (
// Equation(s):
// \Mux0~4_combout  = (cuifregS_3 & (((\registerArray[24][31]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[16][31]~q  & ((!cuifregS_2))))

	.dataa(\registerArray[16][31]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[24][31]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~4 .lut_mask = 16'hCCE2;
defparam \Mux0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y43_N26
cycloneive_lcell_comb \Mux0~5 (
// Equation(s):
// \Mux0~5_combout  = (cuifregS_2 & ((\Mux0~4_combout  & (\registerArray[28][31]~q )) # (!\Mux0~4_combout  & ((\registerArray[20][31]~q ))))) # (!cuifregS_2 & (((\Mux0~4_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[28][31]~q ),
	.datac(\registerArray[20][31]~q ),
	.datad(\Mux0~4_combout ),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~5 .lut_mask = 16'hDDA0;
defparam \Mux0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y40_N7
dffeas \registerArray[22][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][31] .is_wysiwyg = "true";
defparam \registerArray[22][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N5
dffeas \registerArray[26][31] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux372),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][31] .is_wysiwyg = "true";
defparam \registerArray[26][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N4
cycloneive_lcell_comb \Mux0~2 (
// Equation(s):
// \Mux0~2_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & ((\registerArray[26][31]~q ))) # (!cuifregS_3 & (\registerArray[18][31]~q ))))

	.dataa(\registerArray[18][31]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[26][31]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~2 .lut_mask = 16'hFC22;
defparam \Mux0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N6
cycloneive_lcell_comb \Mux0~3 (
// Equation(s):
// \Mux0~3_combout  = (cuifregS_2 & ((\Mux0~2_combout  & (\registerArray[30][31]~q )) # (!\Mux0~2_combout  & ((\registerArray[22][31]~q ))))) # (!cuifregS_2 & (((\Mux0~2_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[30][31]~q ),
	.datac(\registerArray[22][31]~q ),
	.datad(\Mux0~2_combout ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~3 .lut_mask = 16'hDDA0;
defparam \Mux0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N18
cycloneive_lcell_comb \Mux0~6 (
// Equation(s):
// \Mux0~6_combout  = (cuifregS_0 & (cuifregS_1)) # (!cuifregS_0 & ((cuifregS_1 & ((\Mux0~3_combout ))) # (!cuifregS_1 & (\Mux0~5_combout ))))

	.dataa(cuifregS_0),
	.datab(cuifregS_1),
	.datac(\Mux0~5_combout ),
	.datad(\Mux0~3_combout ),
	.cin(gnd),
	.combout(\Mux0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~6 .lut_mask = 16'hDC98;
defparam \Mux0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N30
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// \Mux0~0_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & (\registerArray[21][31]~q )) # (!cuifregS_2 & ((\registerArray[17][31]~q )))))

	.dataa(\registerArray[21][31]~q ),
	.datab(\registerArray[17][31]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'hFA0C;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N16
cycloneive_lcell_comb \Mux0~1 (
// Equation(s):
// \Mux0~1_combout  = (\Mux0~0_combout  & ((\registerArray[29][31]~q ) # ((!cuifregS_3)))) # (!\Mux0~0_combout  & (((\registerArray[25][31]~q  & cuifregS_3))))

	.dataa(\registerArray[29][31]~q ),
	.datab(\registerArray[25][31]~q ),
	.datac(\Mux0~0_combout ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~1 .lut_mask = 16'hACF0;
defparam \Mux0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y43_N2
cycloneive_lcell_comb \Mux0~9 (
// Equation(s):
// \Mux0~9_combout  = (cuifregS_0 & ((\Mux0~6_combout  & (\Mux0~8_combout )) # (!\Mux0~6_combout  & ((\Mux0~1_combout ))))) # (!cuifregS_0 & (((\Mux0~6_combout ))))

	.dataa(cuifregS_0),
	.datab(\Mux0~8_combout ),
	.datac(\Mux0~6_combout ),
	.datad(\Mux0~1_combout ),
	.cin(gnd),
	.combout(\Mux0~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~9 .lut_mask = 16'hDAD0;
defparam \Mux0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N2
cycloneive_lcell_comb \registerArray[26][29]~feeder (
// Equation(s):
// \registerArray[26][29]~feeder_combout  = \Mux39~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux392),
	.cin(gnd),
	.combout(\registerArray[26][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[26][29]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[26][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N3
dffeas \registerArray[26][29] (
	.clk(clk),
	.d(\registerArray[26][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][29] .is_wysiwyg = "true";
defparam \registerArray[26][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N0
cycloneive_lcell_comb \Mux2~2 (
// Equation(s):
// \Mux2~2_combout  = (cuifregS_3 & (((cuifregS_2) # (\registerArray[26][29]~q )))) # (!cuifregS_3 & (\registerArray[18][29]~q  & (!cuifregS_2)))

	.dataa(\registerArray[18][29]~q ),
	.datab(cuifregS_3),
	.datac(cuifregS_2),
	.datad(\registerArray[26][29]~q ),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~2 .lut_mask = 16'hCEC2;
defparam \Mux2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N2
cycloneive_lcell_comb \Mux2~3 (
// Equation(s):
// \Mux2~3_combout  = (cuifregS_2 & ((\Mux2~2_combout  & (\registerArray[30][29]~q )) # (!\Mux2~2_combout  & ((\registerArray[22][29]~q ))))) # (!cuifregS_2 & (((\Mux2~2_combout ))))

	.dataa(\registerArray[30][29]~q ),
	.datab(\registerArray[22][29]~q ),
	.datac(cuifregS_2),
	.datad(\Mux2~2_combout ),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~3 .lut_mask = 16'hAFC0;
defparam \Mux2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N4
cycloneive_lcell_comb \Mux2~6 (
// Equation(s):
// \Mux2~6_combout  = (cuifregS_1 & (((cuifregS_0) # (\Mux2~3_combout )))) # (!cuifregS_1 & (\Mux2~5_combout  & (!cuifregS_0)))

	.dataa(\Mux2~5_combout ),
	.datab(cuifregS_1),
	.datac(cuifregS_0),
	.datad(\Mux2~3_combout ),
	.cin(gnd),
	.combout(\Mux2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~6 .lut_mask = 16'hCEC2;
defparam \Mux2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N4
cycloneive_lcell_comb \Mux2~7 (
// Equation(s):
// \Mux2~7_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[23][29]~q ))) # (!cuifregS_2 & (\registerArray[19][29]~q ))))

	.dataa(\registerArray[19][29]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[23][29]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~7 .lut_mask = 16'hFC22;
defparam \Mux2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N18
cycloneive_lcell_comb \Mux2~8 (
// Equation(s):
// \Mux2~8_combout  = (\Mux2~7_combout  & ((\registerArray[31][29]~q ) # ((!cuifregS_3)))) # (!\Mux2~7_combout  & (((\registerArray[27][29]~q  & cuifregS_3))))

	.dataa(\registerArray[31][29]~q ),
	.datab(\Mux2~7_combout ),
	.datac(\registerArray[27][29]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~8 .lut_mask = 16'hB8CC;
defparam \Mux2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N4
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// \Mux2~0_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[21][29]~q ))) # (!cuifregS_2 & (\registerArray[17][29]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[17][29]~q ),
	.datac(\registerArray[21][29]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'hFA44;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N28
cycloneive_lcell_comb \Mux2~1 (
// Equation(s):
// \Mux2~1_combout  = (cuifregS_3 & ((\Mux2~0_combout  & (\registerArray[29][29]~q )) # (!\Mux2~0_combout  & ((\registerArray[25][29]~q ))))) # (!cuifregS_3 & (((\Mux2~0_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[29][29]~q ),
	.datac(\registerArray[25][29]~q ),
	.datad(\Mux2~0_combout ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~1 .lut_mask = 16'hDDA0;
defparam \Mux2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N14
cycloneive_lcell_comb \Mux2~9 (
// Equation(s):
// \Mux2~9_combout  = (cuifregS_0 & ((\Mux2~6_combout  & (\Mux2~8_combout )) # (!\Mux2~6_combout  & ((\Mux2~1_combout ))))) # (!cuifregS_0 & (\Mux2~6_combout ))

	.dataa(cuifregS_0),
	.datab(\Mux2~6_combout ),
	.datac(\Mux2~8_combout ),
	.datad(\Mux2~1_combout ),
	.cin(gnd),
	.combout(\Mux2~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~9 .lut_mask = 16'hE6C4;
defparam \Mux2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N12
cycloneive_lcell_comb \Mux2~17 (
// Equation(s):
// \Mux2~17_combout  = (cuifregS_0 & (((\registerArray[13][29]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[12][29]~q  & ((!cuifregS_1))))

	.dataa(cuifregS_0),
	.datab(\registerArray[12][29]~q ),
	.datac(\registerArray[13][29]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux2~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~17 .lut_mask = 16'hAAE4;
defparam \Mux2~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N14
cycloneive_lcell_comb \Mux2~18 (
// Equation(s):
// \Mux2~18_combout  = (cuifregS_1 & ((\Mux2~17_combout  & (\registerArray[15][29]~q )) # (!\Mux2~17_combout  & ((\registerArray[14][29]~q ))))) # (!cuifregS_1 & (((\Mux2~17_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[15][29]~q ),
	.datac(\registerArray[14][29]~q ),
	.datad(\Mux2~17_combout ),
	.cin(gnd),
	.combout(\Mux2~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~18 .lut_mask = 16'hDDA0;
defparam \Mux2~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N30
cycloneive_lcell_comb \Mux2~14 (
// Equation(s):
// \Mux2~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][29]~q ))) # (!cuifregS_1 & (\registerArray[1][29]~q ))))

	.dataa(\registerArray[1][29]~q ),
	.datab(\registerArray[3][29]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux2~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~14 .lut_mask = 16'hC0A0;
defparam \Mux2~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N26
cycloneive_lcell_comb \Mux2~15 (
// Equation(s):
// \Mux2~15_combout  = (\Mux2~14_combout ) # ((\registerArray[2][29]~q  & (!cuifregS_0 & cuifregS_1)))

	.dataa(\registerArray[2][29]~q ),
	.datab(cuifregS_0),
	.datac(cuifregS_1),
	.datad(\Mux2~14_combout ),
	.cin(gnd),
	.combout(\Mux2~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~15 .lut_mask = 16'hFF20;
defparam \Mux2~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N3
dffeas \registerArray[5][29] (
	.clk(clk),
	.d(Mux392),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][29] .is_wysiwyg = "true";
defparam \registerArray[5][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N18
cycloneive_lcell_comb \Mux2~12 (
// Equation(s):
// \Mux2~12_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & (\registerArray[5][29]~q )) # (!cuifregS_0 & ((\registerArray[4][29]~q )))))

	.dataa(cuifregS_1),
	.datab(\registerArray[5][29]~q ),
	.datac(cuifregS_0),
	.datad(\registerArray[4][29]~q ),
	.cin(gnd),
	.combout(\Mux2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~12 .lut_mask = 16'hE5E0;
defparam \Mux2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N0
cycloneive_lcell_comb \Mux2~13 (
// Equation(s):
// \Mux2~13_combout  = (cuifregS_1 & ((\Mux2~12_combout  & (\registerArray[7][29]~q )) # (!\Mux2~12_combout  & ((\registerArray[6][29]~q ))))) # (!cuifregS_1 & (((\Mux2~12_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[7][29]~q ),
	.datac(\registerArray[6][29]~q ),
	.datad(\Mux2~12_combout ),
	.cin(gnd),
	.combout(\Mux2~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~13 .lut_mask = 16'hDDA0;
defparam \Mux2~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N8
cycloneive_lcell_comb \Mux2~16 (
// Equation(s):
// \Mux2~16_combout  = (cuifregS_2 & ((cuifregS_3) # ((\Mux2~13_combout )))) # (!cuifregS_2 & (!cuifregS_3 & (\Mux2~15_combout )))

	.dataa(cuifregS_2),
	.datab(cuifregS_3),
	.datac(\Mux2~15_combout ),
	.datad(\Mux2~13_combout ),
	.cin(gnd),
	.combout(\Mux2~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~16 .lut_mask = 16'hBA98;
defparam \Mux2~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N2
cycloneive_lcell_comb \Mux2~10 (
// Equation(s):
// \Mux2~10_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\registerArray[10][29]~q )) # (!cuifregS_1 & ((\registerArray[8][29]~q )))))

	.dataa(\registerArray[10][29]~q ),
	.datab(\registerArray[8][29]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~10 .lut_mask = 16'hFA0C;
defparam \Mux2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N20
cycloneive_lcell_comb \Mux2~11 (
// Equation(s):
// \Mux2~11_combout  = (cuifregS_0 & ((\Mux2~10_combout  & ((\registerArray[11][29]~q ))) # (!\Mux2~10_combout  & (\registerArray[9][29]~q )))) # (!cuifregS_0 & (((\Mux2~10_combout ))))

	.dataa(\registerArray[9][29]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[11][29]~q ),
	.datad(\Mux2~10_combout ),
	.cin(gnd),
	.combout(\Mux2~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~11 .lut_mask = 16'hF388;
defparam \Mux2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y37_N18
cycloneive_lcell_comb \Mux2~19 (
// Equation(s):
// \Mux2~19_combout  = (cuifregS_3 & ((\Mux2~16_combout  & (\Mux2~18_combout )) # (!\Mux2~16_combout  & ((\Mux2~11_combout ))))) # (!cuifregS_3 & (((\Mux2~16_combout ))))

	.dataa(cuifregS_3),
	.datab(\Mux2~18_combout ),
	.datac(\Mux2~16_combout ),
	.datad(\Mux2~11_combout ),
	.cin(gnd),
	.combout(\Mux2~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~19 .lut_mask = 16'hDAD0;
defparam \Mux2~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y36_N17
dffeas \registerArray[13][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][30] .is_wysiwyg = "true";
defparam \registerArray[13][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N16
cycloneive_lcell_comb \Mux1~17 (
// Equation(s):
// \Mux1~17_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & ((\registerArray[13][30]~q ))) # (!cuifregS_0 & (\registerArray[12][30]~q ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[12][30]~q ),
	.datac(\registerArray[13][30]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux1~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~17 .lut_mask = 16'hFA44;
defparam \Mux1~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N18
cycloneive_lcell_comb \Mux1~18 (
// Equation(s):
// \Mux1~18_combout  = (cuifregS_1 & ((\Mux1~17_combout  & (\registerArray[15][30]~q )) # (!\Mux1~17_combout  & ((\registerArray[14][30]~q ))))) # (!cuifregS_1 & (((\Mux1~17_combout ))))

	.dataa(\registerArray[15][30]~q ),
	.datab(cuifregS_1),
	.datac(\registerArray[14][30]~q ),
	.datad(\Mux1~17_combout ),
	.cin(gnd),
	.combout(\Mux1~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~18 .lut_mask = 16'hBBC0;
defparam \Mux1~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N28
cycloneive_lcell_comb \registerArray[5][30]~feeder (
// Equation(s):
// \registerArray[5][30]~feeder_combout  = \Mux38~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux382),
	.cin(gnd),
	.combout(\registerArray[5][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[5][30]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[5][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y31_N29
dffeas \registerArray[5][30] (
	.clk(clk),
	.d(\registerArray[5][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][30] .is_wysiwyg = "true";
defparam \registerArray[5][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N4
cycloneive_lcell_comb \Mux1~10 (
// Equation(s):
// \Mux1~10_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & ((\registerArray[5][30]~q ))) # (!cuifregS_0 & (\registerArray[4][30]~q ))))

	.dataa(\registerArray[4][30]~q ),
	.datab(\registerArray[5][30]~q ),
	.datac(cuifregS_1),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~10 .lut_mask = 16'hFC0A;
defparam \Mux1~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N30
cycloneive_lcell_comb \Mux1~11 (
// Equation(s):
// \Mux1~11_combout  = (\Mux1~10_combout  & (((\registerArray[7][30]~q ) # (!cuifregS_1)))) # (!\Mux1~10_combout  & (\registerArray[6][30]~q  & ((cuifregS_1))))

	.dataa(\registerArray[6][30]~q ),
	.datab(\registerArray[7][30]~q ),
	.datac(\Mux1~10_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux1~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~11 .lut_mask = 16'hCAF0;
defparam \Mux1~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N1
dffeas \registerArray[3][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][30] .is_wysiwyg = "true";
defparam \registerArray[3][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N0
cycloneive_lcell_comb \Mux1~14 (
// Equation(s):
// \Mux1~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][30]~q ))) # (!cuifregS_1 & (\registerArray[1][30]~q ))))

	.dataa(\registerArray[1][30]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[3][30]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux1~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~14 .lut_mask = 16'hC088;
defparam \Mux1~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N22
cycloneive_lcell_comb \Mux1~15 (
// Equation(s):
// \Mux1~15_combout  = (\Mux1~14_combout ) # ((\registerArray[2][30]~q  & (!cuifregS_0 & cuifregS_1)))

	.dataa(\registerArray[2][30]~q ),
	.datab(cuifregS_0),
	.datac(cuifregS_1),
	.datad(\Mux1~14_combout ),
	.cin(gnd),
	.combout(\Mux1~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~15 .lut_mask = 16'hFF20;
defparam \Mux1~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N12
cycloneive_lcell_comb \Mux1~13 (
// Equation(s):
// \Mux1~13_combout  = (\Mux1~12_combout  & ((\registerArray[11][30]~q ) # ((!cuifregS_0)))) # (!\Mux1~12_combout  & (((\registerArray[9][30]~q  & cuifregS_0))))

	.dataa(\Mux1~12_combout ),
	.datab(\registerArray[11][30]~q ),
	.datac(\registerArray[9][30]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux1~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~13 .lut_mask = 16'hD8AA;
defparam \Mux1~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N20
cycloneive_lcell_comb \Mux1~16 (
// Equation(s):
// \Mux1~16_combout  = (cuifregS_3 & ((cuifregS_2) # ((\Mux1~13_combout )))) # (!cuifregS_3 & (!cuifregS_2 & (\Mux1~15_combout )))

	.dataa(cuifregS_3),
	.datab(cuifregS_2),
	.datac(\Mux1~15_combout ),
	.datad(\Mux1~13_combout ),
	.cin(gnd),
	.combout(\Mux1~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~16 .lut_mask = 16'hBA98;
defparam \Mux1~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N26
cycloneive_lcell_comb \Mux1~19 (
// Equation(s):
// \Mux1~19_combout  = (cuifregS_2 & ((\Mux1~16_combout  & (\Mux1~18_combout )) # (!\Mux1~16_combout  & ((\Mux1~11_combout ))))) # (!cuifregS_2 & (((\Mux1~16_combout ))))

	.dataa(\Mux1~18_combout ),
	.datab(cuifregS_2),
	.datac(\Mux1~11_combout ),
	.datad(\Mux1~16_combout ),
	.cin(gnd),
	.combout(\Mux1~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~19 .lut_mask = 16'hBBC0;
defparam \Mux1~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N14
cycloneive_lcell_comb \registerArray[24][30]~feeder (
// Equation(s):
// \registerArray[24][30]~feeder_combout  = \Mux38~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux382),
	.cin(gnd),
	.combout(\registerArray[24][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[24][30]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[24][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y44_N15
dffeas \registerArray[24][30] (
	.clk(clk),
	.d(\registerArray[24][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][30] .is_wysiwyg = "true";
defparam \registerArray[24][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N16
cycloneive_lcell_comb \registerArray[28][30]~feeder (
// Equation(s):
// \registerArray[28][30]~feeder_combout  = \Mux38~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux382),
	.cin(gnd),
	.combout(\registerArray[28][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[28][30]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[28][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N17
dffeas \registerArray[28][30] (
	.clk(clk),
	.d(\registerArray[28][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~67_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[28][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[28][30] .is_wysiwyg = "true";
defparam \registerArray[28][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N6
cycloneive_lcell_comb \Mux1~4 (
// Equation(s):
// \Mux1~4_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & (\registerArray[20][30]~q )) # (!cuifregS_2 & ((\registerArray[16][30]~q )))))

	.dataa(cuifregS_3),
	.datab(\registerArray[20][30]~q ),
	.datac(\registerArray[16][30]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~4 .lut_mask = 16'hEE50;
defparam \Mux1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N0
cycloneive_lcell_comb \Mux1~5 (
// Equation(s):
// \Mux1~5_combout  = (cuifregS_3 & ((\Mux1~4_combout  & ((\registerArray[28][30]~q ))) # (!\Mux1~4_combout  & (\registerArray[24][30]~q )))) # (!cuifregS_3 & (((\Mux1~4_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[24][30]~q ),
	.datac(\registerArray[28][30]~q ),
	.datad(\Mux1~4_combout ),
	.cin(gnd),
	.combout(\Mux1~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~5 .lut_mask = 16'hF588;
defparam \Mux1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N30
cycloneive_lcell_comb \Mux1~6 (
// Equation(s):
// \Mux1~6_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\Mux1~3_combout )) # (!cuifregS_1 & ((\Mux1~5_combout )))))

	.dataa(\Mux1~3_combout ),
	.datab(cuifregS_0),
	.datac(cuifregS_1),
	.datad(\Mux1~5_combout ),
	.cin(gnd),
	.combout(\Mux1~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~6 .lut_mask = 16'hE3E0;
defparam \Mux1~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N16
cycloneive_lcell_comb \Mux1~7 (
// Equation(s):
// \Mux1~7_combout  = (cuifregS_3 & (((\registerArray[27][30]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[19][30]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[19][30]~q ),
	.datac(\registerArray[27][30]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux1~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~7 .lut_mask = 16'hAAE4;
defparam \Mux1~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N23
dffeas \registerArray[23][30] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux382),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][30] .is_wysiwyg = "true";
defparam \registerArray[23][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N22
cycloneive_lcell_comb \Mux1~8 (
// Equation(s):
// \Mux1~8_combout  = (\Mux1~7_combout  & ((\registerArray[31][30]~q ) # ((!cuifregS_2)))) # (!\Mux1~7_combout  & (((\registerArray[23][30]~q  & cuifregS_2))))

	.dataa(\registerArray[31][30]~q ),
	.datab(\Mux1~7_combout ),
	.datac(\registerArray[23][30]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux1~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~8 .lut_mask = 16'hB8CC;
defparam \Mux1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N2
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// \Mux1~0_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & (\registerArray[25][30]~q )) # (!cuifregS_3 & ((\registerArray[17][30]~q )))))

	.dataa(\registerArray[25][30]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[17][30]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'hEE30;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N28
cycloneive_lcell_comb \Mux1~1 (
// Equation(s):
// \Mux1~1_combout  = (cuifregS_2 & ((\Mux1~0_combout  & ((\registerArray[29][30]~q ))) # (!\Mux1~0_combout  & (\registerArray[21][30]~q )))) # (!cuifregS_2 & (((\Mux1~0_combout ))))

	.dataa(\registerArray[21][30]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[29][30]~q ),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~1 .lut_mask = 16'hF388;
defparam \Mux1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y44_N24
cycloneive_lcell_comb \Mux1~9 (
// Equation(s):
// \Mux1~9_combout  = (\Mux1~6_combout  & (((\Mux1~8_combout )) # (!cuifregS_0))) # (!\Mux1~6_combout  & (cuifregS_0 & ((\Mux1~1_combout ))))

	.dataa(\Mux1~6_combout ),
	.datab(cuifregS_0),
	.datac(\Mux1~8_combout ),
	.datad(\Mux1~1_combout ),
	.cin(gnd),
	.combout(\Mux1~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~9 .lut_mask = 16'hE6A2;
defparam \Mux1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N0
cycloneive_lcell_comb \Mux3~7 (
// Equation(s):
// \Mux3~7_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & ((\registerArray[27][28]~q ))) # (!cuifregS_3 & (\registerArray[19][28]~q ))))

	.dataa(\registerArray[19][28]~q ),
	.datab(\registerArray[27][28]~q ),
	.datac(cuifregS_2),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux3~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~7 .lut_mask = 16'hFC0A;
defparam \Mux3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N26
cycloneive_lcell_comb \Mux3~8 (
// Equation(s):
// \Mux3~8_combout  = (cuifregS_2 & ((\Mux3~7_combout  & ((\registerArray[31][28]~q ))) # (!\Mux3~7_combout  & (\registerArray[23][28]~q )))) # (!cuifregS_2 & (((\Mux3~7_combout ))))

	.dataa(\registerArray[23][28]~q ),
	.datab(\registerArray[31][28]~q ),
	.datac(cuifregS_2),
	.datad(\Mux3~7_combout ),
	.cin(gnd),
	.combout(\Mux3~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~8 .lut_mask = 16'hCFA0;
defparam \Mux3~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y40_N4
cycloneive_lcell_comb \registerArray[17][28]~feeder (
// Equation(s):
// \registerArray[17][28]~feeder_combout  = \Mux40~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux402),
	.cin(gnd),
	.combout(\registerArray[17][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[17][28]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[17][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y40_N5
dffeas \registerArray[17][28] (
	.clk(clk),
	.d(\registerArray[17][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][28] .is_wysiwyg = "true";
defparam \registerArray[17][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N28
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (cuifregS_3 & ((\registerArray[25][28]~q ) # ((cuifregS_2)))) # (!cuifregS_3 & (((!cuifregS_2 & \registerArray[17][28]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[25][28]~q ),
	.datac(cuifregS_2),
	.datad(\registerArray[17][28]~q ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hADA8;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N2
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// \Mux3~1_combout  = (cuifregS_2 & ((\Mux3~0_combout  & ((\registerArray[29][28]~q ))) # (!\Mux3~0_combout  & (\registerArray[21][28]~q )))) # (!cuifregS_2 & (((\Mux3~0_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[21][28]~q ),
	.datac(\registerArray[29][28]~q ),
	.datad(\Mux3~0_combout ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'hF588;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N7
dffeas \registerArray[24][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][28] .is_wysiwyg = "true";
defparam \registerArray[24][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N10
cycloneive_lcell_comb \registerArray[16][28]~feeder (
// Equation(s):
// \registerArray[16][28]~feeder_combout  = \Mux40~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux402),
	.cin(gnd),
	.combout(\registerArray[16][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[16][28]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[16][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y34_N11
dffeas \registerArray[16][28] (
	.clk(clk),
	.d(\registerArray[16][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][28] .is_wysiwyg = "true";
defparam \registerArray[16][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N20
cycloneive_lcell_comb \Mux3~4 (
// Equation(s):
// \Mux3~4_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[20][28]~q ))) # (!cuifregS_2 & (\registerArray[16][28]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[16][28]~q ),
	.datac(\registerArray[20][28]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~4 .lut_mask = 16'hFA44;
defparam \Mux3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N6
cycloneive_lcell_comb \Mux3~5 (
// Equation(s):
// \Mux3~5_combout  = (cuifregS_3 & ((\Mux3~4_combout  & (\registerArray[28][28]~q )) # (!\Mux3~4_combout  & ((\registerArray[24][28]~q ))))) # (!cuifregS_3 & (((\Mux3~4_combout ))))

	.dataa(\registerArray[28][28]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[24][28]~q ),
	.datad(\Mux3~4_combout ),
	.cin(gnd),
	.combout(\Mux3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~5 .lut_mask = 16'hBBC0;
defparam \Mux3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N13
dffeas \registerArray[22][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][28] .is_wysiwyg = "true";
defparam \registerArray[22][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N12
cycloneive_lcell_comb \Mux3~2 (
// Equation(s):
// \Mux3~2_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[22][28]~q ))) # (!cuifregS_2 & (\registerArray[18][28]~q ))))

	.dataa(\registerArray[18][28]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[22][28]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~2 .lut_mask = 16'hFC22;
defparam \Mux3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N22
cycloneive_lcell_comb \Mux3~3 (
// Equation(s):
// \Mux3~3_combout  = (cuifregS_3 & ((\Mux3~2_combout  & (\registerArray[30][28]~q )) # (!\Mux3~2_combout  & ((\registerArray[26][28]~q ))))) # (!cuifregS_3 & (((\Mux3~2_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[30][28]~q ),
	.datac(\registerArray[26][28]~q ),
	.datad(\Mux3~2_combout ),
	.cin(gnd),
	.combout(\Mux3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~3 .lut_mask = 16'hDDA0;
defparam \Mux3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N0
cycloneive_lcell_comb \Mux3~6 (
// Equation(s):
// \Mux3~6_combout  = (cuifregS_1 & ((cuifregS_0) # ((\Mux3~3_combout )))) # (!cuifregS_1 & (!cuifregS_0 & (\Mux3~5_combout )))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\Mux3~5_combout ),
	.datad(\Mux3~3_combout ),
	.cin(gnd),
	.combout(\Mux3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~6 .lut_mask = 16'hBA98;
defparam \Mux3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N22
cycloneive_lcell_comb \Mux3~9 (
// Equation(s):
// \Mux3~9_combout  = (cuifregS_0 & ((\Mux3~6_combout  & (\Mux3~8_combout )) # (!\Mux3~6_combout  & ((\Mux3~1_combout ))))) # (!cuifregS_0 & (((\Mux3~6_combout ))))

	.dataa(cuifregS_0),
	.datab(\Mux3~8_combout ),
	.datac(\Mux3~1_combout ),
	.datad(\Mux3~6_combout ),
	.cin(gnd),
	.combout(\Mux3~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~9 .lut_mask = 16'hDDA0;
defparam \Mux3~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N20
cycloneive_lcell_comb \Mux3~17 (
// Equation(s):
// \Mux3~17_combout  = (cuifregS_0 & (((\registerArray[13][28]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[12][28]~q  & ((!cuifregS_1))))

	.dataa(cuifregS_0),
	.datab(\registerArray[12][28]~q ),
	.datac(\registerArray[13][28]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux3~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~17 .lut_mask = 16'hAAE4;
defparam \Mux3~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N10
cycloneive_lcell_comb \Mux3~18 (
// Equation(s):
// \Mux3~18_combout  = (cuifregS_1 & ((\Mux3~17_combout  & (\registerArray[15][28]~q )) # (!\Mux3~17_combout  & ((\registerArray[14][28]~q ))))) # (!cuifregS_1 & (((\Mux3~17_combout ))))

	.dataa(\registerArray[15][28]~q ),
	.datab(cuifregS_1),
	.datac(\registerArray[14][28]~q ),
	.datad(\Mux3~17_combout ),
	.cin(gnd),
	.combout(\Mux3~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~18 .lut_mask = 16'hBBC0;
defparam \Mux3~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N21
dffeas \registerArray[6][28] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux402),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][28] .is_wysiwyg = "true";
defparam \registerArray[6][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N16
cycloneive_lcell_comb \Mux3~10 (
// Equation(s):
// \Mux3~10_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & (\registerArray[5][28]~q )) # (!cuifregS_0 & ((\registerArray[4][28]~q )))))

	.dataa(\registerArray[5][28]~q ),
	.datab(\registerArray[4][28]~q ),
	.datac(cuifregS_1),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux3~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~10 .lut_mask = 16'hFA0C;
defparam \Mux3~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N20
cycloneive_lcell_comb \Mux3~11 (
// Equation(s):
// \Mux3~11_combout  = (cuifregS_1 & ((\Mux3~10_combout  & (\registerArray[7][28]~q )) # (!\Mux3~10_combout  & ((\registerArray[6][28]~q ))))) # (!cuifregS_1 & (((\Mux3~10_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[7][28]~q ),
	.datac(\registerArray[6][28]~q ),
	.datad(\Mux3~10_combout ),
	.cin(gnd),
	.combout(\Mux3~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~11 .lut_mask = 16'hDDA0;
defparam \Mux3~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N28
cycloneive_lcell_comb \Mux3~14 (
// Equation(s):
// \Mux3~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][28]~q ))) # (!cuifregS_1 & (\registerArray[1][28]~q ))))

	.dataa(\registerArray[1][28]~q ),
	.datab(\registerArray[3][28]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux3~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~14 .lut_mask = 16'hC0A0;
defparam \Mux3~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N16
cycloneive_lcell_comb \Mux3~15 (
// Equation(s):
// \Mux3~15_combout  = (\Mux3~14_combout ) # ((cuifregS_1 & (!cuifregS_0 & \registerArray[2][28]~q )))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\registerArray[2][28]~q ),
	.datad(\Mux3~14_combout ),
	.cin(gnd),
	.combout(\Mux3~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~15 .lut_mask = 16'hFF20;
defparam \Mux3~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N2
cycloneive_lcell_comb \Mux3~12 (
// Equation(s):
// \Mux3~12_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][28]~q ))) # (!cuifregS_1 & (\registerArray[8][28]~q ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[8][28]~q ),
	.datac(\registerArray[10][28]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux3~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~12 .lut_mask = 16'hFA44;
defparam \Mux3~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N12
cycloneive_lcell_comb \Mux3~13 (
// Equation(s):
// \Mux3~13_combout  = (cuifregS_0 & ((\Mux3~12_combout  & (\registerArray[11][28]~q )) # (!\Mux3~12_combout  & ((\registerArray[9][28]~q ))))) # (!cuifregS_0 & (((\Mux3~12_combout ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[11][28]~q ),
	.datac(\registerArray[9][28]~q ),
	.datad(\Mux3~12_combout ),
	.cin(gnd),
	.combout(\Mux3~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~13 .lut_mask = 16'hDDA0;
defparam \Mux3~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N18
cycloneive_lcell_comb \Mux3~16 (
// Equation(s):
// \Mux3~16_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & ((\Mux3~13_combout ))) # (!cuifregS_3 & (\Mux3~15_combout ))))

	.dataa(cuifregS_2),
	.datab(\Mux3~15_combout ),
	.datac(cuifregS_3),
	.datad(\Mux3~13_combout ),
	.cin(gnd),
	.combout(\Mux3~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~16 .lut_mask = 16'hF4A4;
defparam \Mux3~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N20
cycloneive_lcell_comb \Mux3~19 (
// Equation(s):
// \Mux3~19_combout  = (cuifregS_2 & ((\Mux3~16_combout  & (\Mux3~18_combout )) # (!\Mux3~16_combout  & ((\Mux3~11_combout ))))) # (!cuifregS_2 & (((\Mux3~16_combout ))))

	.dataa(cuifregS_2),
	.datab(\Mux3~18_combout ),
	.datac(\Mux3~11_combout ),
	.datad(\Mux3~16_combout ),
	.cin(gnd),
	.combout(\Mux3~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~19 .lut_mask = 16'hDDA0;
defparam \Mux3~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N10
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// \Mux4~0_combout  = (cuifregS_2 & ((\registerArray[21][27]~q ) # ((cuifregS_3)))) # (!cuifregS_2 & (((\registerArray[17][27]~q  & !cuifregS_3))))

	.dataa(\registerArray[21][27]~q ),
	.datab(\registerArray[17][27]~q ),
	.datac(cuifregS_2),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'hF0AC;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N20
cycloneive_lcell_comb \Mux4~1 (
// Equation(s):
// \Mux4~1_combout  = (cuifregS_3 & ((\Mux4~0_combout  & (\registerArray[29][27]~q )) # (!\Mux4~0_combout  & ((\registerArray[25][27]~q ))))) # (!cuifregS_3 & (((\Mux4~0_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[29][27]~q ),
	.datac(\registerArray[25][27]~q ),
	.datad(\Mux4~0_combout ),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~1 .lut_mask = 16'hDDA0;
defparam \Mux4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N6
cycloneive_lcell_comb \Mux4~7 (
// Equation(s):
// \Mux4~7_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[23][27]~q ))) # (!cuifregS_2 & (\registerArray[19][27]~q ))))

	.dataa(\registerArray[19][27]~q ),
	.datab(\registerArray[23][27]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux4~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~7 .lut_mask = 16'hFC0A;
defparam \Mux4~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N16
cycloneive_lcell_comb \Mux4~8 (
// Equation(s):
// \Mux4~8_combout  = (cuifregS_3 & ((\Mux4~7_combout  & (\registerArray[31][27]~q )) # (!\Mux4~7_combout  & ((\registerArray[27][27]~q ))))) # (!cuifregS_3 & (((\Mux4~7_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[31][27]~q ),
	.datac(\registerArray[27][27]~q ),
	.datad(\Mux4~7_combout ),
	.cin(gnd),
	.combout(\Mux4~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~8 .lut_mask = 16'hDDA0;
defparam \Mux4~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N31
dffeas \registerArray[22][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][27] .is_wysiwyg = "true";
defparam \registerArray[22][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y42_N29
dffeas \registerArray[26][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][27] .is_wysiwyg = "true";
defparam \registerArray[26][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N28
cycloneive_lcell_comb \Mux4~2 (
// Equation(s):
// \Mux4~2_combout  = (cuifregS_3 & (((\registerArray[26][27]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[18][27]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[18][27]~q ),
	.datac(\registerArray[26][27]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~2 .lut_mask = 16'hAAE4;
defparam \Mux4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N30
cycloneive_lcell_comb \Mux4~3 (
// Equation(s):
// \Mux4~3_combout  = (cuifregS_2 & ((\Mux4~2_combout  & (\registerArray[30][27]~q )) # (!\Mux4~2_combout  & ((\registerArray[22][27]~q ))))) # (!cuifregS_2 & (((\Mux4~2_combout ))))

	.dataa(\registerArray[30][27]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[22][27]~q ),
	.datad(\Mux4~2_combout ),
	.cin(gnd),
	.combout(\Mux4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~3 .lut_mask = 16'hBBC0;
defparam \Mux4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N19
dffeas \registerArray[20][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][27] .is_wysiwyg = "true";
defparam \registerArray[20][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N20
cycloneive_lcell_comb \Mux4~4 (
// Equation(s):
// \Mux4~4_combout  = (cuifregS_3 & (((\registerArray[24][27]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[16][27]~q  & ((!cuifregS_2))))

	.dataa(\registerArray[16][27]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[24][27]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~4 .lut_mask = 16'hCCE2;
defparam \Mux4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N18
cycloneive_lcell_comb \Mux4~5 (
// Equation(s):
// \Mux4~5_combout  = (cuifregS_2 & ((\Mux4~4_combout  & (\registerArray[28][27]~q )) # (!\Mux4~4_combout  & ((\registerArray[20][27]~q ))))) # (!cuifregS_2 & (((\Mux4~4_combout ))))

	.dataa(\registerArray[28][27]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[20][27]~q ),
	.datad(\Mux4~4_combout ),
	.cin(gnd),
	.combout(\Mux4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~5 .lut_mask = 16'hBBC0;
defparam \Mux4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N18
cycloneive_lcell_comb \Mux4~6 (
// Equation(s):
// \Mux4~6_combout  = (cuifregS_0 & (cuifregS_1)) # (!cuifregS_0 & ((cuifregS_1 & (\Mux4~3_combout )) # (!cuifregS_1 & ((\Mux4~5_combout )))))

	.dataa(cuifregS_0),
	.datab(cuifregS_1),
	.datac(\Mux4~3_combout ),
	.datad(\Mux4~5_combout ),
	.cin(gnd),
	.combout(\Mux4~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~6 .lut_mask = 16'hD9C8;
defparam \Mux4~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N12
cycloneive_lcell_comb \Mux4~9 (
// Equation(s):
// \Mux4~9_combout  = (cuifregS_0 & ((\Mux4~6_combout  & ((\Mux4~8_combout ))) # (!\Mux4~6_combout  & (\Mux4~1_combout )))) # (!cuifregS_0 & (((\Mux4~6_combout ))))

	.dataa(\Mux4~1_combout ),
	.datab(cuifregS_0),
	.datac(\Mux4~8_combout ),
	.datad(\Mux4~6_combout ),
	.cin(gnd),
	.combout(\Mux4~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~9 .lut_mask = 16'hF388;
defparam \Mux4~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N24
cycloneive_lcell_comb \Mux4~17 (
// Equation(s):
// \Mux4~17_combout  = (cuifregS_0 & (((\registerArray[13][27]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[12][27]~q  & ((!cuifregS_1))))

	.dataa(cuifregS_0),
	.datab(\registerArray[12][27]~q ),
	.datac(\registerArray[13][27]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux4~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~17 .lut_mask = 16'hAAE4;
defparam \Mux4~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N30
cycloneive_lcell_comb \Mux4~18 (
// Equation(s):
// \Mux4~18_combout  = (cuifregS_1 & ((\Mux4~17_combout  & (\registerArray[15][27]~q )) # (!\Mux4~17_combout  & ((\registerArray[14][27]~q ))))) # (!cuifregS_1 & (((\Mux4~17_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[15][27]~q ),
	.datac(\registerArray[14][27]~q ),
	.datad(\Mux4~17_combout ),
	.cin(gnd),
	.combout(\Mux4~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~18 .lut_mask = 16'hDDA0;
defparam \Mux4~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N6
cycloneive_lcell_comb \Mux4~12 (
// Equation(s):
// \Mux4~12_combout  = (cuifregS_0 & (((\registerArray[5][27]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[4][27]~q  & ((!cuifregS_1))))

	.dataa(cuifregS_0),
	.datab(\registerArray[4][27]~q ),
	.datac(\registerArray[5][27]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux4~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~12 .lut_mask = 16'hAAE4;
defparam \Mux4~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N10
cycloneive_lcell_comb \Mux4~13 (
// Equation(s):
// \Mux4~13_combout  = (cuifregS_1 & ((\Mux4~12_combout  & (\registerArray[7][27]~q )) # (!\Mux4~12_combout  & ((\registerArray[6][27]~q ))))) # (!cuifregS_1 & (((\Mux4~12_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[7][27]~q ),
	.datac(\registerArray[6][27]~q ),
	.datad(\Mux4~12_combout ),
	.cin(gnd),
	.combout(\Mux4~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~13 .lut_mask = 16'hDDA0;
defparam \Mux4~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N22
cycloneive_lcell_comb \Mux4~14 (
// Equation(s):
// \Mux4~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][27]~q ))) # (!cuifregS_1 & (\registerArray[1][27]~q ))))

	.dataa(\registerArray[1][27]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[3][27]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux4~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~14 .lut_mask = 16'hC088;
defparam \Mux4~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N18
cycloneive_lcell_comb \Mux4~15 (
// Equation(s):
// \Mux4~15_combout  = (\Mux4~14_combout ) # ((\registerArray[2][27]~q  & (!cuifregS_0 & cuifregS_1)))

	.dataa(\registerArray[2][27]~q ),
	.datab(cuifregS_0),
	.datac(cuifregS_1),
	.datad(\Mux4~14_combout ),
	.cin(gnd),
	.combout(\Mux4~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~15 .lut_mask = 16'hFF20;
defparam \Mux4~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N8
cycloneive_lcell_comb \Mux4~16 (
// Equation(s):
// \Mux4~16_combout  = (cuifregS_2 & ((cuifregS_3) # ((\Mux4~13_combout )))) # (!cuifregS_2 & (!cuifregS_3 & ((\Mux4~15_combout ))))

	.dataa(cuifregS_2),
	.datab(cuifregS_3),
	.datac(\Mux4~13_combout ),
	.datad(\Mux4~15_combout ),
	.cin(gnd),
	.combout(\Mux4~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~16 .lut_mask = 16'hB9A8;
defparam \Mux4~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N11
dffeas \registerArray[10][27] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux412),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][27] .is_wysiwyg = "true";
defparam \registerArray[10][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N10
cycloneive_lcell_comb \Mux4~10 (
// Equation(s):
// \Mux4~10_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][27]~q ))) # (!cuifregS_1 & (\registerArray[8][27]~q ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[8][27]~q ),
	.datac(\registerArray[10][27]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux4~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~10 .lut_mask = 16'hFA44;
defparam \Mux4~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N24
cycloneive_lcell_comb \Mux4~11 (
// Equation(s):
// \Mux4~11_combout  = (cuifregS_0 & ((\Mux4~10_combout  & (\registerArray[11][27]~q )) # (!\Mux4~10_combout  & ((\registerArray[9][27]~q ))))) # (!cuifregS_0 & (((\Mux4~10_combout ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[11][27]~q ),
	.datac(\registerArray[9][27]~q ),
	.datad(\Mux4~10_combout ),
	.cin(gnd),
	.combout(\Mux4~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~11 .lut_mask = 16'hDDA0;
defparam \Mux4~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N2
cycloneive_lcell_comb \Mux4~19 (
// Equation(s):
// \Mux4~19_combout  = (cuifregS_3 & ((\Mux4~16_combout  & (\Mux4~18_combout )) # (!\Mux4~16_combout  & ((\Mux4~11_combout ))))) # (!cuifregS_3 & (((\Mux4~16_combout ))))

	.dataa(\Mux4~18_combout ),
	.datab(cuifregS_3),
	.datac(\Mux4~16_combout ),
	.datad(\Mux4~11_combout ),
	.cin(gnd),
	.combout(\Mux4~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~19 .lut_mask = 16'hBCB0;
defparam \Mux4~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N20
cycloneive_lcell_comb \Mux5~10 (
// Equation(s):
// \Mux5~10_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & (\registerArray[5][26]~q )) # (!cuifregS_0 & ((\registerArray[4][26]~q )))))

	.dataa(\registerArray[5][26]~q ),
	.datab(cuifregS_1),
	.datac(cuifregS_0),
	.datad(\registerArray[4][26]~q ),
	.cin(gnd),
	.combout(\Mux5~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~10 .lut_mask = 16'hE3E0;
defparam \Mux5~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N14
cycloneive_lcell_comb \Mux5~11 (
// Equation(s):
// \Mux5~11_combout  = (cuifregS_1 & ((\Mux5~10_combout  & (\registerArray[7][26]~q )) # (!\Mux5~10_combout  & ((\registerArray[6][26]~q ))))) # (!cuifregS_1 & (((\Mux5~10_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[7][26]~q ),
	.datac(\registerArray[6][26]~q ),
	.datad(\Mux5~10_combout ),
	.cin(gnd),
	.combout(\Mux5~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~11 .lut_mask = 16'hDDA0;
defparam \Mux5~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y38_N22
cycloneive_lcell_comb \Mux5~14 (
// Equation(s):
// \Mux5~14_combout  = (cuifregS_0 & ((cuifregS_1 & (\registerArray[3][26]~q )) # (!cuifregS_1 & ((\registerArray[1][26]~q )))))

	.dataa(\registerArray[3][26]~q ),
	.datab(\registerArray[1][26]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux5~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~14 .lut_mask = 16'hA0C0;
defparam \Mux5~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N8
cycloneive_lcell_comb \Mux5~15 (
// Equation(s):
// \Mux5~15_combout  = (\Mux5~14_combout ) # ((cuifregS_1 & (!cuifregS_0 & \registerArray[2][26]~q )))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\registerArray[2][26]~q ),
	.datad(\Mux5~14_combout ),
	.cin(gnd),
	.combout(\Mux5~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~15 .lut_mask = 16'hFF20;
defparam \Mux5~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N16
cycloneive_lcell_comb \Mux5~12 (
// Equation(s):
// \Mux5~12_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\registerArray[10][26]~q )) # (!cuifregS_1 & ((\registerArray[8][26]~q )))))

	.dataa(cuifregS_0),
	.datab(\registerArray[10][26]~q ),
	.datac(\registerArray[8][26]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux5~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~12 .lut_mask = 16'hEE50;
defparam \Mux5~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N20
cycloneive_lcell_comb \Mux5~13 (
// Equation(s):
// \Mux5~13_combout  = (cuifregS_0 & ((\Mux5~12_combout  & ((\registerArray[11][26]~q ))) # (!\Mux5~12_combout  & (\registerArray[9][26]~q )))) # (!cuifregS_0 & (((\Mux5~12_combout ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[9][26]~q ),
	.datac(\registerArray[11][26]~q ),
	.datad(\Mux5~12_combout ),
	.cin(gnd),
	.combout(\Mux5~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~13 .lut_mask = 16'hF588;
defparam \Mux5~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N26
cycloneive_lcell_comb \Mux5~16 (
// Equation(s):
// \Mux5~16_combout  = (cuifregS_2 & (cuifregS_3)) # (!cuifregS_2 & ((cuifregS_3 & ((\Mux5~13_combout ))) # (!cuifregS_3 & (\Mux5~15_combout ))))

	.dataa(cuifregS_2),
	.datab(cuifregS_3),
	.datac(\Mux5~15_combout ),
	.datad(\Mux5~13_combout ),
	.cin(gnd),
	.combout(\Mux5~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~16 .lut_mask = 16'hDC98;
defparam \Mux5~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N24
cycloneive_lcell_comb \Mux5~17 (
// Equation(s):
// \Mux5~17_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & ((\registerArray[13][26]~q ))) # (!cuifregS_0 & (\registerArray[12][26]~q ))))

	.dataa(\registerArray[12][26]~q ),
	.datab(\registerArray[13][26]~q ),
	.datac(cuifregS_1),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux5~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~17 .lut_mask = 16'hFC0A;
defparam \Mux5~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N26
cycloneive_lcell_comb \Mux5~18 (
// Equation(s):
// \Mux5~18_combout  = (cuifregS_1 & ((\Mux5~17_combout  & ((\registerArray[15][26]~q ))) # (!\Mux5~17_combout  & (\registerArray[14][26]~q )))) # (!cuifregS_1 & (((\Mux5~17_combout ))))

	.dataa(\registerArray[14][26]~q ),
	.datab(\registerArray[15][26]~q ),
	.datac(cuifregS_1),
	.datad(\Mux5~17_combout ),
	.cin(gnd),
	.combout(\Mux5~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~18 .lut_mask = 16'hCFA0;
defparam \Mux5~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N4
cycloneive_lcell_comb \Mux5~19 (
// Equation(s):
// \Mux5~19_combout  = (cuifregS_2 & ((\Mux5~16_combout  & ((\Mux5~18_combout ))) # (!\Mux5~16_combout  & (\Mux5~11_combout )))) # (!cuifregS_2 & (((\Mux5~16_combout ))))

	.dataa(cuifregS_2),
	.datab(\Mux5~11_combout ),
	.datac(\Mux5~16_combout ),
	.datad(\Mux5~18_combout ),
	.cin(gnd),
	.combout(\Mux5~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~19 .lut_mask = 16'hF858;
defparam \Mux5~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N20
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// \Mux5~0_combout  = (cuifregS_3 & (((\registerArray[25][26]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[17][26]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[17][26]~q ),
	.datac(\registerArray[25][26]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'hAAE4;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N18
cycloneive_lcell_comb \Mux5~1 (
// Equation(s):
// \Mux5~1_combout  = (cuifregS_2 & ((\Mux5~0_combout  & (\registerArray[29][26]~q )) # (!\Mux5~0_combout  & ((\registerArray[21][26]~q ))))) # (!cuifregS_2 & (((\Mux5~0_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[29][26]~q ),
	.datac(\registerArray[21][26]~q ),
	.datad(\Mux5~0_combout ),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~1 .lut_mask = 16'hDDA0;
defparam \Mux5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N28
cycloneive_lcell_comb \Mux5~7 (
// Equation(s):
// \Mux5~7_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & (\registerArray[27][26]~q )) # (!cuifregS_3 & ((\registerArray[19][26]~q )))))

	.dataa(\registerArray[27][26]~q ),
	.datab(\registerArray[19][26]~q ),
	.datac(cuifregS_2),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux5~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~7 .lut_mask = 16'hFA0C;
defparam \Mux5~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y37_N22
cycloneive_lcell_comb \Mux5~8 (
// Equation(s):
// \Mux5~8_combout  = (cuifregS_2 & ((\Mux5~7_combout  & ((\registerArray[31][26]~q ))) # (!\Mux5~7_combout  & (\registerArray[23][26]~q )))) # (!cuifregS_2 & (((\Mux5~7_combout ))))

	.dataa(\registerArray[23][26]~q ),
	.datab(\registerArray[31][26]~q ),
	.datac(cuifregS_2),
	.datad(\Mux5~7_combout ),
	.cin(gnd),
	.combout(\Mux5~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~8 .lut_mask = 16'hCFA0;
defparam \Mux5~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N16
cycloneive_lcell_comb \Mux5~2 (
// Equation(s):
// \Mux5~2_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[22][26]~q ))) # (!cuifregS_2 & (\registerArray[18][26]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[18][26]~q ),
	.datac(\registerArray[22][26]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~2 .lut_mask = 16'hFA44;
defparam \Mux5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N6
cycloneive_lcell_comb \Mux5~3 (
// Equation(s):
// \Mux5~3_combout  = (cuifregS_3 & ((\Mux5~2_combout  & (\registerArray[30][26]~q )) # (!\Mux5~2_combout  & ((\registerArray[26][26]~q ))))) # (!cuifregS_3 & (((\Mux5~2_combout ))))

	.dataa(\registerArray[30][26]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[26][26]~q ),
	.datad(\Mux5~2_combout ),
	.cin(gnd),
	.combout(\Mux5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~3 .lut_mask = 16'hBBC0;
defparam \Mux5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N28
cycloneive_lcell_comb \registerArray[20][26]~feeder (
// Equation(s):
// \registerArray[20][26]~feeder_combout  = \Mux42~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux422),
	.cin(gnd),
	.combout(\registerArray[20][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[20][26]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[20][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N29
dffeas \registerArray[20][26] (
	.clk(clk),
	.d(\registerArray[20][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][26] .is_wysiwyg = "true";
defparam \registerArray[20][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N2
cycloneive_lcell_comb \Mux5~4 (
// Equation(s):
// \Mux5~4_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[20][26]~q ))) # (!cuifregS_2 & (\registerArray[16][26]~q ))))

	.dataa(\registerArray[16][26]~q ),
	.datab(\registerArray[20][26]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~4 .lut_mask = 16'hFC0A;
defparam \Mux5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N28
cycloneive_lcell_comb \Mux5~5 (
// Equation(s):
// \Mux5~5_combout  = (cuifregS_3 & ((\Mux5~4_combout  & ((\registerArray[28][26]~q ))) # (!\Mux5~4_combout  & (\registerArray[24][26]~q )))) # (!cuifregS_3 & (((\Mux5~4_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[24][26]~q ),
	.datac(\registerArray[28][26]~q ),
	.datad(\Mux5~4_combout ),
	.cin(gnd),
	.combout(\Mux5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~5 .lut_mask = 16'hF588;
defparam \Mux5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N12
cycloneive_lcell_comb \Mux5~6 (
// Equation(s):
// \Mux5~6_combout  = (cuifregS_1 & ((cuifregS_0) # ((\Mux5~3_combout )))) # (!cuifregS_1 & (!cuifregS_0 & ((\Mux5~5_combout ))))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\Mux5~3_combout ),
	.datad(\Mux5~5_combout ),
	.cin(gnd),
	.combout(\Mux5~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~6 .lut_mask = 16'hB9A8;
defparam \Mux5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y38_N6
cycloneive_lcell_comb \Mux5~9 (
// Equation(s):
// \Mux5~9_combout  = (cuifregS_0 & ((\Mux5~6_combout  & ((\Mux5~8_combout ))) # (!\Mux5~6_combout  & (\Mux5~1_combout )))) # (!cuifregS_0 & (((\Mux5~6_combout ))))

	.dataa(\Mux5~1_combout ),
	.datab(cuifregS_0),
	.datac(\Mux5~8_combout ),
	.datad(\Mux5~6_combout ),
	.cin(gnd),
	.combout(\Mux5~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~9 .lut_mask = 16'hF388;
defparam \Mux5~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N15
dffeas \registerArray[27][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][25] .is_wysiwyg = "true";
defparam \registerArray[27][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N24
cycloneive_lcell_comb \Mux6~7 (
// Equation(s):
// \Mux6~7_combout  = (cuifregS_2 & (((\registerArray[23][25]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[19][25]~q  & ((!cuifregS_3))))

	.dataa(\registerArray[19][25]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[23][25]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux6~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~7 .lut_mask = 16'hCCE2;
defparam \Mux6~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N14
cycloneive_lcell_comb \Mux6~8 (
// Equation(s):
// \Mux6~8_combout  = (cuifregS_3 & ((\Mux6~7_combout  & (\registerArray[31][25]~q )) # (!\Mux6~7_combout  & ((\registerArray[27][25]~q ))))) # (!cuifregS_3 & (((\Mux6~7_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[31][25]~q ),
	.datac(\registerArray[27][25]~q ),
	.datad(\Mux6~7_combout ),
	.cin(gnd),
	.combout(\Mux6~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~8 .lut_mask = 16'hDDA0;
defparam \Mux6~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N22
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// \Mux6~0_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[21][25]~q ))) # (!cuifregS_2 & (\registerArray[17][25]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[17][25]~q ),
	.datac(\registerArray[21][25]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'hFA44;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N30
cycloneive_lcell_comb \Mux6~1 (
// Equation(s):
// \Mux6~1_combout  = (cuifregS_3 & ((\Mux6~0_combout  & ((\registerArray[29][25]~q ))) # (!\Mux6~0_combout  & (\registerArray[25][25]~q )))) # (!cuifregS_3 & (((\Mux6~0_combout ))))

	.dataa(\registerArray[25][25]~q ),
	.datab(\registerArray[29][25]~q ),
	.datac(cuifregS_3),
	.datad(\Mux6~0_combout ),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~1 .lut_mask = 16'hCFA0;
defparam \Mux6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N27
dffeas \registerArray[24][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][25] .is_wysiwyg = "true";
defparam \registerArray[24][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N26
cycloneive_lcell_comb \Mux6~4 (
// Equation(s):
// \Mux6~4_combout  = (cuifregS_3 & (((\registerArray[24][25]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[16][25]~q  & ((!cuifregS_2))))

	.dataa(\registerArray[16][25]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[24][25]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux6~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~4 .lut_mask = 16'hCCE2;
defparam \Mux6~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N14
cycloneive_lcell_comb \Mux6~5 (
// Equation(s):
// \Mux6~5_combout  = (cuifregS_2 & ((\Mux6~4_combout  & (\registerArray[28][25]~q )) # (!\Mux6~4_combout  & ((\registerArray[20][25]~q ))))) # (!cuifregS_2 & (((\Mux6~4_combout ))))

	.dataa(\registerArray[28][25]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[20][25]~q ),
	.datad(\Mux6~4_combout ),
	.cin(gnd),
	.combout(\Mux6~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~5 .lut_mask = 16'hBBC0;
defparam \Mux6~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N20
cycloneive_lcell_comb \Mux6~6 (
// Equation(s):
// \Mux6~6_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\Mux6~3_combout )) # (!cuifregS_1 & ((\Mux6~5_combout )))))

	.dataa(\Mux6~3_combout ),
	.datab(cuifregS_0),
	.datac(cuifregS_1),
	.datad(\Mux6~5_combout ),
	.cin(gnd),
	.combout(\Mux6~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~6 .lut_mask = 16'hE3E0;
defparam \Mux6~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N22
cycloneive_lcell_comb \Mux6~9 (
// Equation(s):
// \Mux6~9_combout  = (cuifregS_0 & ((\Mux6~6_combout  & (\Mux6~8_combout )) # (!\Mux6~6_combout  & ((\Mux6~1_combout ))))) # (!cuifregS_0 & (((\Mux6~6_combout ))))

	.dataa(\Mux6~8_combout ),
	.datab(cuifregS_0),
	.datac(\Mux6~1_combout ),
	.datad(\Mux6~6_combout ),
	.cin(gnd),
	.combout(\Mux6~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~9 .lut_mask = 16'hBBC0;
defparam \Mux6~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y43_N21
dffeas \registerArray[9][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][25] .is_wysiwyg = "true";
defparam \registerArray[9][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y43_N11
dffeas \registerArray[10][25] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux432),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][25] .is_wysiwyg = "true";
defparam \registerArray[10][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N10
cycloneive_lcell_comb \Mux6~10 (
// Equation(s):
// \Mux6~10_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][25]~q ))) # (!cuifregS_1 & (\registerArray[8][25]~q ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[8][25]~q ),
	.datac(\registerArray[10][25]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux6~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~10 .lut_mask = 16'hFA44;
defparam \Mux6~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N20
cycloneive_lcell_comb \Mux6~11 (
// Equation(s):
// \Mux6~11_combout  = (cuifregS_0 & ((\Mux6~10_combout  & (\registerArray[11][25]~q )) # (!\Mux6~10_combout  & ((\registerArray[9][25]~q ))))) # (!cuifregS_0 & (((\Mux6~10_combout ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[11][25]~q ),
	.datac(\registerArray[9][25]~q ),
	.datad(\Mux6~10_combout ),
	.cin(gnd),
	.combout(\Mux6~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~11 .lut_mask = 16'hDDA0;
defparam \Mux6~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N2
cycloneive_lcell_comb \Mux6~17 (
// Equation(s):
// \Mux6~17_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & ((\registerArray[13][25]~q ))) # (!cuifregS_0 & (\registerArray[12][25]~q ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[12][25]~q ),
	.datac(\registerArray[13][25]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux6~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~17 .lut_mask = 16'hFA44;
defparam \Mux6~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N22
cycloneive_lcell_comb \Mux6~18 (
// Equation(s):
// \Mux6~18_combout  = (\Mux6~17_combout  & ((\registerArray[15][25]~q ) # ((!cuifregS_1)))) # (!\Mux6~17_combout  & (((\registerArray[14][25]~q  & cuifregS_1))))

	.dataa(\registerArray[15][25]~q ),
	.datab(\Mux6~17_combout ),
	.datac(\registerArray[14][25]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux6~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~18 .lut_mask = 16'hB8CC;
defparam \Mux6~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N24
cycloneive_lcell_comb \Mux6~14 (
// Equation(s):
// \Mux6~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][25]~q ))) # (!cuifregS_1 & (\registerArray[1][25]~q ))))

	.dataa(\registerArray[1][25]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[3][25]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux6~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~14 .lut_mask = 16'hC088;
defparam \Mux6~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N4
cycloneive_lcell_comb \Mux6~15 (
// Equation(s):
// \Mux6~15_combout  = (\Mux6~14_combout ) # ((\registerArray[2][25]~q  & (!cuifregS_0 & cuifregS_1)))

	.dataa(\registerArray[2][25]~q ),
	.datab(cuifregS_0),
	.datac(cuifregS_1),
	.datad(\Mux6~14_combout ),
	.cin(gnd),
	.combout(\Mux6~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~15 .lut_mask = 16'hFF20;
defparam \Mux6~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N6
cycloneive_lcell_comb \Mux6~12 (
// Equation(s):
// \Mux6~12_combout  = (cuifregS_0 & (((cuifregS_1) # (\registerArray[5][25]~q )))) # (!cuifregS_0 & (\registerArray[4][25]~q  & (!cuifregS_1)))

	.dataa(cuifregS_0),
	.datab(\registerArray[4][25]~q ),
	.datac(cuifregS_1),
	.datad(\registerArray[5][25]~q ),
	.cin(gnd),
	.combout(\Mux6~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~12 .lut_mask = 16'hAEA4;
defparam \Mux6~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N0
cycloneive_lcell_comb \Mux6~13 (
// Equation(s):
// \Mux6~13_combout  = (cuifregS_1 & ((\Mux6~12_combout  & (\registerArray[7][25]~q )) # (!\Mux6~12_combout  & ((\registerArray[6][25]~q ))))) # (!cuifregS_1 & (((\Mux6~12_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[7][25]~q ),
	.datac(\registerArray[6][25]~q ),
	.datad(\Mux6~12_combout ),
	.cin(gnd),
	.combout(\Mux6~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~13 .lut_mask = 16'hDDA0;
defparam \Mux6~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N10
cycloneive_lcell_comb \Mux6~16 (
// Equation(s):
// \Mux6~16_combout  = (cuifregS_2 & ((cuifregS_3) # ((\Mux6~13_combout )))) # (!cuifregS_2 & (!cuifregS_3 & (\Mux6~15_combout )))

	.dataa(cuifregS_2),
	.datab(cuifregS_3),
	.datac(\Mux6~15_combout ),
	.datad(\Mux6~13_combout ),
	.cin(gnd),
	.combout(\Mux6~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~16 .lut_mask = 16'hBA98;
defparam \Mux6~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y41_N28
cycloneive_lcell_comb \Mux6~19 (
// Equation(s):
// \Mux6~19_combout  = (cuifregS_3 & ((\Mux6~16_combout  & ((\Mux6~18_combout ))) # (!\Mux6~16_combout  & (\Mux6~11_combout )))) # (!cuifregS_3 & (((\Mux6~16_combout ))))

	.dataa(\Mux6~11_combout ),
	.datab(cuifregS_3),
	.datac(\Mux6~18_combout ),
	.datad(\Mux6~16_combout ),
	.cin(gnd),
	.combout(\Mux6~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~19 .lut_mask = 16'hF388;
defparam \Mux6~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N2
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & ((\registerArray[25][24]~q ))) # (!cuifregS_3 & (\registerArray[17][24]~q ))))

	.dataa(\registerArray[17][24]~q ),
	.datab(\registerArray[25][24]~q ),
	.datac(cuifregS_2),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hFC0A;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N10
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// \Mux7~1_combout  = (cuifregS_2 & ((\Mux7~0_combout  & ((\registerArray[29][24]~q ))) # (!\Mux7~0_combout  & (\registerArray[21][24]~q )))) # (!cuifregS_2 & (((\Mux7~0_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[21][24]~q ),
	.datac(\Mux7~0_combout ),
	.datad(\registerArray[29][24]~q ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hF858;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y37_N10
cycloneive_lcell_comb \registerArray[16][24]~feeder (
// Equation(s):
// \registerArray[16][24]~feeder_combout  = \Mux44~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux442),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[16][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[16][24]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[16][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y37_N11
dffeas \registerArray[16][24] (
	.clk(clk),
	.d(\registerArray[16][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][24] .is_wysiwyg = "true";
defparam \registerArray[16][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N2
cycloneive_lcell_comb \Mux7~4 (
// Equation(s):
// \Mux7~4_combout  = (cuifregS_2 & ((\registerArray[20][24]~q ) # ((cuifregS_3)))) # (!cuifregS_2 & (((\registerArray[16][24]~q  & !cuifregS_3))))

	.dataa(\registerArray[20][24]~q ),
	.datab(\registerArray[16][24]~q ),
	.datac(cuifregS_2),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux7~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~4 .lut_mask = 16'hF0AC;
defparam \Mux7~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N4
cycloneive_lcell_comb \Mux7~5 (
// Equation(s):
// \Mux7~5_combout  = (cuifregS_3 & ((\Mux7~4_combout  & (\registerArray[28][24]~q )) # (!\Mux7~4_combout  & ((\registerArray[24][24]~q ))))) # (!cuifregS_3 & (((\Mux7~4_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[28][24]~q ),
	.datac(\registerArray[24][24]~q ),
	.datad(\Mux7~4_combout ),
	.cin(gnd),
	.combout(\Mux7~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~5 .lut_mask = 16'hDDA0;
defparam \Mux7~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N8
cycloneive_lcell_comb \Mux7~2 (
// Equation(s):
// \Mux7~2_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[22][24]~q ))) # (!cuifregS_2 & (\registerArray[18][24]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[18][24]~q ),
	.datac(\registerArray[22][24]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~2 .lut_mask = 16'hFA44;
defparam \Mux7~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N11
dffeas \registerArray[26][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][24] .is_wysiwyg = "true";
defparam \registerArray[26][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N10
cycloneive_lcell_comb \Mux7~3 (
// Equation(s):
// \Mux7~3_combout  = (cuifregS_3 & ((\Mux7~2_combout  & ((\registerArray[30][24]~q ))) # (!\Mux7~2_combout  & (\registerArray[26][24]~q )))) # (!cuifregS_3 & (\Mux7~2_combout ))

	.dataa(cuifregS_3),
	.datab(\Mux7~2_combout ),
	.datac(\registerArray[26][24]~q ),
	.datad(\registerArray[30][24]~q ),
	.cin(gnd),
	.combout(\Mux7~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~3 .lut_mask = 16'hEC64;
defparam \Mux7~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N26
cycloneive_lcell_comb \Mux7~6 (
// Equation(s):
// \Mux7~6_combout  = (cuifregS_0 & (cuifregS_1)) # (!cuifregS_0 & ((cuifregS_1 & ((\Mux7~3_combout ))) # (!cuifregS_1 & (\Mux7~5_combout ))))

	.dataa(cuifregS_0),
	.datab(cuifregS_1),
	.datac(\Mux7~5_combout ),
	.datad(\Mux7~3_combout ),
	.cin(gnd),
	.combout(\Mux7~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~6 .lut_mask = 16'hDC98;
defparam \Mux7~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y41_N21
dffeas \registerArray[23][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][24] .is_wysiwyg = "true";
defparam \registerArray[23][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N12
cycloneive_lcell_comb \Mux7~7 (
// Equation(s):
// \Mux7~7_combout  = (cuifregS_3 & (((\registerArray[27][24]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[19][24]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[19][24]~q ),
	.datac(\registerArray[27][24]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux7~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~7 .lut_mask = 16'hAAE4;
defparam \Mux7~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N20
cycloneive_lcell_comb \Mux7~8 (
// Equation(s):
// \Mux7~8_combout  = (cuifregS_2 & ((\Mux7~7_combout  & (\registerArray[31][24]~q )) # (!\Mux7~7_combout  & ((\registerArray[23][24]~q ))))) # (!cuifregS_2 & (((\Mux7~7_combout ))))

	.dataa(\registerArray[31][24]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[23][24]~q ),
	.datad(\Mux7~7_combout ),
	.cin(gnd),
	.combout(\Mux7~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~8 .lut_mask = 16'hBBC0;
defparam \Mux7~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N22
cycloneive_lcell_comb \Mux7~9 (
// Equation(s):
// \Mux7~9_combout  = (cuifregS_0 & ((\Mux7~6_combout  & ((\Mux7~8_combout ))) # (!\Mux7~6_combout  & (\Mux7~1_combout )))) # (!cuifregS_0 & (((\Mux7~6_combout ))))

	.dataa(\Mux7~1_combout ),
	.datab(cuifregS_0),
	.datac(\Mux7~6_combout ),
	.datad(\Mux7~8_combout ),
	.cin(gnd),
	.combout(\Mux7~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~9 .lut_mask = 16'hF838;
defparam \Mux7~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N24
cycloneive_lcell_comb \Mux7~17 (
// Equation(s):
// \Mux7~17_combout  = (cuifregS_0 & (((\registerArray[13][24]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[12][24]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[12][24]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[13][24]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux7~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~17 .lut_mask = 16'hCCE2;
defparam \Mux7~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N24
cycloneive_lcell_comb \Mux7~18 (
// Equation(s):
// \Mux7~18_combout  = (cuifregS_1 & ((\Mux7~17_combout  & ((\registerArray[15][24]~q ))) # (!\Mux7~17_combout  & (\registerArray[14][24]~q )))) # (!cuifregS_1 & (((\Mux7~17_combout ))))

	.dataa(\registerArray[14][24]~q ),
	.datab(\registerArray[15][24]~q ),
	.datac(cuifregS_1),
	.datad(\Mux7~17_combout ),
	.cin(gnd),
	.combout(\Mux7~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~18 .lut_mask = 16'hCFA0;
defparam \Mux7~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N31
dffeas \registerArray[3][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][24] .is_wysiwyg = "true";
defparam \registerArray[3][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N30
cycloneive_lcell_comb \Mux7~14 (
// Equation(s):
// \Mux7~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][24]~q ))) # (!cuifregS_1 & (\registerArray[1][24]~q ))))

	.dataa(\registerArray[1][24]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[3][24]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux7~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~14 .lut_mask = 16'hC088;
defparam \Mux7~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N20
cycloneive_lcell_comb \Mux7~15 (
// Equation(s):
// \Mux7~15_combout  = (\Mux7~14_combout ) # ((cuifregS_1 & (!cuifregS_0 & \registerArray[2][24]~q )))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\registerArray[2][24]~q ),
	.datad(\Mux7~14_combout ),
	.cin(gnd),
	.combout(\Mux7~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~15 .lut_mask = 16'hFF20;
defparam \Mux7~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y43_N7
dffeas \registerArray[10][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][24] .is_wysiwyg = "true";
defparam \registerArray[10][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N6
cycloneive_lcell_comb \Mux7~12 (
// Equation(s):
// \Mux7~12_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][24]~q ))) # (!cuifregS_1 & (\registerArray[8][24]~q ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[8][24]~q ),
	.datac(\registerArray[10][24]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux7~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~12 .lut_mask = 16'hFA44;
defparam \Mux7~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N24
cycloneive_lcell_comb \Mux7~13 (
// Equation(s):
// \Mux7~13_combout  = (cuifregS_0 & ((\Mux7~12_combout  & (\registerArray[11][24]~q )) # (!\Mux7~12_combout  & ((\registerArray[9][24]~q ))))) # (!cuifregS_0 & (((\Mux7~12_combout ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[11][24]~q ),
	.datac(\registerArray[9][24]~q ),
	.datad(\Mux7~12_combout ),
	.cin(gnd),
	.combout(\Mux7~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~13 .lut_mask = 16'hDDA0;
defparam \Mux7~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N26
cycloneive_lcell_comb \Mux7~16 (
// Equation(s):
// \Mux7~16_combout  = (cuifregS_3 & (((cuifregS_2) # (\Mux7~13_combout )))) # (!cuifregS_3 & (\Mux7~15_combout  & (!cuifregS_2)))

	.dataa(cuifregS_3),
	.datab(\Mux7~15_combout ),
	.datac(cuifregS_2),
	.datad(\Mux7~13_combout ),
	.cin(gnd),
	.combout(\Mux7~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~16 .lut_mask = 16'hAEA4;
defparam \Mux7~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y42_N7
dffeas \registerArray[7][24] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux442),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~77_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[7][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[7][24] .is_wysiwyg = "true";
defparam \registerArray[7][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y42_N20
cycloneive_lcell_comb \Mux7~11 (
// Equation(s):
// \Mux7~11_combout  = (\Mux7~10_combout  & (((\registerArray[7][24]~q )) # (!cuifregS_1))) # (!\Mux7~10_combout  & (cuifregS_1 & (\registerArray[6][24]~q )))

	.dataa(\Mux7~10_combout ),
	.datab(cuifregS_1),
	.datac(\registerArray[6][24]~q ),
	.datad(\registerArray[7][24]~q ),
	.cin(gnd),
	.combout(\Mux7~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~11 .lut_mask = 16'hEA62;
defparam \Mux7~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y37_N0
cycloneive_lcell_comb \Mux7~19 (
// Equation(s):
// \Mux7~19_combout  = (cuifregS_2 & ((\Mux7~16_combout  & (\Mux7~18_combout )) # (!\Mux7~16_combout  & ((\Mux7~11_combout ))))) # (!cuifregS_2 & (((\Mux7~16_combout ))))

	.dataa(cuifregS_2),
	.datab(\Mux7~18_combout ),
	.datac(\Mux7~16_combout ),
	.datad(\Mux7~11_combout ),
	.cin(gnd),
	.combout(\Mux7~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~19 .lut_mask = 16'hDAD0;
defparam \Mux7~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N28
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// \Mux8~0_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[21][23]~q ))) # (!cuifregS_2 & (\registerArray[17][23]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[17][23]~q ),
	.datac(\registerArray[21][23]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hFA44;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N14
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// \Mux8~1_combout  = (\Mux8~0_combout  & ((\registerArray[29][23]~q ) # ((!cuifregS_3)))) # (!\Mux8~0_combout  & (((\registerArray[25][23]~q  & cuifregS_3))))

	.dataa(\registerArray[29][23]~q ),
	.datab(\Mux8~0_combout ),
	.datac(\registerArray[25][23]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'hB8CC;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N12
cycloneive_lcell_comb \registerArray[24][23]~feeder (
// Equation(s):
// \registerArray[24][23]~feeder_combout  = \Mux45~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux452),
	.cin(gnd),
	.combout(\registerArray[24][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[24][23]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[24][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y41_N13
dffeas \registerArray[24][23] (
	.clk(clk),
	.d(\registerArray[24][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][23] .is_wysiwyg = "true";
defparam \registerArray[24][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N16
cycloneive_lcell_comb \Mux8~4 (
// Equation(s):
// \Mux8~4_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & ((\registerArray[24][23]~q ))) # (!cuifregS_3 & (\registerArray[16][23]~q ))))

	.dataa(\registerArray[16][23]~q ),
	.datab(\registerArray[24][23]~q ),
	.datac(cuifregS_2),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux8~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~4 .lut_mask = 16'hFC0A;
defparam \Mux8~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y41_N10
cycloneive_lcell_comb \Mux8~5 (
// Equation(s):
// \Mux8~5_combout  = (cuifregS_2 & ((\Mux8~4_combout  & ((\registerArray[28][23]~q ))) # (!\Mux8~4_combout  & (\registerArray[20][23]~q )))) # (!cuifregS_2 & (((\Mux8~4_combout ))))

	.dataa(\registerArray[20][23]~q ),
	.datab(\registerArray[28][23]~q ),
	.datac(cuifregS_2),
	.datad(\Mux8~4_combout ),
	.cin(gnd),
	.combout(\Mux8~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~5 .lut_mask = 16'hCFA0;
defparam \Mux8~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N8
cycloneive_lcell_comb \Mux8~6 (
// Equation(s):
// \Mux8~6_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\Mux8~3_combout )) # (!cuifregS_1 & ((\Mux8~5_combout )))))

	.dataa(\Mux8~3_combout ),
	.datab(cuifregS_0),
	.datac(\Mux8~5_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux8~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~6 .lut_mask = 16'hEE30;
defparam \Mux8~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N23
dffeas \registerArray[27][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][23] .is_wysiwyg = "true";
defparam \registerArray[27][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N0
cycloneive_lcell_comb \Mux8~7 (
// Equation(s):
// \Mux8~7_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & (\registerArray[23][23]~q )) # (!cuifregS_2 & ((\registerArray[19][23]~q )))))

	.dataa(cuifregS_3),
	.datab(\registerArray[23][23]~q ),
	.datac(\registerArray[19][23]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux8~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~7 .lut_mask = 16'hEE50;
defparam \Mux8~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N22
cycloneive_lcell_comb \Mux8~8 (
// Equation(s):
// \Mux8~8_combout  = (cuifregS_3 & ((\Mux8~7_combout  & (\registerArray[31][23]~q )) # (!\Mux8~7_combout  & ((\registerArray[27][23]~q ))))) # (!cuifregS_3 & (((\Mux8~7_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[31][23]~q ),
	.datac(\registerArray[27][23]~q ),
	.datad(\Mux8~7_combout ),
	.cin(gnd),
	.combout(\Mux8~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~8 .lut_mask = 16'hDDA0;
defparam \Mux8~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N30
cycloneive_lcell_comb \Mux8~9 (
// Equation(s):
// \Mux8~9_combout  = (cuifregS_0 & ((\Mux8~6_combout  & ((\Mux8~8_combout ))) # (!\Mux8~6_combout  & (\Mux8~1_combout )))) # (!cuifregS_0 & (((\Mux8~6_combout ))))

	.dataa(cuifregS_0),
	.datab(\Mux8~1_combout ),
	.datac(\Mux8~6_combout ),
	.datad(\Mux8~8_combout ),
	.cin(gnd),
	.combout(\Mux8~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~9 .lut_mask = 16'hF858;
defparam \Mux8~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N17
dffeas \registerArray[3][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][23] .is_wysiwyg = "true";
defparam \registerArray[3][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N16
cycloneive_lcell_comb \Mux8~14 (
// Equation(s):
// \Mux8~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][23]~q ))) # (!cuifregS_1 & (\registerArray[1][23]~q ))))

	.dataa(\registerArray[1][23]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[3][23]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux8~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~14 .lut_mask = 16'hC088;
defparam \Mux8~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N28
cycloneive_lcell_comb \Mux8~15 (
// Equation(s):
// \Mux8~15_combout  = (\Mux8~14_combout ) # ((cuifregS_1 & (!cuifregS_0 & \registerArray[2][23]~q )))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\registerArray[2][23]~q ),
	.datad(\Mux8~14_combout ),
	.cin(gnd),
	.combout(\Mux8~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~15 .lut_mask = 16'hFF20;
defparam \Mux8~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N1
dffeas \registerArray[5][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][23] .is_wysiwyg = "true";
defparam \registerArray[5][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N0
cycloneive_lcell_comb \Mux8~12 (
// Equation(s):
// \Mux8~12_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & ((\registerArray[5][23]~q ))) # (!cuifregS_0 & (\registerArray[4][23]~q ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[4][23]~q ),
	.datac(\registerArray[5][23]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux8~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~12 .lut_mask = 16'hFA44;
defparam \Mux8~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N10
cycloneive_lcell_comb \Mux8~13 (
// Equation(s):
// \Mux8~13_combout  = (cuifregS_1 & ((\Mux8~12_combout  & ((\registerArray[7][23]~q ))) # (!\Mux8~12_combout  & (\registerArray[6][23]~q )))) # (!cuifregS_1 & (\Mux8~12_combout ))

	.dataa(cuifregS_1),
	.datab(\Mux8~12_combout ),
	.datac(\registerArray[6][23]~q ),
	.datad(\registerArray[7][23]~q ),
	.cin(gnd),
	.combout(\Mux8~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~13 .lut_mask = 16'hEC64;
defparam \Mux8~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N14
cycloneive_lcell_comb \Mux8~16 (
// Equation(s):
// \Mux8~16_combout  = (cuifregS_2 & (((\Mux8~13_combout ) # (cuifregS_3)))) # (!cuifregS_2 & (\Mux8~15_combout  & ((!cuifregS_3))))

	.dataa(cuifregS_2),
	.datab(\Mux8~15_combout ),
	.datac(\Mux8~13_combout ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux8~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~16 .lut_mask = 16'hAAE4;
defparam \Mux8~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N0
cycloneive_lcell_comb \Mux8~17 (
// Equation(s):
// \Mux8~17_combout  = (cuifregS_0 & (((\registerArray[13][23]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[12][23]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[12][23]~q ),
	.datab(\registerArray[13][23]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux8~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~17 .lut_mask = 16'hF0CA;
defparam \Mux8~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N14
cycloneive_lcell_comb \Mux8~18 (
// Equation(s):
// \Mux8~18_combout  = (cuifregS_1 & ((\Mux8~17_combout  & ((\registerArray[15][23]~q ))) # (!\Mux8~17_combout  & (\registerArray[14][23]~q )))) # (!cuifregS_1 & (((\Mux8~17_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[14][23]~q ),
	.datac(\registerArray[15][23]~q ),
	.datad(\Mux8~17_combout ),
	.cin(gnd),
	.combout(\Mux8~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~18 .lut_mask = 16'hF588;
defparam \Mux8~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y43_N15
dffeas \registerArray[10][23] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux452),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][23] .is_wysiwyg = "true";
defparam \registerArray[10][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N14
cycloneive_lcell_comb \Mux8~10 (
// Equation(s):
// \Mux8~10_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][23]~q ))) # (!cuifregS_1 & (\registerArray[8][23]~q ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[8][23]~q ),
	.datac(\registerArray[10][23]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux8~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~10 .lut_mask = 16'hFA44;
defparam \Mux8~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N28
cycloneive_lcell_comb \Mux8~11 (
// Equation(s):
// \Mux8~11_combout  = (\Mux8~10_combout  & ((\registerArray[11][23]~q ) # ((!cuifregS_0)))) # (!\Mux8~10_combout  & (((\registerArray[9][23]~q  & cuifregS_0))))

	.dataa(\registerArray[11][23]~q ),
	.datab(\Mux8~10_combout ),
	.datac(\registerArray[9][23]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux8~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~11 .lut_mask = 16'hB8CC;
defparam \Mux8~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N20
cycloneive_lcell_comb \Mux8~19 (
// Equation(s):
// \Mux8~19_combout  = (cuifregS_3 & ((\Mux8~16_combout  & (\Mux8~18_combout )) # (!\Mux8~16_combout  & ((\Mux8~11_combout ))))) # (!cuifregS_3 & (\Mux8~16_combout ))

	.dataa(cuifregS_3),
	.datab(\Mux8~16_combout ),
	.datac(\Mux8~18_combout ),
	.datad(\Mux8~11_combout ),
	.cin(gnd),
	.combout(\Mux8~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~19 .lut_mask = 16'hE6C4;
defparam \Mux8~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N27
dffeas \registerArray[3][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][22] .is_wysiwyg = "true";
defparam \registerArray[3][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N26
cycloneive_lcell_comb \Mux9~14 (
// Equation(s):
// \Mux9~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][22]~q ))) # (!cuifregS_1 & (\registerArray[1][22]~q ))))

	.dataa(\registerArray[1][22]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[3][22]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux9~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~14 .lut_mask = 16'hC088;
defparam \Mux9~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N0
cycloneive_lcell_comb \Mux9~15 (
// Equation(s):
// \Mux9~15_combout  = (\Mux9~14_combout ) # ((\registerArray[2][22]~q  & (!cuifregS_0 & cuifregS_1)))

	.dataa(\registerArray[2][22]~q ),
	.datab(cuifregS_0),
	.datac(cuifregS_1),
	.datad(\Mux9~14_combout ),
	.cin(gnd),
	.combout(\Mux9~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~15 .lut_mask = 16'hFF20;
defparam \Mux9~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N26
cycloneive_lcell_comb \registerArray[10][22]~feeder (
// Equation(s):
// \registerArray[10][22]~feeder_combout  = \Mux46~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux462),
	.cin(gnd),
	.combout(\registerArray[10][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[10][22]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[10][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y43_N27
dffeas \registerArray[10][22] (
	.clk(clk),
	.d(\registerArray[10][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][22] .is_wysiwyg = "true";
defparam \registerArray[10][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N16
cycloneive_lcell_comb \Mux9~12 (
// Equation(s):
// \Mux9~12_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][22]~q ))) # (!cuifregS_1 & (\registerArray[8][22]~q ))))

	.dataa(\registerArray[8][22]~q ),
	.datab(\registerArray[10][22]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux9~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~12 .lut_mask = 16'hFC0A;
defparam \Mux9~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y43_N10
cycloneive_lcell_comb \Mux9~13 (
// Equation(s):
// \Mux9~13_combout  = (cuifregS_0 & ((\Mux9~12_combout  & ((\registerArray[11][22]~q ))) # (!\Mux9~12_combout  & (\registerArray[9][22]~q )))) # (!cuifregS_0 & (((\Mux9~12_combout ))))

	.dataa(\registerArray[9][22]~q ),
	.datab(\registerArray[11][22]~q ),
	.datac(cuifregS_0),
	.datad(\Mux9~12_combout ),
	.cin(gnd),
	.combout(\Mux9~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~13 .lut_mask = 16'hCFA0;
defparam \Mux9~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N2
cycloneive_lcell_comb \Mux9~16 (
// Equation(s):
// \Mux9~16_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & ((\Mux9~13_combout ))) # (!cuifregS_3 & (\Mux9~15_combout ))))

	.dataa(cuifregS_2),
	.datab(\Mux9~15_combout ),
	.datac(\Mux9~13_combout ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux9~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~16 .lut_mask = 16'hFA44;
defparam \Mux9~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y39_N12
cycloneive_lcell_comb \Mux9~17 (
// Equation(s):
// \Mux9~17_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & (\registerArray[13][22]~q )) # (!cuifregS_0 & ((\registerArray[12][22]~q )))))

	.dataa(\registerArray[13][22]~q ),
	.datab(\registerArray[12][22]~q ),
	.datac(cuifregS_1),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux9~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~17 .lut_mask = 16'hFA0C;
defparam \Mux9~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N14
cycloneive_lcell_comb \Mux9~18 (
// Equation(s):
// \Mux9~18_combout  = (cuifregS_1 & ((\Mux9~17_combout  & (\registerArray[15][22]~q )) # (!\Mux9~17_combout  & ((\registerArray[14][22]~q ))))) # (!cuifregS_1 & (((\Mux9~17_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[15][22]~q ),
	.datac(\registerArray[14][22]~q ),
	.datad(\Mux9~17_combout ),
	.cin(gnd),
	.combout(\Mux9~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~18 .lut_mask = 16'hDDA0;
defparam \Mux9~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N23
dffeas \registerArray[6][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][22] .is_wysiwyg = "true";
defparam \registerArray[6][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N8
cycloneive_lcell_comb \Mux9~10 (
// Equation(s):
// \Mux9~10_combout  = (cuifregS_0 & (((\registerArray[5][22]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[4][22]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[4][22]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[5][22]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux9~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~10 .lut_mask = 16'hCCE2;
defparam \Mux9~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N22
cycloneive_lcell_comb \Mux9~11 (
// Equation(s):
// \Mux9~11_combout  = (cuifregS_1 & ((\Mux9~10_combout  & (\registerArray[7][22]~q )) # (!\Mux9~10_combout  & ((\registerArray[6][22]~q ))))) # (!cuifregS_1 & (((\Mux9~10_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[7][22]~q ),
	.datac(\registerArray[6][22]~q ),
	.datad(\Mux9~10_combout ),
	.cin(gnd),
	.combout(\Mux9~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~11 .lut_mask = 16'hDDA0;
defparam \Mux9~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N4
cycloneive_lcell_comb \Mux9~19 (
// Equation(s):
// \Mux9~19_combout  = (cuifregS_2 & ((\Mux9~16_combout  & (\Mux9~18_combout )) # (!\Mux9~16_combout  & ((\Mux9~11_combout ))))) # (!cuifregS_2 & (\Mux9~16_combout ))

	.dataa(cuifregS_2),
	.datab(\Mux9~16_combout ),
	.datac(\Mux9~18_combout ),
	.datad(\Mux9~11_combout ),
	.cin(gnd),
	.combout(\Mux9~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~19 .lut_mask = 16'hE6C4;
defparam \Mux9~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y41_N13
dffeas \registerArray[23][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][22] .is_wysiwyg = "true";
defparam \registerArray[23][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N4
cycloneive_lcell_comb \Mux9~7 (
// Equation(s):
// \Mux9~7_combout  = (cuifregS_3 & (((\registerArray[27][22]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[19][22]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[19][22]~q ),
	.datac(\registerArray[27][22]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux9~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~7 .lut_mask = 16'hAAE4;
defparam \Mux9~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N12
cycloneive_lcell_comb \Mux9~8 (
// Equation(s):
// \Mux9~8_combout  = (cuifregS_2 & ((\Mux9~7_combout  & (\registerArray[31][22]~q )) # (!\Mux9~7_combout  & ((\registerArray[23][22]~q ))))) # (!cuifregS_2 & (((\Mux9~7_combout ))))

	.dataa(\registerArray[31][22]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[23][22]~q ),
	.datad(\Mux9~7_combout ),
	.cin(gnd),
	.combout(\Mux9~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~8 .lut_mask = 16'hBBC0;
defparam \Mux9~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N8
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// \Mux9~0_combout  = (cuifregS_3 & (((\registerArray[25][22]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[17][22]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[17][22]~q ),
	.datac(\registerArray[25][22]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hAAE4;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N22
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// \Mux9~1_combout  = (\Mux9~0_combout  & ((\registerArray[29][22]~q ) # ((!cuifregS_2)))) # (!\Mux9~0_combout  & (((\registerArray[21][22]~q  & cuifregS_2))))

	.dataa(\registerArray[29][22]~q ),
	.datab(\Mux9~0_combout ),
	.datac(\registerArray[21][22]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'hB8CC;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N28
cycloneive_lcell_comb \Mux9~2 (
// Equation(s):
// \Mux9~2_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[22][22]~q ))) # (!cuifregS_2 & (\registerArray[18][22]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[18][22]~q ),
	.datac(\registerArray[22][22]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux9~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~2 .lut_mask = 16'hFA44;
defparam \Mux9~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N30
cycloneive_lcell_comb \Mux9~3 (
// Equation(s):
// \Mux9~3_combout  = (cuifregS_3 & ((\Mux9~2_combout  & (\registerArray[30][22]~q )) # (!\Mux9~2_combout  & ((\registerArray[26][22]~q ))))) # (!cuifregS_3 & (((\Mux9~2_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[30][22]~q ),
	.datac(\registerArray[26][22]~q ),
	.datad(\Mux9~2_combout ),
	.cin(gnd),
	.combout(\Mux9~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~3 .lut_mask = 16'hDDA0;
defparam \Mux9~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N17
dffeas \registerArray[20][22] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux462),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][22] .is_wysiwyg = "true";
defparam \registerArray[20][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N16
cycloneive_lcell_comb \Mux9~4 (
// Equation(s):
// \Mux9~4_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[20][22]~q ))) # (!cuifregS_2 & (\registerArray[16][22]~q ))))

	.dataa(\registerArray[16][22]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[20][22]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux9~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~4 .lut_mask = 16'hFC22;
defparam \Mux9~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N12
cycloneive_lcell_comb \Mux9~5 (
// Equation(s):
// \Mux9~5_combout  = (cuifregS_3 & ((\Mux9~4_combout  & (\registerArray[28][22]~q )) # (!\Mux9~4_combout  & ((\registerArray[24][22]~q ))))) # (!cuifregS_3 & (((\Mux9~4_combout ))))

	.dataa(\registerArray[28][22]~q ),
	.datab(\registerArray[24][22]~q ),
	.datac(cuifregS_3),
	.datad(\Mux9~4_combout ),
	.cin(gnd),
	.combout(\Mux9~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~5 .lut_mask = 16'hAFC0;
defparam \Mux9~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N16
cycloneive_lcell_comb \Mux9~6 (
// Equation(s):
// \Mux9~6_combout  = (cuifregS_1 & ((cuifregS_0) # ((\Mux9~3_combout )))) # (!cuifregS_1 & (!cuifregS_0 & ((\Mux9~5_combout ))))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\Mux9~3_combout ),
	.datad(\Mux9~5_combout ),
	.cin(gnd),
	.combout(\Mux9~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~6 .lut_mask = 16'hB9A8;
defparam \Mux9~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y41_N18
cycloneive_lcell_comb \Mux9~9 (
// Equation(s):
// \Mux9~9_combout  = (cuifregS_0 & ((\Mux9~6_combout  & (\Mux9~8_combout )) # (!\Mux9~6_combout  & ((\Mux9~1_combout ))))) # (!cuifregS_0 & (((\Mux9~6_combout ))))

	.dataa(cuifregS_0),
	.datab(\Mux9~8_combout ),
	.datac(\Mux9~1_combout ),
	.datad(\Mux9~6_combout ),
	.cin(gnd),
	.combout(\Mux9~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~9 .lut_mask = 16'hDDA0;
defparam \Mux9~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N6
cycloneive_lcell_comb \Mux10~17 (
// Equation(s):
// \Mux10~17_combout  = (cuifregS_0 & (((\registerArray[13][21]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[12][21]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[12][21]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[13][21]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux10~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~17 .lut_mask = 16'hCCE2;
defparam \Mux10~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N12
cycloneive_lcell_comb \Mux10~18 (
// Equation(s):
// \Mux10~18_combout  = (cuifregS_1 & ((\Mux10~17_combout  & (\registerArray[15][21]~q )) # (!\Mux10~17_combout  & ((\registerArray[14][21]~q ))))) # (!cuifregS_1 & (((\Mux10~17_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[15][21]~q ),
	.datac(\registerArray[14][21]~q ),
	.datad(\Mux10~17_combout ),
	.cin(gnd),
	.combout(\Mux10~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~18 .lut_mask = 16'hDDA0;
defparam \Mux10~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y42_N1
dffeas \registerArray[3][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][21] .is_wysiwyg = "true";
defparam \registerArray[3][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N0
cycloneive_lcell_comb \Mux10~14 (
// Equation(s):
// \Mux10~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][21]~q ))) # (!cuifregS_1 & (\registerArray[1][21]~q ))))

	.dataa(\registerArray[1][21]~q ),
	.datab(cuifregS_1),
	.datac(\registerArray[3][21]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux10~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~14 .lut_mask = 16'hE200;
defparam \Mux10~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y42_N20
cycloneive_lcell_comb \Mux10~15 (
// Equation(s):
// \Mux10~15_combout  = (\Mux10~14_combout ) # ((\registerArray[2][21]~q  & (cuifregS_1 & !cuifregS_0)))

	.dataa(\registerArray[2][21]~q ),
	.datab(\Mux10~14_combout ),
	.datac(cuifregS_1),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux10~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~15 .lut_mask = 16'hCCEC;
defparam \Mux10~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y38_N13
dffeas \registerArray[5][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][21] .is_wysiwyg = "true";
defparam \registerArray[5][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N12
cycloneive_lcell_comb \Mux10~12 (
// Equation(s):
// \Mux10~12_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & ((\registerArray[5][21]~q ))) # (!cuifregS_0 & (\registerArray[4][21]~q ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[4][21]~q ),
	.datac(\registerArray[5][21]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux10~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~12 .lut_mask = 16'hFA44;
defparam \Mux10~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N10
cycloneive_lcell_comb \Mux10~13 (
// Equation(s):
// \Mux10~13_combout  = (cuifregS_1 & ((\Mux10~12_combout  & (\registerArray[7][21]~q )) # (!\Mux10~12_combout  & ((\registerArray[6][21]~q ))))) # (!cuifregS_1 & (((\Mux10~12_combout ))))

	.dataa(\registerArray[7][21]~q ),
	.datab(\registerArray[6][21]~q ),
	.datac(cuifregS_1),
	.datad(\Mux10~12_combout ),
	.cin(gnd),
	.combout(\Mux10~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~13 .lut_mask = 16'hAFC0;
defparam \Mux10~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N4
cycloneive_lcell_comb \Mux10~16 (
// Equation(s):
// \Mux10~16_combout  = (cuifregS_2 & ((cuifregS_3) # ((\Mux10~13_combout )))) # (!cuifregS_2 & (!cuifregS_3 & (\Mux10~15_combout )))

	.dataa(cuifregS_2),
	.datab(cuifregS_3),
	.datac(\Mux10~15_combout ),
	.datad(\Mux10~13_combout ),
	.cin(gnd),
	.combout(\Mux10~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~16 .lut_mask = 16'hBA98;
defparam \Mux10~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y42_N4
cycloneive_lcell_comb \registerArray[11][21]~feeder (
// Equation(s):
// \registerArray[11][21]~feeder_combout  = \Mux47~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux472),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[11][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[11][21]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[11][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y42_N5
dffeas \registerArray[11][21] (
	.clk(clk),
	.d(\registerArray[11][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~75_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[11][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[11][21] .is_wysiwyg = "true";
defparam \registerArray[11][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N0
cycloneive_lcell_comb \Mux10~11 (
// Equation(s):
// \Mux10~11_combout  = (\Mux10~10_combout  & ((\registerArray[11][21]~q ) # ((!cuifregS_0)))) # (!\Mux10~10_combout  & (((\registerArray[9][21]~q  & cuifregS_0))))

	.dataa(\Mux10~10_combout ),
	.datab(\registerArray[11][21]~q ),
	.datac(\registerArray[9][21]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux10~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~11 .lut_mask = 16'hD8AA;
defparam \Mux10~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N22
cycloneive_lcell_comb \Mux10~19 (
// Equation(s):
// \Mux10~19_combout  = (cuifregS_3 & ((\Mux10~16_combout  & (\Mux10~18_combout )) # (!\Mux10~16_combout  & ((\Mux10~11_combout ))))) # (!cuifregS_3 & (((\Mux10~16_combout ))))

	.dataa(\Mux10~18_combout ),
	.datab(cuifregS_3),
	.datac(\Mux10~16_combout ),
	.datad(\Mux10~11_combout ),
	.cin(gnd),
	.combout(\Mux10~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~19 .lut_mask = 16'hBCB0;
defparam \Mux10~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N12
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// \Mux10~0_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[21][21]~q ))) # (!cuifregS_2 & (\registerArray[17][21]~q ))))

	.dataa(\registerArray[17][21]~q ),
	.datab(\registerArray[21][21]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hFC0A;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y44_N18
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// \Mux10~1_combout  = (cuifregS_3 & ((\Mux10~0_combout  & (\registerArray[29][21]~q )) # (!\Mux10~0_combout  & ((\registerArray[25][21]~q ))))) # (!cuifregS_3 & (((\Mux10~0_combout ))))

	.dataa(\registerArray[29][21]~q ),
	.datab(\registerArray[25][21]~q ),
	.datac(cuifregS_3),
	.datad(\Mux10~0_combout ),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'hAFC0;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N16
cycloneive_lcell_comb \Mux10~7 (
// Equation(s):
// \Mux10~7_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[23][21]~q ))) # (!cuifregS_2 & (\registerArray[19][21]~q ))))

	.dataa(\registerArray[19][21]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[23][21]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux10~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~7 .lut_mask = 16'hFC22;
defparam \Mux10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N26
cycloneive_lcell_comb \Mux10~8 (
// Equation(s):
// \Mux10~8_combout  = (cuifregS_3 & ((\Mux10~7_combout  & ((\registerArray[31][21]~q ))) # (!\Mux10~7_combout  & (\registerArray[27][21]~q )))) # (!cuifregS_3 & (((\Mux10~7_combout ))))

	.dataa(\registerArray[27][21]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[31][21]~q ),
	.datad(\Mux10~7_combout ),
	.cin(gnd),
	.combout(\Mux10~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~8 .lut_mask = 16'hF388;
defparam \Mux10~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N19
dffeas \registerArray[24][21] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux472),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~66_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[24][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[24][21] .is_wysiwyg = "true";
defparam \registerArray[24][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y31_N22
cycloneive_lcell_comb \registerArray[16][21]~feeder (
// Equation(s):
// \registerArray[16][21]~feeder_combout  = \Mux47~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux472),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[16][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[16][21]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[16][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y31_N23
dffeas \registerArray[16][21] (
	.clk(clk),
	.d(\registerArray[16][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~56_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[16][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[16][21] .is_wysiwyg = "true";
defparam \registerArray[16][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N18
cycloneive_lcell_comb \Mux10~4 (
// Equation(s):
// \Mux10~4_combout  = (cuifregS_3 & ((cuifregS_2) # ((\registerArray[24][21]~q )))) # (!cuifregS_3 & (!cuifregS_2 & ((\registerArray[16][21]~q ))))

	.dataa(cuifregS_3),
	.datab(cuifregS_2),
	.datac(\registerArray[24][21]~q ),
	.datad(\registerArray[16][21]~q ),
	.cin(gnd),
	.combout(\Mux10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~4 .lut_mask = 16'hB9A8;
defparam \Mux10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N10
cycloneive_lcell_comb \Mux10~5 (
// Equation(s):
// \Mux10~5_combout  = (cuifregS_2 & ((\Mux10~4_combout  & (\registerArray[28][21]~q )) # (!\Mux10~4_combout  & ((\registerArray[20][21]~q ))))) # (!cuifregS_2 & (((\Mux10~4_combout ))))

	.dataa(\registerArray[28][21]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[20][21]~q ),
	.datad(\Mux10~4_combout ),
	.cin(gnd),
	.combout(\Mux10~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~5 .lut_mask = 16'hBBC0;
defparam \Mux10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N24
cycloneive_lcell_comb \Mux10~6 (
// Equation(s):
// \Mux10~6_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\Mux10~3_combout )) # (!cuifregS_1 & ((\Mux10~5_combout )))))

	.dataa(\Mux10~3_combout ),
	.datab(cuifregS_0),
	.datac(\Mux10~5_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux10~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~6 .lut_mask = 16'hEE30;
defparam \Mux10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N16
cycloneive_lcell_comb \Mux10~9 (
// Equation(s):
// \Mux10~9_combout  = (cuifregS_0 & ((\Mux10~6_combout  & ((\Mux10~8_combout ))) # (!\Mux10~6_combout  & (\Mux10~1_combout )))) # (!cuifregS_0 & (((\Mux10~6_combout ))))

	.dataa(\Mux10~1_combout ),
	.datab(cuifregS_0),
	.datac(\Mux10~8_combout ),
	.datad(\Mux10~6_combout ),
	.cin(gnd),
	.combout(\Mux10~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~9 .lut_mask = 16'hF388;
defparam \Mux10~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y39_N30
cycloneive_lcell_comb \Mux11~17 (
// Equation(s):
// \Mux11~17_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & ((\registerArray[13][20]~q ))) # (!cuifregS_0 & (\registerArray[12][20]~q ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[12][20]~q ),
	.datac(\registerArray[13][20]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux11~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~17 .lut_mask = 16'hFA44;
defparam \Mux11~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N30
cycloneive_lcell_comb \Mux11~18 (
// Equation(s):
// \Mux11~18_combout  = (cuifregS_1 & ((\Mux11~17_combout  & (\registerArray[15][20]~q )) # (!\Mux11~17_combout  & ((\registerArray[14][20]~q ))))) # (!cuifregS_1 & (((\Mux11~17_combout ))))

	.dataa(\registerArray[15][20]~q ),
	.datab(cuifregS_1),
	.datac(\registerArray[14][20]~q ),
	.datad(\Mux11~17_combout ),
	.cin(gnd),
	.combout(\Mux11~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~18 .lut_mask = 16'hBBC0;
defparam \Mux11~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y44_N12
cycloneive_lcell_comb \Mux11~12 (
// Equation(s):
// \Mux11~12_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\registerArray[10][20]~q )) # (!cuifregS_1 & ((\registerArray[8][20]~q )))))

	.dataa(\registerArray[10][20]~q ),
	.datab(\registerArray[8][20]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux11~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~12 .lut_mask = 16'hFA0C;
defparam \Mux11~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N18
cycloneive_lcell_comb \Mux11~13 (
// Equation(s):
// \Mux11~13_combout  = (cuifregS_0 & ((\Mux11~12_combout  & ((\registerArray[11][20]~q ))) # (!\Mux11~12_combout  & (\registerArray[9][20]~q )))) # (!cuifregS_0 & (((\Mux11~12_combout ))))

	.dataa(\registerArray[9][20]~q ),
	.datab(\registerArray[11][20]~q ),
	.datac(cuifregS_0),
	.datad(\Mux11~12_combout ),
	.cin(gnd),
	.combout(\Mux11~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~13 .lut_mask = 16'hCFA0;
defparam \Mux11~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N8
cycloneive_lcell_comb \Mux11~16 (
// Equation(s):
// \Mux11~16_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & ((\Mux11~13_combout ))) # (!cuifregS_3 & (\Mux11~15_combout ))))

	.dataa(\Mux11~15_combout ),
	.datab(cuifregS_2),
	.datac(cuifregS_3),
	.datad(\Mux11~13_combout ),
	.cin(gnd),
	.combout(\Mux11~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~16 .lut_mask = 16'hF2C2;
defparam \Mux11~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y38_N13
dffeas \registerArray[6][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][20] .is_wysiwyg = "true";
defparam \registerArray[6][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y38_N25
dffeas \registerArray[5][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][20] .is_wysiwyg = "true";
defparam \registerArray[5][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y38_N24
cycloneive_lcell_comb \Mux11~10 (
// Equation(s):
// \Mux11~10_combout  = (cuifregS_0 & (((\registerArray[5][20]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[4][20]~q  & ((!cuifregS_1))))

	.dataa(cuifregS_0),
	.datab(\registerArray[4][20]~q ),
	.datac(\registerArray[5][20]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux11~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~10 .lut_mask = 16'hAAE4;
defparam \Mux11~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N12
cycloneive_lcell_comb \Mux11~11 (
// Equation(s):
// \Mux11~11_combout  = (cuifregS_1 & ((\Mux11~10_combout  & (\registerArray[7][20]~q )) # (!\Mux11~10_combout  & ((\registerArray[6][20]~q ))))) # (!cuifregS_1 & (((\Mux11~10_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[7][20]~q ),
	.datac(\registerArray[6][20]~q ),
	.datad(\Mux11~10_combout ),
	.cin(gnd),
	.combout(\Mux11~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~11 .lut_mask = 16'hDDA0;
defparam \Mux11~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N2
cycloneive_lcell_comb \Mux11~19 (
// Equation(s):
// \Mux11~19_combout  = (cuifregS_2 & ((\Mux11~16_combout  & (\Mux11~18_combout )) # (!\Mux11~16_combout  & ((\Mux11~11_combout ))))) # (!cuifregS_2 & (((\Mux11~16_combout ))))

	.dataa(\Mux11~18_combout ),
	.datab(cuifregS_2),
	.datac(\Mux11~16_combout ),
	.datad(\Mux11~11_combout ),
	.cin(gnd),
	.combout(\Mux11~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~19 .lut_mask = 16'hBCB0;
defparam \Mux11~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y41_N11
dffeas \registerArray[21][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][20] .is_wysiwyg = "true";
defparam \registerArray[21][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N16
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// \Mux11~0_combout  = (cuifregS_3 & (((\registerArray[25][20]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[17][20]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[17][20]~q ),
	.datac(\registerArray[25][20]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hAAE4;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N10
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// \Mux11~1_combout  = (cuifregS_2 & ((\Mux11~0_combout  & (\registerArray[29][20]~q )) # (!\Mux11~0_combout  & ((\registerArray[21][20]~q ))))) # (!cuifregS_2 & (((\Mux11~0_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[29][20]~q ),
	.datac(\registerArray[21][20]~q ),
	.datad(\Mux11~0_combout ),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'hDDA0;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N21
dffeas \registerArray[20][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][20] .is_wysiwyg = "true";
defparam \registerArray[20][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N20
cycloneive_lcell_comb \Mux11~4 (
// Equation(s):
// \Mux11~4_combout  = (cuifregS_2 & ((cuifregS_3) # ((\registerArray[20][20]~q )))) # (!cuifregS_2 & (!cuifregS_3 & ((\registerArray[16][20]~q ))))

	.dataa(cuifregS_2),
	.datab(cuifregS_3),
	.datac(\registerArray[20][20]~q ),
	.datad(\registerArray[16][20]~q ),
	.cin(gnd),
	.combout(\Mux11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~4 .lut_mask = 16'hB9A8;
defparam \Mux11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y38_N14
cycloneive_lcell_comb \Mux11~5 (
// Equation(s):
// \Mux11~5_combout  = (\Mux11~4_combout  & ((\registerArray[28][20]~q ) # ((!cuifregS_3)))) # (!\Mux11~4_combout  & (((\registerArray[24][20]~q  & cuifregS_3))))

	.dataa(\registerArray[28][20]~q ),
	.datab(\Mux11~4_combout ),
	.datac(\registerArray[24][20]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux11~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~5 .lut_mask = 16'hB8CC;
defparam \Mux11~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N24
cycloneive_lcell_comb \Mux11~2 (
// Equation(s):
// \Mux11~2_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[22][20]~q ))) # (!cuifregS_2 & (\registerArray[18][20]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[18][20]~q ),
	.datac(\registerArray[22][20]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~2 .lut_mask = 16'hFA44;
defparam \Mux11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y44_N22
cycloneive_lcell_comb \Mux11~3 (
// Equation(s):
// \Mux11~3_combout  = (\Mux11~2_combout  & ((\registerArray[30][20]~q ) # ((!cuifregS_3)))) # (!\Mux11~2_combout  & (((\registerArray[26][20]~q  & cuifregS_3))))

	.dataa(\registerArray[30][20]~q ),
	.datab(\registerArray[26][20]~q ),
	.datac(\Mux11~2_combout ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~3 .lut_mask = 16'hACF0;
defparam \Mux11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N14
cycloneive_lcell_comb \Mux11~6 (
// Equation(s):
// \Mux11~6_combout  = (cuifregS_1 & ((cuifregS_0) # ((\Mux11~3_combout )))) # (!cuifregS_1 & (!cuifregS_0 & (\Mux11~5_combout )))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\Mux11~5_combout ),
	.datad(\Mux11~3_combout ),
	.cin(gnd),
	.combout(\Mux11~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~6 .lut_mask = 16'hBA98;
defparam \Mux11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y41_N31
dffeas \registerArray[23][20] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux482),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][20] .is_wysiwyg = "true";
defparam \registerArray[23][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N20
cycloneive_lcell_comb \Mux11~7 (
// Equation(s):
// \Mux11~7_combout  = (cuifregS_3 & (((\registerArray[27][20]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[19][20]~q  & ((!cuifregS_2))))

	.dataa(cuifregS_3),
	.datab(\registerArray[19][20]~q ),
	.datac(\registerArray[27][20]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux11~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~7 .lut_mask = 16'hAAE4;
defparam \Mux11~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N30
cycloneive_lcell_comb \Mux11~8 (
// Equation(s):
// \Mux11~8_combout  = (cuifregS_2 & ((\Mux11~7_combout  & (\registerArray[31][20]~q )) # (!\Mux11~7_combout  & ((\registerArray[23][20]~q ))))) # (!cuifregS_2 & (((\Mux11~7_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[31][20]~q ),
	.datac(\registerArray[23][20]~q ),
	.datad(\Mux11~7_combout ),
	.cin(gnd),
	.combout(\Mux11~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~8 .lut_mask = 16'hDDA0;
defparam \Mux11~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y44_N20
cycloneive_lcell_comb \Mux11~9 (
// Equation(s):
// \Mux11~9_combout  = (cuifregS_0 & ((\Mux11~6_combout  & ((\Mux11~8_combout ))) # (!\Mux11~6_combout  & (\Mux11~1_combout )))) # (!cuifregS_0 & (((\Mux11~6_combout ))))

	.dataa(\Mux11~1_combout ),
	.datab(cuifregS_0),
	.datac(\Mux11~6_combout ),
	.datad(\Mux11~8_combout ),
	.cin(gnd),
	.combout(\Mux11~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~9 .lut_mask = 16'hF838;
defparam \Mux11~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N12
cycloneive_lcell_comb \Mux12~7 (
// Equation(s):
// \Mux12~7_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[23][19]~q ))) # (!cuifregS_2 & (\registerArray[19][19]~q ))))

	.dataa(\registerArray[19][19]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[23][19]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux12~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~7 .lut_mask = 16'hFC22;
defparam \Mux12~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N14
cycloneive_lcell_comb \Mux12~8 (
// Equation(s):
// \Mux12~8_combout  = (cuifregS_3 & ((\Mux12~7_combout  & (\registerArray[31][19]~q )) # (!\Mux12~7_combout  & ((\registerArray[27][19]~q ))))) # (!cuifregS_3 & (((\Mux12~7_combout ))))

	.dataa(\registerArray[31][19]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[27][19]~q ),
	.datad(\Mux12~7_combout ),
	.cin(gnd),
	.combout(\Mux12~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~8 .lut_mask = 16'hBBC0;
defparam \Mux12~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N28
cycloneive_lcell_comb \Mux12~2 (
// Equation(s):
// \Mux12~2_combout  = (cuifregS_3 & (((\registerArray[26][19]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[18][19]~q  & ((!cuifregS_2))))

	.dataa(\registerArray[18][19]~q ),
	.datab(\registerArray[26][19]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux12~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~2 .lut_mask = 16'hF0CA;
defparam \Mux12~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N10
cycloneive_lcell_comb \Mux12~3 (
// Equation(s):
// \Mux12~3_combout  = (cuifregS_2 & ((\Mux12~2_combout  & ((\registerArray[30][19]~q ))) # (!\Mux12~2_combout  & (\registerArray[22][19]~q )))) # (!cuifregS_2 & (((\Mux12~2_combout ))))

	.dataa(\registerArray[22][19]~q ),
	.datab(\registerArray[30][19]~q ),
	.datac(cuifregS_2),
	.datad(\Mux12~2_combout ),
	.cin(gnd),
	.combout(\Mux12~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~3 .lut_mask = 16'hCFA0;
defparam \Mux12~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N4
cycloneive_lcell_comb \Mux12~6 (
// Equation(s):
// \Mux12~6_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\Mux12~3_combout ))) # (!cuifregS_1 & (\Mux12~5_combout ))))

	.dataa(\Mux12~5_combout ),
	.datab(cuifregS_0),
	.datac(\Mux12~3_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux12~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~6 .lut_mask = 16'hFC22;
defparam \Mux12~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N24
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (cuifregS_2 & (((\registerArray[21][19]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[17][19]~q  & ((!cuifregS_3))))

	.dataa(\registerArray[17][19]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[21][19]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hCCE2;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N26
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// \Mux12~1_combout  = (cuifregS_3 & ((\Mux12~0_combout  & ((\registerArray[29][19]~q ))) # (!\Mux12~0_combout  & (\registerArray[25][19]~q )))) # (!cuifregS_3 & (((\Mux12~0_combout ))))

	.dataa(\registerArray[25][19]~q ),
	.datab(\registerArray[29][19]~q ),
	.datac(cuifregS_3),
	.datad(\Mux12~0_combout ),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hCFA0;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y43_N22
cycloneive_lcell_comb \Mux12~9 (
// Equation(s):
// \Mux12~9_combout  = (cuifregS_0 & ((\Mux12~6_combout  & (\Mux12~8_combout )) # (!\Mux12~6_combout  & ((\Mux12~1_combout ))))) # (!cuifregS_0 & (((\Mux12~6_combout ))))

	.dataa(\Mux12~8_combout ),
	.datab(cuifregS_0),
	.datac(\Mux12~6_combout ),
	.datad(\Mux12~1_combout ),
	.cin(gnd),
	.combout(\Mux12~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~9 .lut_mask = 16'hBCB0;
defparam \Mux12~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y37_N6
cycloneive_lcell_comb \registerArray[1][19]~feeder (
// Equation(s):
// \registerArray[1][19]~feeder_combout  = \Mux49~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux492),
	.cin(gnd),
	.combout(\registerArray[1][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[1][19]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[1][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y37_N7
dffeas \registerArray[1][19] (
	.clk(clk),
	.d(\registerArray[1][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~79_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[1][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[1][19] .is_wysiwyg = "true";
defparam \registerArray[1][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N14
cycloneive_lcell_comb \Mux12~14 (
// Equation(s):
// \Mux12~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][19]~q ))) # (!cuifregS_1 & (\registerArray[1][19]~q ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[1][19]~q ),
	.datac(cuifregS_1),
	.datad(\registerArray[3][19]~q ),
	.cin(gnd),
	.combout(\Mux12~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~14 .lut_mask = 16'hA808;
defparam \Mux12~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N20
cycloneive_lcell_comb \Mux12~15 (
// Equation(s):
// \Mux12~15_combout  = (\Mux12~14_combout ) # ((!cuifregS_0 & (cuifregS_1 & \registerArray[2][19]~q )))

	.dataa(cuifregS_0),
	.datab(cuifregS_1),
	.datac(\Mux12~14_combout ),
	.datad(\registerArray[2][19]~q ),
	.cin(gnd),
	.combout(\Mux12~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~15 .lut_mask = 16'hF4F0;
defparam \Mux12~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N14
cycloneive_lcell_comb \Mux12~12 (
// Equation(s):
// \Mux12~12_combout  = (cuifregS_0 & ((\registerArray[5][19]~q ) # ((cuifregS_1)))) # (!cuifregS_0 & (((\registerArray[4][19]~q  & !cuifregS_1))))

	.dataa(\registerArray[5][19]~q ),
	.datab(\registerArray[4][19]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux12~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~12 .lut_mask = 16'hF0AC;
defparam \Mux12~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N10
cycloneive_lcell_comb \Mux12~13 (
// Equation(s):
// \Mux12~13_combout  = (cuifregS_1 & ((\Mux12~12_combout  & (\registerArray[7][19]~q )) # (!\Mux12~12_combout  & ((\registerArray[6][19]~q ))))) # (!cuifregS_1 & (((\Mux12~12_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[7][19]~q ),
	.datac(\registerArray[6][19]~q ),
	.datad(\Mux12~12_combout ),
	.cin(gnd),
	.combout(\Mux12~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~13 .lut_mask = 16'hDDA0;
defparam \Mux12~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N10
cycloneive_lcell_comb \Mux12~16 (
// Equation(s):
// \Mux12~16_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\Mux12~13_combout ))) # (!cuifregS_2 & (\Mux12~15_combout ))))

	.dataa(cuifregS_3),
	.datab(\Mux12~15_combout ),
	.datac(cuifregS_2),
	.datad(\Mux12~13_combout ),
	.cin(gnd),
	.combout(\Mux12~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~16 .lut_mask = 16'hF4A4;
defparam \Mux12~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y39_N17
dffeas \registerArray[9][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~72_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[9][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[9][19] .is_wysiwyg = "true";
defparam \registerArray[9][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y39_N3
dffeas \registerArray[10][19] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux492),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][19] .is_wysiwyg = "true";
defparam \registerArray[10][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N2
cycloneive_lcell_comb \Mux12~10 (
// Equation(s):
// \Mux12~10_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][19]~q ))) # (!cuifregS_1 & (\registerArray[8][19]~q ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[8][19]~q ),
	.datac(\registerArray[10][19]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux12~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~10 .lut_mask = 16'hFA44;
defparam \Mux12~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N16
cycloneive_lcell_comb \Mux12~11 (
// Equation(s):
// \Mux12~11_combout  = (cuifregS_0 & ((\Mux12~10_combout  & (\registerArray[11][19]~q )) # (!\Mux12~10_combout  & ((\registerArray[9][19]~q ))))) # (!cuifregS_0 & (((\Mux12~10_combout ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[11][19]~q ),
	.datac(\registerArray[9][19]~q ),
	.datad(\Mux12~10_combout ),
	.cin(gnd),
	.combout(\Mux12~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~11 .lut_mask = 16'hDDA0;
defparam \Mux12~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N24
cycloneive_lcell_comb \Mux12~17 (
// Equation(s):
// \Mux12~17_combout  = (cuifregS_1 & (((cuifregS_0)))) # (!cuifregS_1 & ((cuifregS_0 & (\registerArray[13][19]~q )) # (!cuifregS_0 & ((\registerArray[12][19]~q )))))

	.dataa(\registerArray[13][19]~q ),
	.datab(\registerArray[12][19]~q ),
	.datac(cuifregS_1),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux12~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~17 .lut_mask = 16'hFA0C;
defparam \Mux12~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y43_N22
cycloneive_lcell_comb \Mux12~18 (
// Equation(s):
// \Mux12~18_combout  = (cuifregS_1 & ((\Mux12~17_combout  & (\registerArray[15][19]~q )) # (!\Mux12~17_combout  & ((\registerArray[14][19]~q ))))) # (!cuifregS_1 & (((\Mux12~17_combout ))))

	.dataa(\registerArray[15][19]~q ),
	.datab(\registerArray[14][19]~q ),
	.datac(cuifregS_1),
	.datad(\Mux12~17_combout ),
	.cin(gnd),
	.combout(\Mux12~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~18 .lut_mask = 16'hAFC0;
defparam \Mux12~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y43_N16
cycloneive_lcell_comb \Mux12~19 (
// Equation(s):
// \Mux12~19_combout  = (\Mux12~16_combout  & (((\Mux12~18_combout )) # (!cuifregS_3))) # (!\Mux12~16_combout  & (cuifregS_3 & (\Mux12~11_combout )))

	.dataa(\Mux12~16_combout ),
	.datab(cuifregS_3),
	.datac(\Mux12~11_combout ),
	.datad(\Mux12~18_combout ),
	.cin(gnd),
	.combout(\Mux12~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~19 .lut_mask = 16'hEA62;
defparam \Mux12~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N16
cycloneive_lcell_comb \registerArray[20][18]~feeder (
// Equation(s):
// \registerArray[20][18]~feeder_combout  = \Mux50~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux502),
	.cin(gnd),
	.combout(\registerArray[20][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[20][18]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[20][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y40_N17
dffeas \registerArray[20][18] (
	.clk(clk),
	.d(\registerArray[20][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][18] .is_wysiwyg = "true";
defparam \registerArray[20][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y40_N0
cycloneive_lcell_comb \Mux13~4 (
// Equation(s):
// \Mux13~4_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & (\registerArray[20][18]~q )) # (!cuifregS_2 & ((\registerArray[16][18]~q )))))

	.dataa(cuifregS_3),
	.datab(\registerArray[20][18]~q ),
	.datac(\registerArray[16][18]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux13~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~4 .lut_mask = 16'hEE50;
defparam \Mux13~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y41_N2
cycloneive_lcell_comb \Mux13~5 (
// Equation(s):
// \Mux13~5_combout  = (cuifregS_3 & ((\Mux13~4_combout  & (\registerArray[28][18]~q )) # (!\Mux13~4_combout  & ((\registerArray[24][18]~q ))))) # (!cuifregS_3 & (((\Mux13~4_combout ))))

	.dataa(\registerArray[28][18]~q ),
	.datab(cuifregS_3),
	.datac(\registerArray[24][18]~q ),
	.datad(\Mux13~4_combout ),
	.cin(gnd),
	.combout(\Mux13~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~5 .lut_mask = 16'hBBC0;
defparam \Mux13~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N26
cycloneive_lcell_comb \Mux13~6 (
// Equation(s):
// \Mux13~6_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\Mux13~3_combout )) # (!cuifregS_1 & ((\Mux13~5_combout )))))

	.dataa(\Mux13~3_combout ),
	.datab(cuifregS_0),
	.datac(cuifregS_1),
	.datad(\Mux13~5_combout ),
	.cin(gnd),
	.combout(\Mux13~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~6 .lut_mask = 16'hE3E0;
defparam \Mux13~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N20
cycloneive_lcell_comb \registerArray[23][18]~feeder (
// Equation(s):
// \registerArray[23][18]~feeder_combout  = \Mux50~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux502),
	.cin(gnd),
	.combout(\registerArray[23][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[23][18]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[23][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y42_N21
dffeas \registerArray[23][18] (
	.clk(clk),
	.d(\registerArray[23][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][18] .is_wysiwyg = "true";
defparam \registerArray[23][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N20
cycloneive_lcell_comb \Mux13~7 (
// Equation(s):
// \Mux13~7_combout  = (cuifregS_3 & ((\registerArray[27][18]~q ) # ((cuifregS_2)))) # (!cuifregS_3 & (((\registerArray[19][18]~q  & !cuifregS_2))))

	.dataa(\registerArray[27][18]~q ),
	.datab(\registerArray[19][18]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux13~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~7 .lut_mask = 16'hF0AC;
defparam \Mux13~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y39_N26
cycloneive_lcell_comb \Mux13~8 (
// Equation(s):
// \Mux13~8_combout  = (cuifregS_2 & ((\Mux13~7_combout  & ((\registerArray[31][18]~q ))) # (!\Mux13~7_combout  & (\registerArray[23][18]~q )))) # (!cuifregS_2 & (((\Mux13~7_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[23][18]~q ),
	.datac(\registerArray[31][18]~q ),
	.datad(\Mux13~7_combout ),
	.cin(gnd),
	.combout(\Mux13~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~8 .lut_mask = 16'hF588;
defparam \Mux13~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y41_N26
cycloneive_lcell_comb \registerArray[17][18]~feeder (
// Equation(s):
// \registerArray[17][18]~feeder_combout  = \Mux50~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux502),
	.cin(gnd),
	.combout(\registerArray[17][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[17][18]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[17][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y41_N27
dffeas \registerArray[17][18] (
	.clk(clk),
	.d(\registerArray[17][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][18] .is_wysiwyg = "true";
defparam \registerArray[17][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N24
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// \Mux13~0_combout  = (cuifregS_3 & ((\registerArray[25][18]~q ) # ((cuifregS_2)))) # (!cuifregS_3 & (((\registerArray[17][18]~q  & !cuifregS_2))))

	.dataa(\registerArray[25][18]~q ),
	.datab(\registerArray[17][18]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hF0AC;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y41_N2
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// \Mux13~1_combout  = (cuifregS_2 & ((\Mux13~0_combout  & ((\registerArray[29][18]~q ))) # (!\Mux13~0_combout  & (\registerArray[21][18]~q )))) # (!cuifregS_2 & (((\Mux13~0_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[21][18]~q ),
	.datac(\registerArray[29][18]~q ),
	.datad(\Mux13~0_combout ),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'hF588;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N16
cycloneive_lcell_comb \Mux13~9 (
// Equation(s):
// \Mux13~9_combout  = (\Mux13~6_combout  & (((\Mux13~8_combout )) # (!cuifregS_0))) # (!\Mux13~6_combout  & (cuifregS_0 & ((\Mux13~1_combout ))))

	.dataa(\Mux13~6_combout ),
	.datab(cuifregS_0),
	.datac(\Mux13~8_combout ),
	.datad(\Mux13~1_combout ),
	.cin(gnd),
	.combout(\Mux13~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~9 .lut_mask = 16'hE6A2;
defparam \Mux13~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N22
cycloneive_lcell_comb \Mux13~17 (
// Equation(s):
// \Mux13~17_combout  = (cuifregS_0 & ((\registerArray[13][18]~q ) # ((cuifregS_1)))) # (!cuifregS_0 & (((\registerArray[12][18]~q  & !cuifregS_1))))

	.dataa(\registerArray[13][18]~q ),
	.datab(\registerArray[12][18]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux13~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~17 .lut_mask = 16'hF0AC;
defparam \Mux13~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y42_N24
cycloneive_lcell_comb \Mux13~18 (
// Equation(s):
// \Mux13~18_combout  = (\Mux13~17_combout  & (((\registerArray[15][18]~q ) # (!cuifregS_1)))) # (!\Mux13~17_combout  & (\registerArray[14][18]~q  & ((cuifregS_1))))

	.dataa(\registerArray[14][18]~q ),
	.datab(\registerArray[15][18]~q ),
	.datac(\Mux13~17_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux13~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~18 .lut_mask = 16'hCAF0;
defparam \Mux13~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N1
dffeas \registerArray[6][18] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux502),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][18] .is_wysiwyg = "true";
defparam \registerArray[6][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N6
cycloneive_lcell_comb \Mux13~10 (
// Equation(s):
// \Mux13~10_combout  = (cuifregS_0 & ((\registerArray[5][18]~q ) # ((cuifregS_1)))) # (!cuifregS_0 & (((\registerArray[4][18]~q  & !cuifregS_1))))

	.dataa(\registerArray[5][18]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[4][18]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux13~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~10 .lut_mask = 16'hCCB8;
defparam \Mux13~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N0
cycloneive_lcell_comb \Mux13~11 (
// Equation(s):
// \Mux13~11_combout  = (cuifregS_1 & ((\Mux13~10_combout  & (\registerArray[7][18]~q )) # (!\Mux13~10_combout  & ((\registerArray[6][18]~q ))))) # (!cuifregS_1 & (((\Mux13~10_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[7][18]~q ),
	.datac(\registerArray[6][18]~q ),
	.datad(\Mux13~10_combout ),
	.cin(gnd),
	.combout(\Mux13~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~11 .lut_mask = 16'hDDA0;
defparam \Mux13~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N10
cycloneive_lcell_comb \Mux13~14 (
// Equation(s):
// \Mux13~14_combout  = (cuifregS_0 & ((cuifregS_1 & (\registerArray[3][18]~q )) # (!cuifregS_1 & ((\registerArray[1][18]~q )))))

	.dataa(\registerArray[3][18]~q ),
	.datab(cuifregS_1),
	.datac(cuifregS_0),
	.datad(\registerArray[1][18]~q ),
	.cin(gnd),
	.combout(\Mux13~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~14 .lut_mask = 16'hB080;
defparam \Mux13~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N8
cycloneive_lcell_comb \Mux13~15 (
// Equation(s):
// \Mux13~15_combout  = (\Mux13~14_combout ) # ((\registerArray[2][18]~q  & (!cuifregS_0 & cuifregS_1)))

	.dataa(\registerArray[2][18]~q ),
	.datab(cuifregS_0),
	.datac(cuifregS_1),
	.datad(\Mux13~14_combout ),
	.cin(gnd),
	.combout(\Mux13~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~15 .lut_mask = 16'hFF20;
defparam \Mux13~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N18
cycloneive_lcell_comb \registerArray[10][18]~feeder (
// Equation(s):
// \registerArray[10][18]~feeder_combout  = \Mux50~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux502),
	.cin(gnd),
	.combout(\registerArray[10][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[10][18]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[10][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y41_N19
dffeas \registerArray[10][18] (
	.clk(clk),
	.d(\registerArray[10][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~73_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[10][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[10][18] .is_wysiwyg = "true";
defparam \registerArray[10][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N0
cycloneive_lcell_comb \Mux13~12 (
// Equation(s):
// \Mux13~12_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\registerArray[10][18]~q ))) # (!cuifregS_1 & (\registerArray[8][18]~q ))))

	.dataa(\registerArray[8][18]~q ),
	.datab(\registerArray[10][18]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux13~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~12 .lut_mask = 16'hFC0A;
defparam \Mux13~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y41_N10
cycloneive_lcell_comb \Mux13~13 (
// Equation(s):
// \Mux13~13_combout  = (cuifregS_0 & ((\Mux13~12_combout  & ((\registerArray[11][18]~q ))) # (!\Mux13~12_combout  & (\registerArray[9][18]~q )))) # (!cuifregS_0 & (((\Mux13~12_combout ))))

	.dataa(\registerArray[9][18]~q ),
	.datab(\registerArray[11][18]~q ),
	.datac(cuifregS_0),
	.datad(\Mux13~12_combout ),
	.cin(gnd),
	.combout(\Mux13~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~13 .lut_mask = 16'hCFA0;
defparam \Mux13~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N6
cycloneive_lcell_comb \Mux13~16 (
// Equation(s):
// \Mux13~16_combout  = (cuifregS_3 & ((cuifregS_2) # ((\Mux13~13_combout )))) # (!cuifregS_3 & (!cuifregS_2 & (\Mux13~15_combout )))

	.dataa(cuifregS_3),
	.datab(cuifregS_2),
	.datac(\Mux13~15_combout ),
	.datad(\Mux13~13_combout ),
	.cin(gnd),
	.combout(\Mux13~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~16 .lut_mask = 16'hBA98;
defparam \Mux13~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y42_N28
cycloneive_lcell_comb \Mux13~19 (
// Equation(s):
// \Mux13~19_combout  = (cuifregS_2 & ((\Mux13~16_combout  & (\Mux13~18_combout )) # (!\Mux13~16_combout  & ((\Mux13~11_combout ))))) # (!cuifregS_2 & (((\Mux13~16_combout ))))

	.dataa(\Mux13~18_combout ),
	.datab(cuifregS_2),
	.datac(\Mux13~11_combout ),
	.datad(\Mux13~16_combout ),
	.cin(gnd),
	.combout(\Mux13~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~19 .lut_mask = 16'hBBC0;
defparam \Mux13~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N14
cycloneive_lcell_comb \registerArray[13][17]~feeder (
// Equation(s):
// \registerArray[13][17]~feeder_combout  = \Mux51~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux512),
	.cin(gnd),
	.combout(\registerArray[13][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[13][17]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[13][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N15
dffeas \registerArray[13][17] (
	.clk(clk),
	.d(\registerArray[13][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~82_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[13][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[13][17] .is_wysiwyg = "true";
defparam \registerArray[13][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N4
cycloneive_lcell_comb \Mux14~17 (
// Equation(s):
// \Mux14~17_combout  = (cuifregS_0 & (((\registerArray[13][17]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[12][17]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[12][17]~q ),
	.datab(\registerArray[13][17]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux14~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~17 .lut_mask = 16'hF0CA;
defparam \Mux14~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N6
cycloneive_lcell_comb \Mux14~18 (
// Equation(s):
// \Mux14~18_combout  = (\Mux14~17_combout  & ((\registerArray[15][17]~q ) # ((!cuifregS_1)))) # (!\Mux14~17_combout  & (((\registerArray[14][17]~q  & cuifregS_1))))

	.dataa(\registerArray[15][17]~q ),
	.datab(\registerArray[14][17]~q ),
	.datac(\Mux14~17_combout ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux14~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~18 .lut_mask = 16'hACF0;
defparam \Mux14~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y39_N4
cycloneive_lcell_comb \Mux14~11 (
// Equation(s):
// \Mux14~11_combout  = (\Mux14~10_combout  & ((\registerArray[11][17]~q ) # ((!cuifregS_0)))) # (!\Mux14~10_combout  & (((\registerArray[9][17]~q  & cuifregS_0))))

	.dataa(\Mux14~10_combout ),
	.datab(\registerArray[11][17]~q ),
	.datac(\registerArray[9][17]~q ),
	.datad(cuifregS_0),
	.cin(gnd),
	.combout(\Mux14~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~11 .lut_mask = 16'hD8AA;
defparam \Mux14~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y37_N13
dffeas \registerArray[3][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~78_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[3][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[3][17] .is_wysiwyg = "true";
defparam \registerArray[3][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y37_N12
cycloneive_lcell_comb \Mux14~14 (
// Equation(s):
// \Mux14~14_combout  = (cuifregS_0 & ((cuifregS_1 & ((\registerArray[3][17]~q ))) # (!cuifregS_1 & (\registerArray[1][17]~q ))))

	.dataa(\registerArray[1][17]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[3][17]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux14~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~14 .lut_mask = 16'hC088;
defparam \Mux14~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N4
cycloneive_lcell_comb \Mux14~15 (
// Equation(s):
// \Mux14~15_combout  = (\Mux14~14_combout ) # ((\registerArray[2][17]~q  & (!cuifregS_0 & cuifregS_1)))

	.dataa(\registerArray[2][17]~q ),
	.datab(cuifregS_0),
	.datac(cuifregS_1),
	.datad(\Mux14~14_combout ),
	.cin(gnd),
	.combout(\Mux14~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~15 .lut_mask = 16'hFF20;
defparam \Mux14~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N10
cycloneive_lcell_comb \registerArray[4][17]~feeder (
// Equation(s):
// \registerArray[4][17]~feeder_combout  = \Mux51~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux512),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[4][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[4][17]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[4][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N11
dffeas \registerArray[4][17] (
	.clk(clk),
	.d(\registerArray[4][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~59_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[4][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[4][17] .is_wysiwyg = "true";
defparam \registerArray[4][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N4
cycloneive_lcell_comb \Mux14~12 (
// Equation(s):
// \Mux14~12_combout  = (cuifregS_0 & (((\registerArray[5][17]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[4][17]~q  & ((!cuifregS_1))))

	.dataa(cuifregS_0),
	.datab(\registerArray[4][17]~q ),
	.datac(\registerArray[5][17]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux14~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~12 .lut_mask = 16'hAAE4;
defparam \Mux14~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y38_N24
cycloneive_lcell_comb \Mux14~13 (
// Equation(s):
// \Mux14~13_combout  = (cuifregS_1 & ((\Mux14~12_combout  & (\registerArray[7][17]~q )) # (!\Mux14~12_combout  & ((\registerArray[6][17]~q ))))) # (!cuifregS_1 & (((\Mux14~12_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[7][17]~q ),
	.datac(\registerArray[6][17]~q ),
	.datad(\Mux14~12_combout ),
	.cin(gnd),
	.combout(\Mux14~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~13 .lut_mask = 16'hDDA0;
defparam \Mux14~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N2
cycloneive_lcell_comb \Mux14~16 (
// Equation(s):
// \Mux14~16_combout  = (cuifregS_3 & (cuifregS_2)) # (!cuifregS_3 & ((cuifregS_2 & ((\Mux14~13_combout ))) # (!cuifregS_2 & (\Mux14~15_combout ))))

	.dataa(cuifregS_3),
	.datab(cuifregS_2),
	.datac(\Mux14~15_combout ),
	.datad(\Mux14~13_combout ),
	.cin(gnd),
	.combout(\Mux14~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~16 .lut_mask = 16'hDC98;
defparam \Mux14~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N8
cycloneive_lcell_comb \Mux14~19 (
// Equation(s):
// \Mux14~19_combout  = (cuifregS_3 & ((\Mux14~16_combout  & (\Mux14~18_combout )) # (!\Mux14~16_combout  & ((\Mux14~11_combout ))))) # (!cuifregS_3 & (((\Mux14~16_combout ))))

	.dataa(\Mux14~18_combout ),
	.datab(cuifregS_3),
	.datac(\Mux14~11_combout ),
	.datad(\Mux14~16_combout ),
	.cin(gnd),
	.combout(\Mux14~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~19 .lut_mask = 16'hBBC0;
defparam \Mux14~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y41_N19
dffeas \registerArray[27][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~68_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[27][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[27][17] .is_wysiwyg = "true";
defparam \registerArray[27][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y41_N2
cycloneive_lcell_comb \Mux14~7 (
// Equation(s):
// \Mux14~7_combout  = (cuifregS_2 & (((\registerArray[23][17]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[19][17]~q  & ((!cuifregS_3))))

	.dataa(cuifregS_2),
	.datab(\registerArray[19][17]~q ),
	.datac(\registerArray[23][17]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux14~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~7 .lut_mask = 16'hAAE4;
defparam \Mux14~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y41_N30
cycloneive_lcell_comb \Mux14~8 (
// Equation(s):
// \Mux14~8_combout  = (cuifregS_3 & ((\Mux14~7_combout  & (\registerArray[31][17]~q )) # (!\Mux14~7_combout  & ((\registerArray[27][17]~q ))))) # (!cuifregS_3 & (((\Mux14~7_combout ))))

	.dataa(\registerArray[31][17]~q ),
	.datab(\registerArray[27][17]~q ),
	.datac(cuifregS_3),
	.datad(\Mux14~7_combout ),
	.cin(gnd),
	.combout(\Mux14~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~8 .lut_mask = 16'hAFC0;
defparam \Mux14~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y37_N30
cycloneive_lcell_comb \registerArray[17][17]~feeder (
// Equation(s):
// \registerArray[17][17]~feeder_combout  = \Mux51~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux512),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[17][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[17][17]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[17][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y37_N31
dffeas \registerArray[17][17] (
	.clk(clk),
	.d(\registerArray[17][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~53_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[17][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[17][17] .is_wysiwyg = "true";
defparam \registerArray[17][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N24
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// \Mux14~0_combout  = (cuifregS_3 & (((cuifregS_2)))) # (!cuifregS_3 & ((cuifregS_2 & ((\registerArray[21][17]~q ))) # (!cuifregS_2 & (\registerArray[17][17]~q ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[17][17]~q ),
	.datac(\registerArray[21][17]~q ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hFA44;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y41_N6
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// \Mux14~1_combout  = (cuifregS_3 & ((\Mux14~0_combout  & (\registerArray[29][17]~q )) # (!\Mux14~0_combout  & ((\registerArray[25][17]~q ))))) # (!cuifregS_3 & (((\Mux14~0_combout ))))

	.dataa(cuifregS_3),
	.datab(\registerArray[29][17]~q ),
	.datac(\registerArray[25][17]~q ),
	.datad(\Mux14~0_combout ),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hDDA0;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y42_N11
dffeas \registerArray[22][17] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux512),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~62_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[22][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[22][17] .is_wysiwyg = "true";
defparam \registerArray[22][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N0
cycloneive_lcell_comb \registerArray[26][17]~feeder (
// Equation(s):
// \registerArray[26][17]~feeder_combout  = \Mux51~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux512),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[26][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[26][17]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[26][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N1
dffeas \registerArray[26][17] (
	.clk(clk),
	.d(\registerArray[26][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][17] .is_wysiwyg = "true";
defparam \registerArray[26][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N22
cycloneive_lcell_comb \Mux14~2 (
// Equation(s):
// \Mux14~2_combout  = (cuifregS_3 & (((\registerArray[26][17]~q ) # (cuifregS_2)))) # (!cuifregS_3 & (\registerArray[18][17]~q  & ((!cuifregS_2))))

	.dataa(\registerArray[18][17]~q ),
	.datab(\registerArray[26][17]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux14~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~2 .lut_mask = 16'hF0CA;
defparam \Mux14~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y42_N10
cycloneive_lcell_comb \Mux14~3 (
// Equation(s):
// \Mux14~3_combout  = (cuifregS_2 & ((\Mux14~2_combout  & (\registerArray[30][17]~q )) # (!\Mux14~2_combout  & ((\registerArray[22][17]~q ))))) # (!cuifregS_2 & (((\Mux14~2_combout ))))

	.dataa(\registerArray[30][17]~q ),
	.datab(cuifregS_2),
	.datac(\registerArray[22][17]~q ),
	.datad(\Mux14~2_combout ),
	.cin(gnd),
	.combout(\Mux14~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~3 .lut_mask = 16'hBBC0;
defparam \Mux14~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N28
cycloneive_lcell_comb \Mux14~6 (
// Equation(s):
// \Mux14~6_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & ((\Mux14~3_combout ))) # (!cuifregS_1 & (\Mux14~5_combout ))))

	.dataa(\Mux14~5_combout ),
	.datab(cuifregS_0),
	.datac(cuifregS_1),
	.datad(\Mux14~3_combout ),
	.cin(gnd),
	.combout(\Mux14~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~6 .lut_mask = 16'hF2C2;
defparam \Mux14~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y40_N10
cycloneive_lcell_comb \Mux14~9 (
// Equation(s):
// \Mux14~9_combout  = (cuifregS_0 & ((\Mux14~6_combout  & (\Mux14~8_combout )) # (!\Mux14~6_combout  & ((\Mux14~1_combout ))))) # (!cuifregS_0 & (((\Mux14~6_combout ))))

	.dataa(\Mux14~8_combout ),
	.datab(cuifregS_0),
	.datac(\Mux14~1_combout ),
	.datad(\Mux14~6_combout ),
	.cin(gnd),
	.combout(\Mux14~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~9 .lut_mask = 16'hBBC0;
defparam \Mux14~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y34_N13
dffeas \registerArray[6][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~76_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[6][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[6][0] .is_wysiwyg = "true";
defparam \registerArray[6][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N24
cycloneive_lcell_comb \registerArray[5][0]~feeder (
// Equation(s):
// \registerArray[5][0]~feeder_combout  = \Mux68~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux68),
	.cin(gnd),
	.combout(\registerArray[5][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[5][0]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[5][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N25
dffeas \registerArray[5][0] (
	.clk(clk),
	.d(\registerArray[5][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~58_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[5][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[5][0] .is_wysiwyg = "true";
defparam \registerArray[5][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N16
cycloneive_lcell_comb \Mux31~10 (
// Equation(s):
// \Mux31~10_combout  = (cuifregS_0 & (((\registerArray[5][0]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[4][0]~q  & ((!cuifregS_1))))

	.dataa(\registerArray[4][0]~q ),
	.datab(\registerArray[5][0]~q ),
	.datac(cuifregS_0),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux31~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~10 .lut_mask = 16'hF0CA;
defparam \Mux31~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N12
cycloneive_lcell_comb \Mux31~11 (
// Equation(s):
// \Mux31~11_combout  = (cuifregS_1 & ((\Mux31~10_combout  & (\registerArray[7][0]~q )) # (!\Mux31~10_combout  & ((\registerArray[6][0]~q ))))) # (!cuifregS_1 & (((\Mux31~10_combout ))))

	.dataa(cuifregS_1),
	.datab(\registerArray[7][0]~q ),
	.datac(\registerArray[6][0]~q ),
	.datad(\Mux31~10_combout ),
	.cin(gnd),
	.combout(\Mux31~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~11 .lut_mask = 16'hDDA0;
defparam \Mux31~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y35_N23
dffeas \registerArray[8][0] (
	.clk(clk),
	.d(gnd),
	.asdata(Mux68),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~74_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[8][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[8][0] .is_wysiwyg = "true";
defparam \registerArray[8][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y35_N22
cycloneive_lcell_comb \Mux31~12 (
// Equation(s):
// \Mux31~12_combout  = (cuifregS_0 & (((cuifregS_1)))) # (!cuifregS_0 & ((cuifregS_1 & (\registerArray[10][0]~q )) # (!cuifregS_1 & ((\registerArray[8][0]~q )))))

	.dataa(\registerArray[10][0]~q ),
	.datab(cuifregS_0),
	.datac(\registerArray[8][0]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux31~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~12 .lut_mask = 16'hEE30;
defparam \Mux31~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N22
cycloneive_lcell_comb \Mux31~13 (
// Equation(s):
// \Mux31~13_combout  = (cuifregS_0 & ((\Mux31~12_combout  & ((\registerArray[11][0]~q ))) # (!\Mux31~12_combout  & (\registerArray[9][0]~q )))) # (!cuifregS_0 & (((\Mux31~12_combout ))))

	.dataa(cuifregS_0),
	.datab(\registerArray[9][0]~q ),
	.datac(\registerArray[11][0]~q ),
	.datad(\Mux31~12_combout ),
	.cin(gnd),
	.combout(\Mux31~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~13 .lut_mask = 16'hF588;
defparam \Mux31~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y37_N12
cycloneive_lcell_comb \Mux31~14 (
// Equation(s):
// \Mux31~14_combout  = (cuifregS_0 & ((cuifregS_1 & (\registerArray[3][0]~q )) # (!cuifregS_1 & ((\registerArray[1][0]~q )))))

	.dataa(cuifregS_1),
	.datab(cuifregS_0),
	.datac(\registerArray[3][0]~q ),
	.datad(\registerArray[1][0]~q ),
	.cin(gnd),
	.combout(\Mux31~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~14 .lut_mask = 16'hC480;
defparam \Mux31~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N12
cycloneive_lcell_comb \Mux31~15 (
// Equation(s):
// \Mux31~15_combout  = (\Mux31~14_combout ) # ((!cuifregS_0 & (cuifregS_1 & \registerArray[2][0]~q )))

	.dataa(cuifregS_0),
	.datab(cuifregS_1),
	.datac(\registerArray[2][0]~q ),
	.datad(\Mux31~14_combout ),
	.cin(gnd),
	.combout(\Mux31~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~15 .lut_mask = 16'hFF40;
defparam \Mux31~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N22
cycloneive_lcell_comb \Mux31~16 (
// Equation(s):
// \Mux31~16_combout  = (cuifregS_2 & (cuifregS_3)) # (!cuifregS_2 & ((cuifregS_3 & (\Mux31~13_combout )) # (!cuifregS_3 & ((\Mux31~15_combout )))))

	.dataa(cuifregS_2),
	.datab(cuifregS_3),
	.datac(\Mux31~13_combout ),
	.datad(\Mux31~15_combout ),
	.cin(gnd),
	.combout(\Mux31~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~16 .lut_mask = 16'hD9C8;
defparam \Mux31~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y36_N28
cycloneive_lcell_comb \Mux31~17 (
// Equation(s):
// \Mux31~17_combout  = (cuifregS_0 & (((\registerArray[13][0]~q ) # (cuifregS_1)))) # (!cuifregS_0 & (\registerArray[12][0]~q  & ((!cuifregS_1))))

	.dataa(cuifregS_0),
	.datab(\registerArray[12][0]~q ),
	.datac(\registerArray[13][0]~q ),
	.datad(cuifregS_1),
	.cin(gnd),
	.combout(\Mux31~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~17 .lut_mask = 16'hAAE4;
defparam \Mux31~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N26
cycloneive_lcell_comb \Mux31~18 (
// Equation(s):
// \Mux31~18_combout  = (cuifregS_1 & ((\Mux31~17_combout  & ((\registerArray[15][0]~q ))) # (!\Mux31~17_combout  & (\registerArray[14][0]~q )))) # (!cuifregS_1 & (((\Mux31~17_combout ))))

	.dataa(\registerArray[14][0]~q ),
	.datab(\registerArray[15][0]~q ),
	.datac(cuifregS_1),
	.datad(\Mux31~17_combout ),
	.cin(gnd),
	.combout(\Mux31~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~18 .lut_mask = 16'hCFA0;
defparam \Mux31~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N4
cycloneive_lcell_comb \Mux31~19 (
// Equation(s):
// \Mux31~19_combout  = (cuifregS_2 & ((\Mux31~16_combout  & ((\Mux31~18_combout ))) # (!\Mux31~16_combout  & (\Mux31~11_combout )))) # (!cuifregS_2 & (((\Mux31~16_combout ))))

	.dataa(cuifregS_2),
	.datab(\Mux31~11_combout ),
	.datac(\Mux31~16_combout ),
	.datad(\Mux31~18_combout ),
	.cin(gnd),
	.combout(\Mux31~19_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~19 .lut_mask = 16'hF858;
defparam \Mux31~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N18
cycloneive_lcell_comb \registerArray[23][0]~feeder (
// Equation(s):
// \registerArray[23][0]~feeder_combout  = \Mux68~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux68),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[23][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[23][0]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[23][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y40_N19
dffeas \registerArray[23][0] (
	.clk(clk),
	.d(\registerArray[23][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~69_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[23][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[23][0] .is_wysiwyg = "true";
defparam \registerArray[23][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N20
cycloneive_lcell_comb \Mux31~7 (
// Equation(s):
// \Mux31~7_combout  = (cuifregS_2 & (((cuifregS_3)))) # (!cuifregS_2 & ((cuifregS_3 & ((\registerArray[27][0]~q ))) # (!cuifregS_3 & (\registerArray[19][0]~q ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[19][0]~q ),
	.datac(\registerArray[27][0]~q ),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux31~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~7 .lut_mask = 16'hFA44;
defparam \Mux31~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y40_N12
cycloneive_lcell_comb \Mux31~8 (
// Equation(s):
// \Mux31~8_combout  = (cuifregS_2 & ((\Mux31~7_combout  & ((\registerArray[31][0]~q ))) # (!\Mux31~7_combout  & (\registerArray[23][0]~q )))) # (!cuifregS_2 & (((\Mux31~7_combout ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[23][0]~q ),
	.datac(\registerArray[31][0]~q ),
	.datad(\Mux31~7_combout ),
	.cin(gnd),
	.combout(\Mux31~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~8 .lut_mask = 16'hF588;
defparam \Mux31~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N8
cycloneive_lcell_comb \registerArray[20][0]~feeder (
// Equation(s):
// \registerArray[20][0]~feeder_combout  = \Mux68~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux68),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[20][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[20][0]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[20][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y39_N9
dffeas \registerArray[20][0] (
	.clk(clk),
	.d(\registerArray[20][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~55_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[20][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[20][0] .is_wysiwyg = "true";
defparam \registerArray[20][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y39_N10
cycloneive_lcell_comb \Mux31~4 (
// Equation(s):
// \Mux31~4_combout  = (cuifregS_2 & ((\registerArray[20][0]~q ) # ((cuifregS_3)))) # (!cuifregS_2 & (((!cuifregS_3 & \registerArray[16][0]~q ))))

	.dataa(cuifregS_2),
	.datab(\registerArray[20][0]~q ),
	.datac(cuifregS_3),
	.datad(\registerArray[16][0]~q ),
	.cin(gnd),
	.combout(\Mux31~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~4 .lut_mask = 16'hADA8;
defparam \Mux31~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N14
cycloneive_lcell_comb \Mux31~5 (
// Equation(s):
// \Mux31~5_combout  = (cuifregS_3 & ((\Mux31~4_combout  & ((\registerArray[28][0]~q ))) # (!\Mux31~4_combout  & (\registerArray[24][0]~q )))) # (!cuifregS_3 & (((\Mux31~4_combout ))))

	.dataa(\registerArray[24][0]~q ),
	.datab(\registerArray[28][0]~q ),
	.datac(cuifregS_3),
	.datad(\Mux31~4_combout ),
	.cin(gnd),
	.combout(\Mux31~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~5 .lut_mask = 16'hCFA0;
defparam \Mux31~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y40_N26
cycloneive_lcell_comb \Mux31~2 (
// Equation(s):
// \Mux31~2_combout  = (cuifregS_2 & (((\registerArray[22][0]~q ) # (cuifregS_3)))) # (!cuifregS_2 & (\registerArray[18][0]~q  & ((!cuifregS_3))))

	.dataa(\registerArray[18][0]~q ),
	.datab(\registerArray[22][0]~q ),
	.datac(cuifregS_2),
	.datad(cuifregS_3),
	.cin(gnd),
	.combout(\Mux31~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~2 .lut_mask = 16'hF0CA;
defparam \Mux31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N8
cycloneive_lcell_comb \registerArray[26][0]~feeder (
// Equation(s):
// \registerArray[26][0]~feeder_combout  = \Mux68~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux68),
	.datad(gnd),
	.cin(gnd),
	.combout(\registerArray[26][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[26][0]~feeder .lut_mask = 16'hF0F0;
defparam \registerArray[26][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y40_N9
dffeas \registerArray[26][0] (
	.clk(clk),
	.d(\registerArray[26][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~63_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[26][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[26][0] .is_wysiwyg = "true";
defparam \registerArray[26][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y40_N4
cycloneive_lcell_comb \Mux31~3 (
// Equation(s):
// \Mux31~3_combout  = (cuifregS_3 & ((\Mux31~2_combout  & (\registerArray[30][0]~q )) # (!\Mux31~2_combout  & ((\registerArray[26][0]~q ))))) # (!cuifregS_3 & (((\Mux31~2_combout ))))

	.dataa(\registerArray[30][0]~q ),
	.datab(cuifregS_3),
	.datac(\Mux31~2_combout ),
	.datad(\registerArray[26][0]~q ),
	.cin(gnd),
	.combout(\Mux31~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~3 .lut_mask = 16'hBCB0;
defparam \Mux31~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N8
cycloneive_lcell_comb \Mux31~6 (
// Equation(s):
// \Mux31~6_combout  = (cuifregS_0 & (cuifregS_1)) # (!cuifregS_0 & ((cuifregS_1 & ((\Mux31~3_combout ))) # (!cuifregS_1 & (\Mux31~5_combout ))))

	.dataa(cuifregS_0),
	.datab(cuifregS_1),
	.datac(\Mux31~5_combout ),
	.datad(\Mux31~3_combout ),
	.cin(gnd),
	.combout(\Mux31~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~6 .lut_mask = 16'hDC98;
defparam \Mux31~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y36_N20
cycloneive_lcell_comb \registerArray[21][0]~feeder (
// Equation(s):
// \registerArray[21][0]~feeder_combout  = \Mux68~1_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux68),
	.cin(gnd),
	.combout(\registerArray[21][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \registerArray[21][0]~feeder .lut_mask = 16'hFF00;
defparam \registerArray[21][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y36_N21
dffeas \registerArray[21][0] (
	.clk(clk),
	.d(\registerArray[21][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(n_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~52_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\registerArray[21][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \registerArray[21][0] .is_wysiwyg = "true";
defparam \registerArray[21][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N4
cycloneive_lcell_comb \Mux31~0 (
// Equation(s):
// \Mux31~0_combout  = (cuifregS_3 & ((\registerArray[25][0]~q ) # ((cuifregS_2)))) # (!cuifregS_3 & (((\registerArray[17][0]~q  & !cuifregS_2))))

	.dataa(\registerArray[25][0]~q ),
	.datab(\registerArray[17][0]~q ),
	.datac(cuifregS_3),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~0 .lut_mask = 16'hF0AC;
defparam \Mux31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y40_N26
cycloneive_lcell_comb \Mux31~1 (
// Equation(s):
// \Mux31~1_combout  = (\Mux31~0_combout  & ((\registerArray[29][0]~q ) # ((!cuifregS_2)))) # (!\Mux31~0_combout  & (((\registerArray[21][0]~q  & cuifregS_2))))

	.dataa(\registerArray[29][0]~q ),
	.datab(\registerArray[21][0]~q ),
	.datac(\Mux31~0_combout ),
	.datad(cuifregS_2),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~1 .lut_mask = 16'hACF0;
defparam \Mux31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y40_N10
cycloneive_lcell_comb \Mux31~9 (
// Equation(s):
// \Mux31~9_combout  = (cuifregS_0 & ((\Mux31~6_combout  & (\Mux31~8_combout )) # (!\Mux31~6_combout  & ((\Mux31~1_combout ))))) # (!cuifregS_0 & (((\Mux31~6_combout ))))

	.dataa(cuifregS_0),
	.datab(\Mux31~8_combout ),
	.datac(\Mux31~6_combout ),
	.datad(\Mux31~1_combout ),
	.cin(gnd),
	.combout(\Mux31~9_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~9 .lut_mask = 16'hDAD0;
defparam \Mux31~9 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module request_unit (
	ruifdmemREN,
	ruifdmemWEN,
	always1,
	dcifimemload_30,
	dcifimemload_31,
	dcifimemload_29,
	Equal2,
	dcifdhit,
	CPUCLK,
	nRST,
	devpor,
	devclrn,
	devoe);
output 	ruifdmemREN;
output 	ruifdmemWEN;
input 	always1;
input 	dcifimemload_30;
input 	dcifimemload_31;
input 	dcifimemload_29;
input 	Equal2;
input 	dcifdhit;
input 	CPUCLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \dmemREN~0_combout ;
wire \dmemREN~1_combout ;
wire \dmemWEN~0_combout ;


// Location: FF_X59_Y36_N25
dffeas \ruif.dmemREN (
	.clk(CPUCLK),
	.d(\dmemREN~1_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ruifdmemREN),
	.prn(vcc));
// synopsys translate_off
defparam \ruif.dmemREN .is_wysiwyg = "true";
defparam \ruif.dmemREN .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y36_N15
dffeas \ruif.dmemWEN (
	.clk(CPUCLK),
	.d(\dmemWEN~0_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always1),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ruifdmemWEN),
	.prn(vcc));
// synopsys translate_off
defparam \ruif.dmemWEN .is_wysiwyg = "true";
defparam \ruif.dmemWEN .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N28
cycloneive_lcell_comb \dmemREN~0 (
// Equation(s):
// \dmemREN~0_combout  = (dcifimemload_31 & (Equal21 & (dcifdhit & !dcifimemload_30)))

	.dataa(dcifimemload_31),
	.datab(Equal2),
	.datac(dcifdhit),
	.datad(dcifimemload_30),
	.cin(gnd),
	.combout(\dmemREN~0_combout ),
	.cout());
// synopsys translate_off
defparam \dmemREN~0 .lut_mask = 16'h0080;
defparam \dmemREN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N24
cycloneive_lcell_comb \dmemREN~1 (
// Equation(s):
// \dmemREN~1_combout  = (!dcifimemload_29 & \dmemREN~0_combout )

	.dataa(gnd),
	.datab(dcifimemload_29),
	.datac(gnd),
	.datad(\dmemREN~0_combout ),
	.cin(gnd),
	.combout(\dmemREN~1_combout ),
	.cout());
// synopsys translate_off
defparam \dmemREN~1 .lut_mask = 16'h3300;
defparam \dmemREN~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y36_N14
cycloneive_lcell_comb \dmemWEN~0 (
// Equation(s):
// \dmemWEN~0_combout  = (dcifimemload_29 & \dmemREN~0_combout )

	.dataa(gnd),
	.datab(dcifimemload_29),
	.datac(gnd),
	.datad(\dmemREN~0_combout ),
	.cin(gnd),
	.combout(\dmemWEN~0_combout ),
	.cout());
// synopsys translate_off
defparam \dmemWEN~0 .lut_mask = 16'hCC00;
defparam \dmemWEN~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module memory_control (
	ruifdmemREN,
	ruifdmemWEN,
	iwait,
	devpor,
	devclrn,
	devoe);
input 	ruifdmemREN;
input 	ruifdmemWEN;
output 	iwait;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X59_Y35_N2
cycloneive_lcell_comb \iwait~0 (
// Equation(s):
// iwait = (ruifdmemWEN) # (ruifdmemREN)

	.dataa(ruifdmemWEN),
	.datab(gnd),
	.datac(gnd),
	.datad(ruifdmemREN),
	.cin(gnd),
	.combout(iwait),
	.cout());
// synopsys translate_off
defparam \iwait~0 .lut_mask = 16'hFFAA;
defparam \iwait~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule
