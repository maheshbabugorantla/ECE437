/*
	Mahesh Babu Gorantla
	mgorantl@purdue.edu

	Holds the Program Counter Logic Interface Signals
*/

`ifndef PC_LOGIC_IF_VH
`define PC_LOGIC_IF_VH

interface pc_logic_if;

	// Types
	`include "cpu_types_pkg.vh"

	
endinterface

`endif