/*
	Author: Mahesh Babu Gorantla, mgorantl@purdue.edu
	mg Account: mg226
	module: alu
	Description: This source code is used to design the alu for Lab-1 => This is a purely Combinational Block
*/

`include "../include/cpu_types_pkg.vh"
`include "../include/alu_if.vh"

import cpu_types_pkg::*;

module alu(
	alu_if.alu my_alu
);

	always_comb
	begin: OPERATION
		
	end

	always_comb
	begin: FLAGS

	end	

endmodule
